

module top(

	);



endmodule