module pe_tile(input [0 : 0] reset, input [31 : 0] config_data, input [31 : 0] config_addr, input [15 : 0] tile_id, input [0 : 0] clk);
endmodule