module switch_box(
                  output left_0,
                  input  left_1,
                  output left_2,
                  input  left_3,

                  input  right_0,
                  output right_1,
                  input  right_2,
                  output right_3,

                  input  top_0,
                  output top_1,
                  input  top_2,
                  output top_3,
                  
                  output bottom_0,
                  input  bottom_1,
                  output bottom_2,
                  input  bottom_3
                  );
   

endmodule // switch_box
