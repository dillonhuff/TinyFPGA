`include "pe_tile"
`include "io1in_pad"
`include "io1out_pad"


module top(
	input clk,
	input reset,
	input [31:0] config_addr,
	input [31:0] config_data,
	input in_wire_0,
	input in_wire_1,
	input in_wire_2,
	input in_wire_3,
	input in_wire_4,
	input in_wire_5,
	input in_wire_6,
	input in_wire_7,
	input in_wire_8,
	input in_wire_9,
	input in_wire_10,
	input in_wire_11,
	input in_wire_12,
	input in_wire_13,
	input in_wire_14,
	input in_wire_15,
	output out_wire_0,
	output out_wire_1,
	output out_wire_2,
	output out_wire_3,
	output out_wire_4,
	output out_wire_5,
	output out_wire_6,
	output out_wire_7,
	output out_wire_8,
	output out_wire_9,
	output out_wire_10,
	output out_wire_11,
	output out_wire_12,
	output out_wire_13,
	output out_wire_14,
	output out_wire_15
	);

	wire input_to_grid_0;
	wire input_to_grid_1;
	wire input_to_grid_2;
	wire input_to_grid_3;
	wire input_to_grid_4;
	wire input_to_grid_5;
	wire input_to_grid_6;
	wire input_to_grid_7;
	wire input_to_grid_8;
	wire input_to_grid_9;
	wire input_to_grid_10;
	wire input_to_grid_11;
	wire input_to_grid_12;
	wire input_to_grid_13;
	wire input_to_grid_14;
	wire input_to_grid_15;


	wire grid_to_output_0;
	wire grid_to_output_1;
	wire grid_to_output_2;
	wire grid_to_output_3;
	wire grid_to_output_4;
	wire grid_to_output_5;
	wire grid_to_output_6;
	wire grid_to_output_7;
	wire grid_to_output_8;
	wire grid_to_output_9;
	wire grid_to_output_10;
	wire grid_to_output_11;
	wire grid_to_output_12;
	wire grid_to_output_13;
	wire grid_to_output_14;
	wire grid_to_output_15;


	io1in_pad in_pad_0(
		.clk(clk),
		.top_pin(in_wire_0),
		.pin(input_to_grid_0)
	);

	io1in_pad in_pad_1(
		.clk(clk),
		.top_pin(in_wire_1),
		.pin(input_to_grid_1)
	);

	io1in_pad in_pad_2(
		.clk(clk),
		.top_pin(in_wire_2),
		.pin(input_to_grid_2)
	);

	io1in_pad in_pad_3(
		.clk(clk),
		.top_pin(in_wire_3),
		.pin(input_to_grid_3)
	);

	io1in_pad in_pad_4(
		.clk(clk),
		.top_pin(in_wire_4),
		.pin(input_to_grid_4)
	);

	io1in_pad in_pad_5(
		.clk(clk),
		.top_pin(in_wire_5),
		.pin(input_to_grid_5)
	);

	io1in_pad in_pad_6(
		.clk(clk),
		.top_pin(in_wire_6),
		.pin(input_to_grid_6)
	);

	io1in_pad in_pad_7(
		.clk(clk),
		.top_pin(in_wire_7),
		.pin(input_to_grid_7)
	);

	io1in_pad in_pad_8(
		.clk(clk),
		.top_pin(in_wire_8),
		.pin(input_to_grid_8)
	);

	io1in_pad in_pad_9(
		.clk(clk),
		.top_pin(in_wire_9),
		.pin(input_to_grid_9)
	);

	io1in_pad in_pad_10(
		.clk(clk),
		.top_pin(in_wire_10),
		.pin(input_to_grid_10)
	);

	io1in_pad in_pad_11(
		.clk(clk),
		.top_pin(in_wire_11),
		.pin(input_to_grid_11)
	);

	io1in_pad in_pad_12(
		.clk(clk),
		.top_pin(in_wire_12),
		.pin(input_to_grid_12)
	);

	io1in_pad in_pad_13(
		.clk(clk),
		.top_pin(in_wire_13),
		.pin(input_to_grid_13)
	);

	io1in_pad in_pad_14(
		.clk(clk),
		.top_pin(in_wire_14),
		.pin(input_to_grid_14)
	);

	io1in_pad in_pad_15(
		.clk(clk),
		.top_pin(in_wire_15),
		.pin(input_to_grid_15)
	);

	io1out_pad out_pad_0(
		.clk(clk),
		.top_pin(out_wire_0),
		.pin(grid_to_output_0)
	);

	io1out_pad out_pad_1(
		.clk(clk),
		.top_pin(out_wire_1),
		.pin(grid_to_output_1)
	);

	io1out_pad out_pad_2(
		.clk(clk),
		.top_pin(out_wire_2),
		.pin(grid_to_output_2)
	);

	io1out_pad out_pad_3(
		.clk(clk),
		.top_pin(out_wire_3),
		.pin(grid_to_output_3)
	);

	io1out_pad out_pad_4(
		.clk(clk),
		.top_pin(out_wire_4),
		.pin(grid_to_output_4)
	);

	io1out_pad out_pad_5(
		.clk(clk),
		.top_pin(out_wire_5),
		.pin(grid_to_output_5)
	);

	io1out_pad out_pad_6(
		.clk(clk),
		.top_pin(out_wire_6),
		.pin(grid_to_output_6)
	);

	io1out_pad out_pad_7(
		.clk(clk),
		.top_pin(out_wire_7),
		.pin(grid_to_output_7)
	);

	io1out_pad out_pad_8(
		.clk(clk),
		.top_pin(out_wire_8),
		.pin(grid_to_output_8)
	);

	io1out_pad out_pad_9(
		.clk(clk),
		.top_pin(out_wire_9),
		.pin(grid_to_output_9)
	);

	io1out_pad out_pad_10(
		.clk(clk),
		.top_pin(out_wire_10),
		.pin(grid_to_output_10)
	);

	io1out_pad out_pad_11(
		.clk(clk),
		.top_pin(out_wire_11),
		.pin(grid_to_output_11)
	);

	io1out_pad out_pad_12(
		.clk(clk),
		.top_pin(out_wire_12),
		.pin(grid_to_output_12)
	);

	io1out_pad out_pad_13(
		.clk(clk),
		.top_pin(out_wire_13),
		.pin(grid_to_output_13)
	);

	io1out_pad out_pad_14(
		.clk(clk),
		.top_pin(out_wire_14),
		.pin(grid_to_output_14)
	);

	io1out_pad out_pad_15(
		.clk(clk),
		.top_pin(out_wire_15),
		.pin(grid_to_output_15)
	);

	// PE tile grid
	pe_tile pe_tile_0_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1)
	);

	pe_tile pe_tile_0_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(2)
	);

	pe_tile pe_tile_0_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(3)
	);

	pe_tile pe_tile_0_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(4)
	);

	pe_tile pe_tile_0_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(5)
	);

	pe_tile pe_tile_0_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(6)
	);

	pe_tile pe_tile_0_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(7)
	);

	pe_tile pe_tile_0_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(8)
	);

	pe_tile pe_tile_0_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(9)
	);

	pe_tile pe_tile_0_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(10)
	);

	pe_tile pe_tile_0_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(11)
	);

	pe_tile pe_tile_0_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(12)
	);

	pe_tile pe_tile_0_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(13)
	);

	pe_tile pe_tile_0_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(14)
	);

	pe_tile pe_tile_0_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(15)
	);

	pe_tile pe_tile_0_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(16)
	);

	pe_tile pe_tile_1_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(17)
	);

	pe_tile pe_tile_1_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(18)
	);

	pe_tile pe_tile_1_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(19)
	);

	pe_tile pe_tile_1_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(20)
	);

	pe_tile pe_tile_1_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(21)
	);

	pe_tile pe_tile_1_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(22)
	);

	pe_tile pe_tile_1_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(23)
	);

	pe_tile pe_tile_1_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(24)
	);

	pe_tile pe_tile_1_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(25)
	);

	pe_tile pe_tile_1_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(26)
	);

	pe_tile pe_tile_1_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(27)
	);

	pe_tile pe_tile_1_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(28)
	);

	pe_tile pe_tile_1_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(29)
	);

	pe_tile pe_tile_1_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(30)
	);

	pe_tile pe_tile_1_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(31)
	);

	pe_tile pe_tile_1_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(32)
	);

	pe_tile pe_tile_2_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(33)
	);

	pe_tile pe_tile_2_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(34)
	);

	pe_tile pe_tile_2_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(35)
	);

	pe_tile pe_tile_2_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(36)
	);

	pe_tile pe_tile_2_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(37)
	);

	pe_tile pe_tile_2_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(38)
	);

	pe_tile pe_tile_2_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(39)
	);

	pe_tile pe_tile_2_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(40)
	);

	pe_tile pe_tile_2_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(41)
	);

	pe_tile pe_tile_2_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(42)
	);

	pe_tile pe_tile_2_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(43)
	);

	pe_tile pe_tile_2_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(44)
	);

	pe_tile pe_tile_2_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(45)
	);

	pe_tile pe_tile_2_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(46)
	);

	pe_tile pe_tile_2_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(47)
	);

	pe_tile pe_tile_2_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(48)
	);

	pe_tile pe_tile_3_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(49)
	);

	pe_tile pe_tile_3_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(50)
	);

	pe_tile pe_tile_3_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(51)
	);

	pe_tile pe_tile_3_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(52)
	);

	pe_tile pe_tile_3_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(53)
	);

	pe_tile pe_tile_3_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(54)
	);

	pe_tile pe_tile_3_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(55)
	);

	pe_tile pe_tile_3_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(56)
	);

	pe_tile pe_tile_3_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(57)
	);

	pe_tile pe_tile_3_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(58)
	);

	pe_tile pe_tile_3_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(59)
	);

	pe_tile pe_tile_3_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(60)
	);

	pe_tile pe_tile_3_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(61)
	);

	pe_tile pe_tile_3_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(62)
	);

	pe_tile pe_tile_3_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(63)
	);

	pe_tile pe_tile_3_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(64)
	);

	pe_tile pe_tile_4_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(65)
	);

	pe_tile pe_tile_4_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(66)
	);

	pe_tile pe_tile_4_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(67)
	);

	pe_tile pe_tile_4_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(68)
	);

	pe_tile pe_tile_4_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(69)
	);

	pe_tile pe_tile_4_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(70)
	);

	pe_tile pe_tile_4_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(71)
	);

	pe_tile pe_tile_4_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(72)
	);

	pe_tile pe_tile_4_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(73)
	);

	pe_tile pe_tile_4_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(74)
	);

	pe_tile pe_tile_4_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(75)
	);

	pe_tile pe_tile_4_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(76)
	);

	pe_tile pe_tile_4_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(77)
	);

	pe_tile pe_tile_4_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(78)
	);

	pe_tile pe_tile_4_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(79)
	);

	pe_tile pe_tile_4_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(80)
	);

	pe_tile pe_tile_5_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(81)
	);

	pe_tile pe_tile_5_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(82)
	);

	pe_tile pe_tile_5_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(83)
	);

	pe_tile pe_tile_5_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(84)
	);

	pe_tile pe_tile_5_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(85)
	);

	pe_tile pe_tile_5_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(86)
	);

	pe_tile pe_tile_5_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(87)
	);

	pe_tile pe_tile_5_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(88)
	);

	pe_tile pe_tile_5_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(89)
	);

	pe_tile pe_tile_5_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(90)
	);

	pe_tile pe_tile_5_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(91)
	);

	pe_tile pe_tile_5_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(92)
	);

	pe_tile pe_tile_5_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(93)
	);

	pe_tile pe_tile_5_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(94)
	);

	pe_tile pe_tile_5_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(95)
	);

	pe_tile pe_tile_5_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(96)
	);

	pe_tile pe_tile_6_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(97)
	);

	pe_tile pe_tile_6_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(98)
	);

	pe_tile pe_tile_6_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(99)
	);

	pe_tile pe_tile_6_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(100)
	);

	pe_tile pe_tile_6_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(101)
	);

	pe_tile pe_tile_6_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(102)
	);

	pe_tile pe_tile_6_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(103)
	);

	pe_tile pe_tile_6_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(104)
	);

	pe_tile pe_tile_6_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(105)
	);

	pe_tile pe_tile_6_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(106)
	);

	pe_tile pe_tile_6_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(107)
	);

	pe_tile pe_tile_6_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(108)
	);

	pe_tile pe_tile_6_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(109)
	);

	pe_tile pe_tile_6_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(110)
	);

	pe_tile pe_tile_6_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(111)
	);

	pe_tile pe_tile_6_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(112)
	);

	pe_tile pe_tile_7_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(113)
	);

	pe_tile pe_tile_7_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(114)
	);

	pe_tile pe_tile_7_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(115)
	);

	pe_tile pe_tile_7_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(116)
	);

	pe_tile pe_tile_7_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(117)
	);

	pe_tile pe_tile_7_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(118)
	);

	pe_tile pe_tile_7_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(119)
	);

	pe_tile pe_tile_7_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(120)
	);

	pe_tile pe_tile_7_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(121)
	);

	pe_tile pe_tile_7_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(122)
	);

	pe_tile pe_tile_7_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(123)
	);

	pe_tile pe_tile_7_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(124)
	);

	pe_tile pe_tile_7_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(125)
	);

	pe_tile pe_tile_7_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(126)
	);

	pe_tile pe_tile_7_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(127)
	);

	pe_tile pe_tile_7_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(128)
	);

	pe_tile pe_tile_8_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(129)
	);

	pe_tile pe_tile_8_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(130)
	);

	pe_tile pe_tile_8_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(131)
	);

	pe_tile pe_tile_8_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(132)
	);

	pe_tile pe_tile_8_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(133)
	);

	pe_tile pe_tile_8_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(134)
	);

	pe_tile pe_tile_8_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(135)
	);

	pe_tile pe_tile_8_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(136)
	);

	pe_tile pe_tile_8_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(137)
	);

	pe_tile pe_tile_8_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(138)
	);

	pe_tile pe_tile_8_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(139)
	);

	pe_tile pe_tile_8_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(140)
	);

	pe_tile pe_tile_8_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(141)
	);

	pe_tile pe_tile_8_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(142)
	);

	pe_tile pe_tile_8_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(143)
	);

	pe_tile pe_tile_8_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(144)
	);

	pe_tile pe_tile_9_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(145)
	);

	pe_tile pe_tile_9_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(146)
	);

	pe_tile pe_tile_9_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(147)
	);

	pe_tile pe_tile_9_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(148)
	);

	pe_tile pe_tile_9_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(149)
	);

	pe_tile pe_tile_9_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(150)
	);

	pe_tile pe_tile_9_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(151)
	);

	pe_tile pe_tile_9_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(152)
	);

	pe_tile pe_tile_9_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(153)
	);

	pe_tile pe_tile_9_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(154)
	);

	pe_tile pe_tile_9_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(155)
	);

	pe_tile pe_tile_9_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(156)
	);

	pe_tile pe_tile_9_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(157)
	);

	pe_tile pe_tile_9_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(158)
	);

	pe_tile pe_tile_9_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(159)
	);

	pe_tile pe_tile_9_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(160)
	);

	pe_tile pe_tile_10_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(161)
	);

	pe_tile pe_tile_10_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(162)
	);

	pe_tile pe_tile_10_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(163)
	);

	pe_tile pe_tile_10_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(164)
	);

	pe_tile pe_tile_10_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(165)
	);

	pe_tile pe_tile_10_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(166)
	);

	pe_tile pe_tile_10_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(167)
	);

	pe_tile pe_tile_10_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(168)
	);

	pe_tile pe_tile_10_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(169)
	);

	pe_tile pe_tile_10_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(170)
	);

	pe_tile pe_tile_10_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(171)
	);

	pe_tile pe_tile_10_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(172)
	);

	pe_tile pe_tile_10_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(173)
	);

	pe_tile pe_tile_10_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(174)
	);

	pe_tile pe_tile_10_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(175)
	);

	pe_tile pe_tile_10_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(176)
	);

	pe_tile pe_tile_11_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(177)
	);

	pe_tile pe_tile_11_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(178)
	);

	pe_tile pe_tile_11_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(179)
	);

	pe_tile pe_tile_11_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(180)
	);

	pe_tile pe_tile_11_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(181)
	);

	pe_tile pe_tile_11_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(182)
	);

	pe_tile pe_tile_11_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(183)
	);

	pe_tile pe_tile_11_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(184)
	);

	pe_tile pe_tile_11_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(185)
	);

	pe_tile pe_tile_11_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(186)
	);

	pe_tile pe_tile_11_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(187)
	);

	pe_tile pe_tile_11_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(188)
	);

	pe_tile pe_tile_11_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(189)
	);

	pe_tile pe_tile_11_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(190)
	);

	pe_tile pe_tile_11_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(191)
	);

	pe_tile pe_tile_11_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(192)
	);

	pe_tile pe_tile_12_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(193)
	);

	pe_tile pe_tile_12_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(194)
	);

	pe_tile pe_tile_12_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(195)
	);

	pe_tile pe_tile_12_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(196)
	);

	pe_tile pe_tile_12_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(197)
	);

	pe_tile pe_tile_12_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(198)
	);

	pe_tile pe_tile_12_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(199)
	);

	pe_tile pe_tile_12_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(200)
	);

	pe_tile pe_tile_12_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(201)
	);

	pe_tile pe_tile_12_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(202)
	);

	pe_tile pe_tile_12_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(203)
	);

	pe_tile pe_tile_12_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(204)
	);

	pe_tile pe_tile_12_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(205)
	);

	pe_tile pe_tile_12_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(206)
	);

	pe_tile pe_tile_12_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(207)
	);

	pe_tile pe_tile_12_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(208)
	);

	pe_tile pe_tile_13_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(209)
	);

	pe_tile pe_tile_13_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(210)
	);

	pe_tile pe_tile_13_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(211)
	);

	pe_tile pe_tile_13_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(212)
	);

	pe_tile pe_tile_13_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(213)
	);

	pe_tile pe_tile_13_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(214)
	);

	pe_tile pe_tile_13_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(215)
	);

	pe_tile pe_tile_13_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(216)
	);

	pe_tile pe_tile_13_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(217)
	);

	pe_tile pe_tile_13_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(218)
	);

	pe_tile pe_tile_13_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(219)
	);

	pe_tile pe_tile_13_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(220)
	);

	pe_tile pe_tile_13_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(221)
	);

	pe_tile pe_tile_13_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(222)
	);

	pe_tile pe_tile_13_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(223)
	);

	pe_tile pe_tile_13_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(224)
	);

	pe_tile pe_tile_14_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(225)
	);

	pe_tile pe_tile_14_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(226)
	);

	pe_tile pe_tile_14_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(227)
	);

	pe_tile pe_tile_14_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(228)
	);

	pe_tile pe_tile_14_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(229)
	);

	pe_tile pe_tile_14_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(230)
	);

	pe_tile pe_tile_14_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(231)
	);

	pe_tile pe_tile_14_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(232)
	);

	pe_tile pe_tile_14_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(233)
	);

	pe_tile pe_tile_14_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(234)
	);

	pe_tile pe_tile_14_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(235)
	);

	pe_tile pe_tile_14_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(236)
	);

	pe_tile pe_tile_14_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(237)
	);

	pe_tile pe_tile_14_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(238)
	);

	pe_tile pe_tile_14_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(239)
	);

	pe_tile pe_tile_14_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(240)
	);

	pe_tile pe_tile_15_0(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(241)
	);

	pe_tile pe_tile_15_1(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(242)
	);

	pe_tile pe_tile_15_2(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(243)
	);

	pe_tile pe_tile_15_3(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(244)
	);

	pe_tile pe_tile_15_4(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(245)
	);

	pe_tile pe_tile_15_5(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(246)
	);

	pe_tile pe_tile_15_6(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(247)
	);

	pe_tile pe_tile_15_7(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(248)
	);

	pe_tile pe_tile_15_8(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(249)
	);

	pe_tile pe_tile_15_9(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(250)
	);

	pe_tile pe_tile_15_10(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(251)
	);

	pe_tile pe_tile_15_11(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(252)
	);

	pe_tile pe_tile_15_12(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(253)
	);

	pe_tile pe_tile_15_13(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(254)
	);

	pe_tile pe_tile_15_14(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(255)
	);

	pe_tile pe_tile_15_15(
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(256)
	);



endmodule