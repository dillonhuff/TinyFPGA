module pe_tile();
   
endmodule
