`ifndef pe_tile_included
`define pe_tile_included 1
`include "pe_tile"
`endif

`ifndef io1in_pad_included
`define io1in_pad_included 1
`include "io1in_pad"
`endif

`ifndef io1out_pad_included
`define io1out_pad_included 1
`include "io1out_pad"
`endif



module top(
	input [0 : 0] reset,
	input [31 : 0] config_data,
	input [0 : 0] in_wire_2,
	input [0 : 0] in_wire_1,
	input [0 : 0] clk,
	input [0 : 0] in_wire_0,
	input [31 : 0] config_addr,
	output [0 : 0] out_wire_2,
	output [0 : 0] out_wire_1,
	output [0 : 0] out_wire_0
	);

	// Internal wires
	wire [1 - 1 : 0] wire_8;
	wire [1 - 1 : 0] wire_9;
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_0_2;
	wire [1 - 1 : 0] wire_42;
	wire [1 - 1 : 0] wire_0;
	wire [1 - 1 : 0] wire_1;
	wire [1 - 1 : 0] wire_2;
	wire [1 - 1 : 0] wire_3;
	wire [1 - 1 : 0] wire_4;
	wire [1 - 1 : 0] wire_5;
	wire [1 - 1 : 0] wire_6;
	wire [1 - 1 : 0] wire_7;
	wire [1 - 1 : 0] wire_47;
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_0_1;
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_0_0;
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_0_3;
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_0_2;
	wire [1 - 1 : 0] wire_22;
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_0_1_const;
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_1_0_const;
	wire [1 - 1 : 0] clk;
	wire [32 - 1 : 0] config_addr;
	wire [1 - 1 : 0] vertical_tile_0_0_to_tile_1_0_1;
	wire [1 - 1 : 0] vertical_tile_0_0_to_tile_1_0_0;
	wire [1 - 1 : 0] vertical_tile_0_0_to_tile_1_0_3;
	wire [1 - 1 : 0] vertical_tile_0_0_to_tile_1_0_2;
	wire [1 - 1 : 0] in_pad_2_pin_to_pe_tile_0_2_in_wire_3_0;
	wire [1 - 1 : 0] out_wire_2;
	wire [1 - 1 : 0] out_wire_1;
	wire [1 - 1 : 0] out_wire_0;
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_2_0_3;
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_0_2_0;
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_0_2_3;
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_0_2_2;
	wire [1 - 1 : 0] pe_tile_0_1_in_wire_3_3_const;
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_0_2_const;
	wire [1 - 1 : 0] pe_tile_2_0_in_wire_1_3_const;
	wire [1 - 1 : 0] pe_tile_0_0in_wire_2_1_const;
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_0_0_const;
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_2_1_3;
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_2_1_2;
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_2_1_1;
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_2_1_0;
	wire [1 - 1 : 0] pe_tile_0_0_in_wire_3_3_const;
	wire [1 - 1 : 0] out_pad_0_pin_to_pe_tile_2_0_out_wire_1_0;
	reg [1 - 1 : 0] pe_tile_0_2_id_wire;
	wire [1 - 1 : 0] in_wire_2;
	wire [1 - 1 : 0] in_wire_1;
	wire [1 - 1 : 0] in_wire_0;
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_0_3_const;
	wire [1 - 1 : 0] horizontal_tile_1_0_to_tile_1_1_1;
	wire [1 - 1 : 0] horizontal_tile_1_0_to_tile_1_1_0;
	wire [1 - 1 : 0] horizontal_tile_1_0_to_tile_1_1_3;
	wire [1 - 1 : 0] horizontal_tile_1_0_to_tile_1_1_2;
	wire [1 - 1 : 0] pe_tile_2_1_in_wire_1_2_const;
	wire [1 - 1 : 0] reset;
	wire [1 - 1 : 0] pe_tile_1_2_in_wire_0_2_const;
	wire [1 - 1 : 0] pe_tile_1_0in_wire_2_3_const;
	wire [1 - 1 : 0] wire_24;
	reg [1 - 1 : 0] pe_tile_0_1_id_wire;
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_0_1_1;
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_0_1_0;
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_0_1_3;
	wire [1 - 1 : 0] vertical_tile_1_1_to_tile_0_1_2;
	wire [1 - 1 : 0] horizontal_tile_0_2_to_tile_0_1_3;
	wire [1 - 1 : 0] horizontal_tile_0_2_to_tile_0_1_2;
	wire [1 - 1 : 0] horizontal_tile_0_2_to_tile_0_1_1;
	wire [1 - 1 : 0] horizontal_tile_0_2_to_tile_0_1_0;
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_0_1_const;
	wire [1 - 1 : 0] wire_49;
	wire [1 - 1 : 0] wire_48;
	wire [1 - 1 : 0] wire_43;
	reg [1 - 1 : 0] pe_tile_0_0_id_wire;
	wire [1 - 1 : 0] horizontal_tile_2_0_to_tile_2_1_1;
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_0_0;
	wire [1 - 1 : 0] horizontal_tile_2_0_to_tile_2_1_3;
	wire [1 - 1 : 0] horizontal_tile_2_0_to_tile_2_1_2;
	wire [1 - 1 : 0] wire_45;
	wire [1 - 1 : 0] pe_tile_1_0in_wire_2_0_const;
	wire [1 - 1 : 0] pe_tile_2_1_in_wire_1_3_const;
	wire [1 - 1 : 0] wire_46;
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_2_3;
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_2_2;
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_2_1;
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_2_0;
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_0_0_1;
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_0_0_0;
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_0_0_3;
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_0_0_2;
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_3_2_const;
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_3_1_const;
	wire [1 - 1 : 0] vertical_tile_2_1_to_tile_1_1_3;
	wire [1 - 1 : 0] vertical_tile_2_1_to_tile_1_1_2;
	wire [1 - 1 : 0] vertical_tile_2_1_to_tile_1_1_1;
	wire [1 - 1 : 0] vertical_tile_2_1_to_tile_1_1_0;
	wire [1 - 1 : 0] wire_52;
	wire [1 - 1 : 0] wire_53;
	wire [1 - 1 : 0] wire_50;
	reg [1 - 1 : 0] pe_tile_2_0_id_wire;
	wire [1 - 1 : 0] pe_tile_0_0_in_wire_3_1_const;
	wire [1 - 1 : 0] in_pad_1_pin_to_pe_tile_0_1_in_wire_3_0;
	wire [1 - 1 : 0] pe_tile_2_0_in_wire_1_2_const;
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_0_0_const;
	wire [1 - 1 : 0] pe_tile_2_0_in_wire_1_0_const;
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_1_1_const;
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_2_2_3;
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_2_2_2;
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_2_2_1;
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_2_2_0;
	wire [1 - 1 : 0] pe_tile_2_1_in_wire_1_1_const;
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_1_3_const;
	wire [1 - 1 : 0] wire_51;
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_0_3_const;
	wire [1 - 1 : 0] wire_23;
	wire [1 - 1 : 0] wire_12;
	wire [1 - 1 : 0] wire_21;
	wire [1 - 1 : 0] wire_20;
	wire [1 - 1 : 0] wire_27;
	wire [1 - 1 : 0] wire_26;
	wire [1 - 1 : 0] wire_25;
	wire [1 - 1 : 0] pe_tile_0_1_in_wire_3_2_const;
	wire [1 - 1 : 0] pe_tile_2_2_in_wire_1_2_const;
	wire [1 - 1 : 0] wire_29;
	wire [1 - 1 : 0] wire_28;
	wire [1 - 1 : 0] wire_10;
	wire [1 - 1 : 0] wire_11;
	wire [1 - 1 : 0] pe_tile_1_2_in_wire_0_0_const;
	wire [1 - 1 : 0] pe_tile_2_0in_wire_2_1_const;
	wire [1 - 1 : 0] pe_tile_0_1_in_wire_3_1_const;
	wire [1 - 1 : 0] vertical_tile_2_0_to_tile_1_0_3;
	wire [1 - 1 : 0] vertical_tile_2_0_to_tile_1_0_2;
	wire [1 - 1 : 0] vertical_tile_2_0_to_tile_1_0_1;
	wire [1 - 1 : 0] vertical_tile_2_0_to_tile_1_0_0;
	wire [1 - 1 : 0] pe_tile_1_2_in_wire_0_3_const;
	reg [1 - 1 : 0] pe_tile_1_1_id_wire;
	wire [1 - 1 : 0] vertical_tile_2_2_to_tile_1_2_3;
	wire [1 - 1 : 0] vertical_tile_2_2_to_tile_1_2_2;
	wire [1 - 1 : 0] vertical_tile_2_2_to_tile_1_2_1;
	wire [1 - 1 : 0] vertical_tile_0_1_to_tile_1_1_2;
	wire [1 - 1 : 0] wire_34;
	wire [1 - 1 : 0] wire_35;
	wire [1 - 1 : 0] wire_36;
	wire [1 - 1 : 0] wire_37;
	wire [1 - 1 : 0] wire_38;
	wire [1 - 1 : 0] wire_39;
	reg [1 - 1 : 0] pe_tile_2_2_id_wire;
	wire [1 - 1 : 0] vertical_tile_0_2_to_tile_1_2_1;
	wire [1 - 1 : 0] vertical_tile_0_2_to_tile_1_2_0;
	wire [1 - 1 : 0] vertical_tile_0_2_to_tile_1_2_3;
	wire [1 - 1 : 0] vertical_tile_0_2_to_tile_1_2_2;
	reg [1 - 1 : 0] pe_tile_2_1_id_wire;
	wire [1 - 1 : 0] pe_tile_0_0in_wire_2_0_const;
	wire [1 - 1 : 0] pe_tile_2_1_in_wire_1_0_const;
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_2_0;
	wire [1 - 1 : 0] horizontal_tile_2_2_to_tile_2_1_3;
	wire [1 - 1 : 0] horizontal_tile_2_2_to_tile_2_1_2;
	wire [1 - 1 : 0] horizontal_tile_2_2_to_tile_2_1_1;
	wire [1 - 1 : 0] horizontal_tile_2_2_to_tile_2_1_0;
	wire [1 - 1 : 0] pe_tile_1_0in_wire_2_2_const;
	wire [1 - 1 : 0] in_pad_0_pin_to_pe_tile_0_0_in_wire_3_0;
	wire [1 - 1 : 0] pe_tile_2_0in_wire_2_0_const;
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_3_3_const;
	wire [1 - 1 : 0] vertical_tile_1_2_to_tile_0_2_1;
	wire [1 - 1 : 0] pe_tile_0_2_in_wire_0_2_const;
	wire [1 - 1 : 0] pe_tile_0_0_in_wire_3_2_const;
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_2_0_2;
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_0_1;
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_0_0;
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_0_3;
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_0_2;
	wire [32 - 1 : 0] config_data;
	wire [1 - 1 : 0] wire_30;
	wire [1 - 1 : 0] pe_tile_0_0in_wire_2_3_const;
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_2_0_0;
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_2_3;
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_2_2;
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_2_1;
	wire [1 - 1 : 0] horizontal_tile_1_1_to_tile_1_2_0;
	wire [1 - 1 : 0] pe_tile_2_0in_wire_2_3_const;
	wire [1 - 1 : 0] out_pad_1_pin_to_pe_tile_2_1_out_wire_1_0;
	wire [1 - 1 : 0] pe_tile_2_0in_wire_2_2_const;
	wire [1 - 1 : 0] wire_41;
	wire [1 - 1 : 0] wire_31;
	wire [1 - 1 : 0] pe_tile_1_2_in_wire_0_1_const;
	wire [1 - 1 : 0] out_pad_2_pin_to_pe_tile_2_2_out_wire_1_0;
	wire [1 - 1 : 0] pe_tile_2_0_in_wire_1_1_const;
	wire [1 - 1 : 0] wire_13;
	wire [1 - 1 : 0] pe_tile_0_0in_wire_2_2_const;
	wire [1 - 1 : 0] horizontal_tile_1_2_to_tile_1_1_3;
	wire [1 - 1 : 0] horizontal_tile_1_2_to_tile_1_1_2;
	wire [1 - 1 : 0] horizontal_tile_1_2_to_tile_1_1_1;
	wire [1 - 1 : 0] horizontal_tile_1_2_to_tile_1_1_0;
	wire [1 - 1 : 0] wire_40;
	reg [1 - 1 : 0] pe_tile_1_0_id_wire;
	wire [1 - 1 : 0] wire_32;
	reg [1 - 1 : 0] pe_tile_1_2_id_wire;
	wire [1 - 1 : 0] wire_18;
	wire [1 - 1 : 0] wire_19;
	wire [1 - 1 : 0] vertical_tile_1_0_to_tile_2_0_1;
	wire [1 - 1 : 0] pe_tile_1_0in_wire_2_1_const;
	wire [1 - 1 : 0] horizontal_tile_0_0_to_tile_0_1_1;
	wire [1 - 1 : 0] horizontal_tile_0_0_to_tile_0_1_0;
	wire [1 - 1 : 0] horizontal_tile_0_0_to_tile_0_1_3;
	wire [1 - 1 : 0] horizontal_tile_0_0_to_tile_0_1_2;
	wire [1 - 1 : 0] wire_16;
	wire [1 - 1 : 0] wire_17;
	wire [1 - 1 : 0] wire_14;
	wire [1 - 1 : 0] wire_15;
	wire [1 - 1 : 0] vertical_tile_0_1_to_tile_1_1_1;
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_2_3;
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_2_2;
	wire [1 - 1 : 0] horizontal_tile_0_1_to_tile_0_2_1;
	wire [1 - 1 : 0] vertical_tile_0_1_to_tile_1_1_0;
	wire [1 - 1 : 0] wire_33;
	wire [1 - 1 : 0] vertical_tile_0_1_to_tile_1_1_3;
	wire [1 - 1 : 0] wire_44;
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_0_1;
	wire [1 - 1 : 0] vertical_tile_2_2_to_tile_1_2_0;
	wire [1 - 1 : 0] horizontal_tile_2_0_to_tile_2_1_0;
	wire [1 - 1 : 0] horizontal_tile_2_1_to_tile_2_0_3;
	// End of wire declarations

	io1out_pad out_pad_2(
		.top_pin(out_wire_2),
		.clk(clk),
		.pin(out_pad_2_pin_to_pe_tile_2_2_out_wire_1_0)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0_in_wire_3_3_const_2(
		.out(pe_tile_0_0_in_wire_3_3_const),
		.in(wire_2)
	);

	io1out_pad out_pad_0(
		.top_pin(out_wire_0),
		.clk(clk),
		.pin(out_pad_0_pin_to_pe_tile_2_0_out_wire_1_0)
	);

	io1out_pad out_pad_1(
		.top_pin(out_wire_1),
		.clk(clk),
		.pin(out_pad_1_pin_to_pe_tile_2_1_out_wire_1_0)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_0in_wire_2_1_const_21(
		.out(pe_tile_1_0in_wire_2_1_const),
		.in(wire_21)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_1_in_wire_3_2_const_9(
		.out(pe_tile_0_1_in_wire_3_2_const),
		.in(wire_9)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_1_in_wire_1_0_const_40(
		.out(pe_tile_2_1_in_wire_1_0_const),
		.in(wire_40)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_2_in_wire_3_3_const_14_const(
		.out(wire_14)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0in_wire_2_3_const_38(
		.out(pe_tile_2_0in_wire_2_3_const),
		.in(wire_38)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0_in_wire_1_0_const_31(
		.out(pe_tile_2_0_in_wire_1_0_const),
		.in(wire_31)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_0_in_wire_3_3_const_2_const(
		.out(wire_2)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_id_wire_19(
		.out(pe_tile_0_2_id_wire),
		.in(wire_19)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_2_in_wire_0_0_const_26(
		.out(pe_tile_1_2_in_wire_0_0_const),
		.in(wire_26)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_1_in_wire_3_3_const_10(
		.out(pe_tile_0_1_in_wire_3_3_const),
		.in(wire_10)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_2_in_wire_0_2_const_51_const(
		.out(wire_51)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_2_in_wire_0_1_const_50_const(
		.out(wire_50)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_0_in_wire_3_1_const_0_const(
		.out(wire_0)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0in_wire_2_1_const_4(
		.out(pe_tile_0_0in_wire_2_1_const),
		.in(wire_4)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_1_in_wire_1_2_const_42(
		.out(pe_tile_2_1_in_wire_1_2_const),
		.in(wire_42)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_1_2_const_47(
		.out(pe_tile_2_2_in_wire_1_2_const),
		.in(wire_47)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_0in_wire_2_0_const_20(
		.out(pe_tile_1_0in_wire_2_0_const),
		.in(wire_20)
	);

	const_mod #(.width(1), .value(3))  assign_pe_tile_0_2_id_wire_19_const(
		.out(wire_19)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_2_in_wire_0_3_const_52_const(
		.out(wire_52)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_2_in_wire_1_2_const_47_const(
		.out(wire_47)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_1_0in_wire_2_0_const_20_const(
		.out(wire_20)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0in_wire_2_1_const_36(
		.out(pe_tile_2_0in_wire_2_1_const),
		.in(wire_36)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_0_in_wire_1_0_const_31_const(
		.out(wire_31)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_0_2_const_17(
		.out(pe_tile_0_2_in_wire_0_2_const),
		.in(wire_17)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_1_id_wire_11(
		.out(pe_tile_0_1_id_wire),
		.in(wire_11)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_1_id_wire_25(
		.out(pe_tile_1_1_id_wire),
		.in(wire_25)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_2_in_wire_3_1_const_12_const(
		.out(wire_12)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_2_in_wire_0_0_const_49_const(
		.out(wire_49)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_0in_wire_2_2_const_37_const(
		.out(wire_37)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_1_0in_wire_2_3_const_23_const(
		.out(wire_23)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0in_wire_2_0_const_3(
		.out(pe_tile_0_0in_wire_2_0_const),
		.in(wire_3)
	);

	pe_tile_right pe_tile_1_2(
		.out_wire_3_0(vertical_tile_1_2_to_tile_0_2_0),
		.out_wire_3_1(vertical_tile_1_2_to_tile_0_2_1),
		.out_wire_3_2(vertical_tile_1_2_to_tile_0_2_2),
		.out_wire_3_3(vertical_tile_1_2_to_tile_0_2_3),
		.in_wire_3_0(vertical_tile_0_2_to_tile_1_2_0),
		.in_wire_3_1(vertical_tile_0_2_to_tile_1_2_1),
		.in_wire_3_2(vertical_tile_0_2_to_tile_1_2_2),
		.in_wire_3_3(vertical_tile_0_2_to_tile_1_2_3),
		.out_wire_1_0(vertical_tile_1_2_to_tile_2_2_0),
		.out_wire_1_1(vertical_tile_1_2_to_tile_2_2_1),
		.out_wire_1_2(vertical_tile_1_2_to_tile_2_2_2),
		.out_wire_1_3(vertical_tile_1_2_to_tile_2_2_3),
		.in_wire_1_0(vertical_tile_2_2_to_tile_1_2_0),
		.in_wire_1_1(vertical_tile_2_2_to_tile_1_2_1),
		.in_wire_1_2(vertical_tile_2_2_to_tile_1_2_2),
		.in_wire_1_3(vertical_tile_2_2_to_tile_1_2_3),
		.out_wire_2_0(horizontal_tile_1_2_to_tile_1_1_0),
		.out_wire_2_1(horizontal_tile_1_2_to_tile_1_1_1),
		.out_wire_2_2(horizontal_tile_1_2_to_tile_1_1_2),
		.out_wire_2_3(horizontal_tile_1_2_to_tile_1_1_3),
		.in_wire_2_0(horizontal_tile_1_1_to_tile_1_2_0),
		.in_wire_2_1(horizontal_tile_1_1_to_tile_1_2_1),
		.in_wire_2_2(horizontal_tile_1_1_to_tile_1_2_2),
		.in_wire_2_3(horizontal_tile_1_1_to_tile_1_2_3),
		.in_wire_0_0(pe_tile_1_2_in_wire_0_0_const),
		.in_wire_0_1(pe_tile_1_2_in_wire_0_1_const),
		.in_wire_0_2(pe_tile_1_2_in_wire_0_2_const),
		.in_wire_0_3(pe_tile_1_2_in_wire_0_3_const),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_1_2_id_wire)
	);

	pe_tile_left pe_tile_1_0(
		.out_wire_3_0(vertical_tile_1_0_to_tile_0_0_0),
		.out_wire_3_1(vertical_tile_1_0_to_tile_0_0_1),
		.out_wire_3_2(vertical_tile_1_0_to_tile_0_0_2),
		.out_wire_3_3(vertical_tile_1_0_to_tile_0_0_3),
		.in_wire_3_0(vertical_tile_0_0_to_tile_1_0_0),
		.in_wire_3_1(vertical_tile_0_0_to_tile_1_0_1),
		.in_wire_3_2(vertical_tile_0_0_to_tile_1_0_2),
		.in_wire_3_3(vertical_tile_0_0_to_tile_1_0_3),
		.out_wire_1_0(vertical_tile_1_0_to_tile_2_0_0),
		.out_wire_1_1(vertical_tile_1_0_to_tile_2_0_1),
		.out_wire_1_2(vertical_tile_1_0_to_tile_2_0_2),
		.out_wire_1_3(vertical_tile_1_0_to_tile_2_0_3),
		.in_wire_1_0(vertical_tile_2_0_to_tile_1_0_0),
		.in_wire_1_1(vertical_tile_2_0_to_tile_1_0_1),
		.in_wire_1_2(vertical_tile_2_0_to_tile_1_0_2),
		.in_wire_1_3(vertical_tile_2_0_to_tile_1_0_3),
		.in_wire_2_0(pe_tile_1_0in_wire_2_0_const),
		.in_wire_2_1(pe_tile_1_0in_wire_2_1_const),
		.in_wire_2_2(pe_tile_1_0in_wire_2_2_const),
		.in_wire_2_3(pe_tile_1_0in_wire_2_3_const),
		.out_wire_0_0(horizontal_tile_1_0_to_tile_1_1_0),
		.out_wire_0_1(horizontal_tile_1_0_to_tile_1_1_1),
		.out_wire_0_2(horizontal_tile_1_0_to_tile_1_1_2),
		.out_wire_0_3(horizontal_tile_1_0_to_tile_1_1_3),
		.in_wire_0_0(horizontal_tile_1_1_to_tile_1_0_0),
		.in_wire_0_1(horizontal_tile_1_1_to_tile_1_0_1),
		.in_wire_0_2(horizontal_tile_1_1_to_tile_1_0_2),
		.in_wire_0_3(horizontal_tile_1_1_to_tile_1_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_1_0_id_wire)
	);

	pe_tile pe_tile_1_1(
		.out_wire_3_0(vertical_tile_1_1_to_tile_0_1_0),
		.out_wire_3_1(vertical_tile_1_1_to_tile_0_1_1),
		.out_wire_3_2(vertical_tile_1_1_to_tile_0_1_2),
		.out_wire_3_3(vertical_tile_1_1_to_tile_0_1_3),
		.in_wire_3_0(vertical_tile_0_1_to_tile_1_1_0),
		.in_wire_3_1(vertical_tile_0_1_to_tile_1_1_1),
		.in_wire_3_2(vertical_tile_0_1_to_tile_1_1_2),
		.in_wire_3_3(vertical_tile_0_1_to_tile_1_1_3),
		.out_wire_1_0(vertical_tile_1_1_to_tile_2_1_0),
		.out_wire_1_1(vertical_tile_1_1_to_tile_2_1_1),
		.out_wire_1_2(vertical_tile_1_1_to_tile_2_1_2),
		.out_wire_1_3(vertical_tile_1_1_to_tile_2_1_3),
		.in_wire_1_0(vertical_tile_2_1_to_tile_1_1_0),
		.in_wire_1_1(vertical_tile_2_1_to_tile_1_1_1),
		.in_wire_1_2(vertical_tile_2_1_to_tile_1_1_2),
		.in_wire_1_3(vertical_tile_2_1_to_tile_1_1_3),
		.out_wire_2_0(horizontal_tile_1_1_to_tile_1_0_0),
		.out_wire_2_1(horizontal_tile_1_1_to_tile_1_0_1),
		.out_wire_2_2(horizontal_tile_1_1_to_tile_1_0_2),
		.out_wire_2_3(horizontal_tile_1_1_to_tile_1_0_3),
		.in_wire_2_0(horizontal_tile_1_0_to_tile_1_1_0),
		.in_wire_2_1(horizontal_tile_1_0_to_tile_1_1_1),
		.in_wire_2_2(horizontal_tile_1_0_to_tile_1_1_2),
		.in_wire_2_3(horizontal_tile_1_0_to_tile_1_1_3),
		.out_wire_0_0(horizontal_tile_1_1_to_tile_1_2_0),
		.out_wire_0_1(horizontal_tile_1_1_to_tile_1_2_1),
		.out_wire_0_2(horizontal_tile_1_1_to_tile_1_2_2),
		.out_wire_0_3(horizontal_tile_1_1_to_tile_1_2_3),
		.in_wire_0_0(horizontal_tile_1_2_to_tile_1_1_0),
		.in_wire_0_1(horizontal_tile_1_2_to_tile_1_1_1),
		.in_wire_0_2(horizontal_tile_1_2_to_tile_1_1_2),
		.in_wire_0_3(horizontal_tile_1_2_to_tile_1_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_1_1_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0in_wire_2_0_const_35(
		.out(pe_tile_2_0in_wire_2_0_const),
		.in(wire_35)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0in_wire_2_3_const_6(
		.out(pe_tile_0_0in_wire_2_3_const),
		.in(wire_6)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_2_in_wire_1_0_const_45_const(
		.out(wire_45)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_0_1_const_50(
		.out(pe_tile_2_2_in_wire_0_1_const),
		.in(wire_50)
	);

	const_mod #(.width(1), .value(5))  assign_pe_tile_1_1_id_wire_25_const(
		.out(wire_25)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_2_in_wire_1_3_const_48_const(
		.out(wire_48)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_1_in_wire_1_1_const_41_const(
		.out(wire_41)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_1_in_wire_1_0_const_40_const(
		.out(wire_40)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_1_0in_wire_2_2_const_22_const(
		.out(wire_22)
	);

	const_mod #(.width(1), .value(7))  assign_pe_tile_2_0_id_wire_39_const(
		.out(wire_39)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0_id_wire_7(
		.out(pe_tile_0_0_id_wire),
		.in(wire_7)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0_in_wire_1_1_const_32(
		.out(pe_tile_2_0_in_wire_1_1_const),
		.in(wire_32)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_0in_wire_2_1_const_36_const(
		.out(wire_36)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_1_in_wire_3_1_const_8_const(
		.out(wire_8)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_1_2_in_wire_0_3_const_29_const(
		.out(wire_29)
	);

	const_mod #(.width(1), .value(2))  assign_pe_tile_0_1_id_wire_11_const(
		.out(wire_11)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_1_3_const_48(
		.out(pe_tile_2_2_in_wire_1_3_const),
		.in(wire_48)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_2_in_wire_1_1_const_46_const(
		.out(wire_46)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_0_2_const_51(
		.out(pe_tile_2_2_in_wire_0_2_const),
		.in(wire_51)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_0_0_const_49(
		.out(pe_tile_2_2_in_wire_0_0_const),
		.in(wire_49)
	);

	pe_tile_bottom_left pe_tile_2_0(
		.out_wire_3_0(vertical_tile_2_0_to_tile_1_0_0),
		.out_wire_3_1(vertical_tile_2_0_to_tile_1_0_1),
		.out_wire_3_2(vertical_tile_2_0_to_tile_1_0_2),
		.out_wire_3_3(vertical_tile_2_0_to_tile_1_0_3),
		.in_wire_3_0(vertical_tile_1_0_to_tile_2_0_0),
		.in_wire_3_1(vertical_tile_1_0_to_tile_2_0_1),
		.in_wire_3_2(vertical_tile_1_0_to_tile_2_0_2),
		.in_wire_3_3(vertical_tile_1_0_to_tile_2_0_3),
		.out_wire_1_0(out_pad_0_pin_to_pe_tile_2_0_out_wire_1_0),
		.in_wire_1_0(pe_tile_2_0_in_wire_1_0_const),
		.in_wire_1_1(pe_tile_2_0_in_wire_1_1_const),
		.in_wire_1_2(pe_tile_2_0_in_wire_1_2_const),
		.in_wire_1_3(pe_tile_2_0_in_wire_1_3_const),
		.in_wire_2_0(pe_tile_2_0in_wire_2_0_const),
		.in_wire_2_1(pe_tile_2_0in_wire_2_1_const),
		.in_wire_2_2(pe_tile_2_0in_wire_2_2_const),
		.in_wire_2_3(pe_tile_2_0in_wire_2_3_const),
		.out_wire_0_0(horizontal_tile_2_0_to_tile_2_1_0),
		.out_wire_0_1(horizontal_tile_2_0_to_tile_2_1_1),
		.out_wire_0_2(horizontal_tile_2_0_to_tile_2_1_2),
		.out_wire_0_3(horizontal_tile_2_0_to_tile_2_1_3),
		.in_wire_0_0(horizontal_tile_2_1_to_tile_2_0_0),
		.in_wire_0_1(horizontal_tile_2_1_to_tile_2_0_1),
		.in_wire_0_2(horizontal_tile_2_1_to_tile_2_0_2),
		.in_wire_0_3(horizontal_tile_2_1_to_tile_2_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_2_0_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_1_in_wire_1_1_const_41(
		.out(pe_tile_2_1_in_wire_1_1_const),
		.in(wire_41)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_1_id_wire_44(
		.out(pe_tile_2_1_id_wire),
		.in(wire_44)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_0_in_wire_1_2_const_33_const(
		.out(wire_33)
	);

	pe_tile_bottom_right pe_tile_2_2(
		.out_wire_3_0(vertical_tile_2_2_to_tile_1_2_0),
		.out_wire_3_1(vertical_tile_2_2_to_tile_1_2_1),
		.out_wire_3_2(vertical_tile_2_2_to_tile_1_2_2),
		.out_wire_3_3(vertical_tile_2_2_to_tile_1_2_3),
		.in_wire_3_0(vertical_tile_1_2_to_tile_2_2_0),
		.in_wire_3_1(vertical_tile_1_2_to_tile_2_2_1),
		.in_wire_3_2(vertical_tile_1_2_to_tile_2_2_2),
		.in_wire_3_3(vertical_tile_1_2_to_tile_2_2_3),
		.out_wire_1_0(out_pad_2_pin_to_pe_tile_2_2_out_wire_1_0),
		.in_wire_1_0(pe_tile_2_2_in_wire_1_0_const),
		.in_wire_1_1(pe_tile_2_2_in_wire_1_1_const),
		.in_wire_1_2(pe_tile_2_2_in_wire_1_2_const),
		.in_wire_1_3(pe_tile_2_2_in_wire_1_3_const),
		.out_wire_2_0(horizontal_tile_2_2_to_tile_2_1_0),
		.out_wire_2_1(horizontal_tile_2_2_to_tile_2_1_1),
		.out_wire_2_2(horizontal_tile_2_2_to_tile_2_1_2),
		.out_wire_2_3(horizontal_tile_2_2_to_tile_2_1_3),
		.in_wire_2_0(horizontal_tile_2_1_to_tile_2_2_0),
		.in_wire_2_1(horizontal_tile_2_1_to_tile_2_2_1),
		.in_wire_2_2(horizontal_tile_2_1_to_tile_2_2_2),
		.in_wire_2_3(horizontal_tile_2_1_to_tile_2_2_3),
		.in_wire_0_0(pe_tile_2_2_in_wire_0_0_const),
		.in_wire_0_1(pe_tile_2_2_in_wire_0_1_const),
		.in_wire_0_2(pe_tile_2_2_in_wire_0_2_const),
		.in_wire_0_3(pe_tile_2_2_in_wire_0_3_const),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_2_2_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_1_in_wire_3_1_const_8(
		.out(pe_tile_0_1_in_wire_3_1_const),
		.in(wire_8)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_0in_wire_2_2_const_5_const(
		.out(wire_5)
	);

	const_mod #(.width(1), .value(4))  assign_pe_tile_1_0_id_wire_24_const(
		.out(wire_24)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0in_wire_2_2_const_5(
		.out(pe_tile_0_0in_wire_2_2_const),
		.in(wire_5)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_0in_wire_2_2_const_22(
		.out(pe_tile_1_0in_wire_2_2_const),
		.in(wire_22)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_2_in_wire_0_2_const_28(
		.out(pe_tile_1_2_in_wire_0_2_const),
		.in(wire_28)
	);

	pe_tile_top_right pe_tile_0_2(
		.in_wire_3_0(in_pad_2_pin_to_pe_tile_0_2_in_wire_3_0),
		.in_wire_3_1(pe_tile_0_2_in_wire_3_1_const),
		.in_wire_3_2(pe_tile_0_2_in_wire_3_2_const),
		.in_wire_3_3(pe_tile_0_2_in_wire_3_3_const),
		.out_wire_1_0(vertical_tile_0_2_to_tile_1_2_0),
		.out_wire_1_1(vertical_tile_0_2_to_tile_1_2_1),
		.out_wire_1_2(vertical_tile_0_2_to_tile_1_2_2),
		.out_wire_1_3(vertical_tile_0_2_to_tile_1_2_3),
		.in_wire_1_0(vertical_tile_1_2_to_tile_0_2_0),
		.in_wire_1_1(vertical_tile_1_2_to_tile_0_2_1),
		.in_wire_1_2(vertical_tile_1_2_to_tile_0_2_2),
		.in_wire_1_3(vertical_tile_1_2_to_tile_0_2_3),
		.out_wire_2_0(horizontal_tile_0_2_to_tile_0_1_0),
		.out_wire_2_1(horizontal_tile_0_2_to_tile_0_1_1),
		.out_wire_2_2(horizontal_tile_0_2_to_tile_0_1_2),
		.out_wire_2_3(horizontal_tile_0_2_to_tile_0_1_3),
		.in_wire_2_0(horizontal_tile_0_1_to_tile_0_2_0),
		.in_wire_2_1(horizontal_tile_0_1_to_tile_0_2_1),
		.in_wire_2_2(horizontal_tile_0_1_to_tile_0_2_2),
		.in_wire_2_3(horizontal_tile_0_1_to_tile_0_2_3),
		.in_wire_0_0(pe_tile_0_2_in_wire_0_0_const),
		.in_wire_0_1(pe_tile_0_2_in_wire_0_1_const),
		.in_wire_0_2(pe_tile_0_2_in_wire_0_2_const),
		.in_wire_0_3(pe_tile_0_2_in_wire_0_3_const),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_0_2_id_wire)
	);

	pe_tile_top pe_tile_0_1(
		.in_wire_3_0(in_pad_1_pin_to_pe_tile_0_1_in_wire_3_0),
		.in_wire_3_1(pe_tile_0_1_in_wire_3_1_const),
		.in_wire_3_2(pe_tile_0_1_in_wire_3_2_const),
		.in_wire_3_3(pe_tile_0_1_in_wire_3_3_const),
		.out_wire_1_0(vertical_tile_0_1_to_tile_1_1_0),
		.out_wire_1_1(vertical_tile_0_1_to_tile_1_1_1),
		.out_wire_1_2(vertical_tile_0_1_to_tile_1_1_2),
		.out_wire_1_3(vertical_tile_0_1_to_tile_1_1_3),
		.in_wire_1_0(vertical_tile_1_1_to_tile_0_1_0),
		.in_wire_1_1(vertical_tile_1_1_to_tile_0_1_1),
		.in_wire_1_2(vertical_tile_1_1_to_tile_0_1_2),
		.in_wire_1_3(vertical_tile_1_1_to_tile_0_1_3),
		.out_wire_2_0(horizontal_tile_0_1_to_tile_0_0_0),
		.out_wire_2_1(horizontal_tile_0_1_to_tile_0_0_1),
		.out_wire_2_2(horizontal_tile_0_1_to_tile_0_0_2),
		.out_wire_2_3(horizontal_tile_0_1_to_tile_0_0_3),
		.in_wire_2_0(horizontal_tile_0_0_to_tile_0_1_0),
		.in_wire_2_1(horizontal_tile_0_0_to_tile_0_1_1),
		.in_wire_2_2(horizontal_tile_0_0_to_tile_0_1_2),
		.in_wire_2_3(horizontal_tile_0_0_to_tile_0_1_3),
		.out_wire_0_0(horizontal_tile_0_1_to_tile_0_2_0),
		.out_wire_0_1(horizontal_tile_0_1_to_tile_0_2_1),
		.out_wire_0_2(horizontal_tile_0_1_to_tile_0_2_2),
		.out_wire_0_3(horizontal_tile_0_1_to_tile_0_2_3),
		.in_wire_0_0(horizontal_tile_0_2_to_tile_0_1_0),
		.in_wire_0_1(horizontal_tile_0_2_to_tile_0_1_1),
		.in_wire_0_2(horizontal_tile_0_2_to_tile_0_1_2),
		.in_wire_0_3(horizontal_tile_0_2_to_tile_0_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_0_1_id_wire)
	);

	pe_tile_top_left pe_tile_0_0(
		.in_wire_3_0(in_pad_0_pin_to_pe_tile_0_0_in_wire_3_0),
		.in_wire_3_1(pe_tile_0_0_in_wire_3_1_const),
		.in_wire_3_2(pe_tile_0_0_in_wire_3_2_const),
		.in_wire_3_3(pe_tile_0_0_in_wire_3_3_const),
		.out_wire_1_0(vertical_tile_0_0_to_tile_1_0_0),
		.out_wire_1_1(vertical_tile_0_0_to_tile_1_0_1),
		.out_wire_1_2(vertical_tile_0_0_to_tile_1_0_2),
		.out_wire_1_3(vertical_tile_0_0_to_tile_1_0_3),
		.in_wire_1_0(vertical_tile_1_0_to_tile_0_0_0),
		.in_wire_1_1(vertical_tile_1_0_to_tile_0_0_1),
		.in_wire_1_2(vertical_tile_1_0_to_tile_0_0_2),
		.in_wire_1_3(vertical_tile_1_0_to_tile_0_0_3),
		.in_wire_2_0(pe_tile_0_0in_wire_2_0_const),
		.in_wire_2_1(pe_tile_0_0in_wire_2_1_const),
		.in_wire_2_2(pe_tile_0_0in_wire_2_2_const),
		.in_wire_2_3(pe_tile_0_0in_wire_2_3_const),
		.out_wire_0_0(horizontal_tile_0_0_to_tile_0_1_0),
		.out_wire_0_1(horizontal_tile_0_0_to_tile_0_1_1),
		.out_wire_0_2(horizontal_tile_0_0_to_tile_0_1_2),
		.out_wire_0_3(horizontal_tile_0_0_to_tile_0_1_3),
		.in_wire_0_0(horizontal_tile_0_1_to_tile_0_0_0),
		.in_wire_0_1(horizontal_tile_0_1_to_tile_0_0_1),
		.in_wire_0_2(horizontal_tile_0_1_to_tile_0_0_2),
		.in_wire_0_3(horizontal_tile_0_1_to_tile_0_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_0_0_id_wire)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_2_in_wire_0_3_const_29(
		.out(pe_tile_1_2_in_wire_0_3_const),
		.in(wire_29)
	);

	pe_tile_bottom pe_tile_2_1(
		.out_wire_3_0(vertical_tile_2_1_to_tile_1_1_0),
		.out_wire_3_1(vertical_tile_2_1_to_tile_1_1_1),
		.out_wire_3_2(vertical_tile_2_1_to_tile_1_1_2),
		.out_wire_3_3(vertical_tile_2_1_to_tile_1_1_3),
		.in_wire_3_0(vertical_tile_1_1_to_tile_2_1_0),
		.in_wire_3_1(vertical_tile_1_1_to_tile_2_1_1),
		.in_wire_3_2(vertical_tile_1_1_to_tile_2_1_2),
		.in_wire_3_3(vertical_tile_1_1_to_tile_2_1_3),
		.out_wire_1_0(out_pad_1_pin_to_pe_tile_2_1_out_wire_1_0),
		.in_wire_1_0(pe_tile_2_1_in_wire_1_0_const),
		.in_wire_1_1(pe_tile_2_1_in_wire_1_1_const),
		.in_wire_1_2(pe_tile_2_1_in_wire_1_2_const),
		.in_wire_1_3(pe_tile_2_1_in_wire_1_3_const),
		.out_wire_2_0(horizontal_tile_2_1_to_tile_2_0_0),
		.out_wire_2_1(horizontal_tile_2_1_to_tile_2_0_1),
		.out_wire_2_2(horizontal_tile_2_1_to_tile_2_0_2),
		.out_wire_2_3(horizontal_tile_2_1_to_tile_2_0_3),
		.in_wire_2_0(horizontal_tile_2_0_to_tile_2_1_0),
		.in_wire_2_1(horizontal_tile_2_0_to_tile_2_1_1),
		.in_wire_2_2(horizontal_tile_2_0_to_tile_2_1_2),
		.in_wire_2_3(horizontal_tile_2_0_to_tile_2_1_3),
		.out_wire_0_0(horizontal_tile_2_1_to_tile_2_2_0),
		.out_wire_0_1(horizontal_tile_2_1_to_tile_2_2_1),
		.out_wire_0_2(horizontal_tile_2_1_to_tile_2_2_2),
		.out_wire_0_3(horizontal_tile_2_1_to_tile_2_2_3),
		.in_wire_0_0(horizontal_tile_2_2_to_tile_2_1_0),
		.in_wire_0_1(horizontal_tile_2_2_to_tile_2_1_1),
		.in_wire_0_2(horizontal_tile_2_2_to_tile_2_1_2),
		.in_wire_0_3(horizontal_tile_2_2_to_tile_2_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(pe_tile_2_1_id_wire)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_0in_wire_2_3_const_6_const(
		.out(wire_6)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_2_in_wire_3_2_const_13_const(
		.out(wire_13)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_0in_wire_2_0_const_35_const(
		.out(wire_35)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0_in_wire_3_1_const_0(
		.out(pe_tile_0_0_in_wire_3_1_const),
		.in(wire_0)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_1_in_wire_3_3_const_10_const(
		.out(wire_10)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_0in_wire_2_0_const_3_const(
		.out(wire_3)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_1_0_const_45(
		.out(pe_tile_2_2_in_wire_1_0_const),
		.in(wire_45)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_2_in_wire_0_0_const_15_const(
		.out(wire_15)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_3_3_const_14(
		.out(pe_tile_0_2_in_wire_3_3_const),
		.in(wire_14)
	);

	const_mod #(.width(1), .value(8))  assign_pe_tile_2_1_id_wire_44_const(
		.out(wire_44)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_0_in_wire_3_2_const_1_const(
		.out(wire_1)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_2_in_wire_0_3_const_18_const(
		.out(wire_18)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_3_1_const_12(
		.out(pe_tile_0_2_in_wire_3_1_const),
		.in(wire_12)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_0_in_wire_3_2_const_1(
		.out(pe_tile_0_0_in_wire_3_2_const),
		.in(wire_1)
	);

	const_mod #(.width(1), .value(1))  assign_pe_tile_0_0_id_wire_7_const(
		.out(wire_7)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_2_in_wire_0_2_const_17_const(
		.out(wire_17)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_1_in_wire_1_3_const_43(
		.out(pe_tile_2_1_in_wire_1_3_const),
		.in(wire_43)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_id_wire_53(
		.out(pe_tile_2_2_id_wire),
		.in(wire_53)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_0_3_const_18(
		.out(pe_tile_0_2_in_wire_0_3_const),
		.in(wire_18)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_1_in_wire_3_2_const_9_const(
		.out(wire_9)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_0_1_const_16(
		.out(pe_tile_0_2_in_wire_0_1_const),
		.in(wire_16)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0_id_wire_39(
		.out(pe_tile_2_0_id_wire),
		.in(wire_39)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_0_in_wire_1_3_const_34_const(
		.out(wire_34)
	);

	const_mod #(.width(1), .value(9))  assign_pe_tile_2_2_id_wire_53_const(
		.out(wire_53)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_0_in_wire_1_1_const_32_const(
		.out(wire_32)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0_in_wire_1_3_const_34(
		.out(pe_tile_2_0_in_wire_1_3_const),
		.in(wire_34)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_1_in_wire_1_2_const_42_const(
		.out(wire_42)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_0in_wire_2_1_const_4_const(
		.out(wire_4)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_2_in_wire_0_1_const_27(
		.out(pe_tile_1_2_in_wire_0_1_const),
		.in(wire_27)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_0in_wire_2_3_const_38_const(
		.out(wire_38)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_0_0_const_15(
		.out(pe_tile_0_2_in_wire_0_0_const),
		.in(wire_15)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_1_1_const_46(
		.out(pe_tile_2_2_in_wire_1_1_const),
		.in(wire_46)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_2_1_in_wire_1_3_const_43_const(
		.out(wire_43)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_1_2_in_wire_0_2_const_28_const(
		.out(wire_28)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0_in_wire_1_2_const_33(
		.out(pe_tile_2_0_in_wire_1_2_const),
		.in(wire_33)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_1_2_in_wire_0_0_const_26_const(
		.out(wire_26)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_0in_wire_2_2_const_37(
		.out(pe_tile_2_0in_wire_2_2_const),
		.in(wire_37)
	);

	const_mod #(.width(1), .value(6))  assign_pe_tile_1_2_id_wire_30_const(
		.out(wire_30)
	);

	assign_mod #(.width(1))  assign_pe_tile_0_2_in_wire_3_2_const_13(
		.out(pe_tile_0_2_in_wire_3_2_const),
		.in(wire_13)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_0_2_in_wire_0_1_const_16_const(
		.out(wire_16)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_1_0in_wire_2_1_const_21_const(
		.out(wire_21)
	);

	const_mod #(.width(1), .value(1'b0))  assign_pe_tile_1_2_in_wire_0_1_const_27_const(
		.out(wire_27)
	);

	assign_mod #(.width(1))  assign_pe_tile_2_2_in_wire_0_3_const_52(
		.out(pe_tile_2_2_in_wire_0_3_const),
		.in(wire_52)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_0in_wire_2_3_const_23(
		.out(pe_tile_1_0in_wire_2_3_const),
		.in(wire_23)
	);

	io1in_pad in_pad_2(
		.clk(clk),
		.top_pin(in_wire_2),
		.pin(in_pad_2_pin_to_pe_tile_0_2_in_wire_3_0)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_0_id_wire_24(
		.out(pe_tile_1_0_id_wire),
		.in(wire_24)
	);

	io1in_pad in_pad_0(
		.clk(clk),
		.top_pin(in_wire_0),
		.pin(in_pad_0_pin_to_pe_tile_0_0_in_wire_3_0)
	);

	io1in_pad in_pad_1(
		.clk(clk),
		.top_pin(in_wire_1),
		.pin(in_pad_1_pin_to_pe_tile_0_1_in_wire_3_0)
	);

	assign_mod #(.width(1))  assign_pe_tile_1_2_id_wire_30(
		.out(pe_tile_1_2_id_wire),
		.in(wire_30)
	);



endmodule