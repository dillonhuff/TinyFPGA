module connect_box(input clk,
                   input rst);

   
endmodule
