module pe_tile(input clk,
               input rst);

   
endmodule
