`ifndef pe_tile_included
`define pe_tile_included 1
`include "pe_tile"
`endif
`ifndef io1in_pad_included
`define io1in_pad_included 1
`include "io1in_pad"
`endif
`ifndef io1out_pad_included
`define io1out_pad_included 1
`include "io1out_pad"
`endif


module top(
	input clk,
	input reset,
	input [31:0] config_addr,
	input [31:0] config_data,
	input in_wire_0,
	input in_wire_1,
	input in_wire_2,
	input in_wire_3,
	input in_wire_4,
	input in_wire_5,
	input in_wire_6,
	input in_wire_7,
	input in_wire_8,
	input in_wire_9,
	input in_wire_10,
	input in_wire_11,
	input in_wire_12,
	input in_wire_13,
	input in_wire_14,
	input in_wire_15,
	input in_wire_16,
	input in_wire_17,
	input in_wire_18,
	input in_wire_19,
	input in_wire_20,
	input in_wire_21,
	input in_wire_22,
	input in_wire_23,
	input in_wire_24,
	input in_wire_25,
	input in_wire_26,
	input in_wire_27,
	input in_wire_28,
	input in_wire_29,
	input in_wire_30,
	input in_wire_31,
	output out_wire_0,
	output out_wire_1,
	output out_wire_2,
	output out_wire_3,
	output out_wire_4,
	output out_wire_5,
	output out_wire_6,
	output out_wire_7,
	output out_wire_8,
	output out_wire_9,
	output out_wire_10,
	output out_wire_11,
	output out_wire_12,
	output out_wire_13,
	output out_wire_14,
	output out_wire_15,
	output out_wire_16,
	output out_wire_17,
	output out_wire_18,
	output out_wire_19,
	output out_wire_20,
	output out_wire_21,
	output out_wire_22,
	output out_wire_23,
	output out_wire_24,
	output out_wire_25,
	output out_wire_26,
	output out_wire_27,
	output out_wire_28,
	output out_wire_29,
	output out_wire_30,
	output out_wire_31
	);

	wire input_to_grid_0;
	wire input_to_grid_1;
	wire input_to_grid_2;
	wire input_to_grid_3;
	wire input_to_grid_4;
	wire input_to_grid_5;
	wire input_to_grid_6;
	wire input_to_grid_7;
	wire input_to_grid_8;
	wire input_to_grid_9;
	wire input_to_grid_10;
	wire input_to_grid_11;
	wire input_to_grid_12;
	wire input_to_grid_13;
	wire input_to_grid_14;
	wire input_to_grid_15;
	wire input_to_grid_16;
	wire input_to_grid_17;
	wire input_to_grid_18;
	wire input_to_grid_19;
	wire input_to_grid_20;
	wire input_to_grid_21;
	wire input_to_grid_22;
	wire input_to_grid_23;
	wire input_to_grid_24;
	wire input_to_grid_25;
	wire input_to_grid_26;
	wire input_to_grid_27;
	wire input_to_grid_28;
	wire input_to_grid_29;
	wire input_to_grid_30;
	wire input_to_grid_31;


	wire grid_to_output_0;
	wire grid_to_output_1;
	wire grid_to_output_2;
	wire grid_to_output_3;
	wire grid_to_output_4;
	wire grid_to_output_5;
	wire grid_to_output_6;
	wire grid_to_output_7;
	wire grid_to_output_8;
	wire grid_to_output_9;
	wire grid_to_output_10;
	wire grid_to_output_11;
	wire grid_to_output_12;
	wire grid_to_output_13;
	wire grid_to_output_14;
	wire grid_to_output_15;
	wire grid_to_output_16;
	wire grid_to_output_17;
	wire grid_to_output_18;
	wire grid_to_output_19;
	wire grid_to_output_20;
	wire grid_to_output_21;
	wire grid_to_output_22;
	wire grid_to_output_23;
	wire grid_to_output_24;
	wire grid_to_output_25;
	wire grid_to_output_26;
	wire grid_to_output_27;
	wire grid_to_output_28;
	wire grid_to_output_29;
	wire grid_to_output_30;
	wire grid_to_output_31;


	// input pads
	io1in_pad in_pad_0(
		.clk(clk),
		.top_pin(in_wire_0),
		.pin(input_to_grid_0)
	);

	io1in_pad in_pad_1(
		.clk(clk),
		.top_pin(in_wire_1),
		.pin(input_to_grid_1)
	);

	io1in_pad in_pad_2(
		.clk(clk),
		.top_pin(in_wire_2),
		.pin(input_to_grid_2)
	);

	io1in_pad in_pad_3(
		.clk(clk),
		.top_pin(in_wire_3),
		.pin(input_to_grid_3)
	);

	io1in_pad in_pad_4(
		.clk(clk),
		.top_pin(in_wire_4),
		.pin(input_to_grid_4)
	);

	io1in_pad in_pad_5(
		.clk(clk),
		.top_pin(in_wire_5),
		.pin(input_to_grid_5)
	);

	io1in_pad in_pad_6(
		.clk(clk),
		.top_pin(in_wire_6),
		.pin(input_to_grid_6)
	);

	io1in_pad in_pad_7(
		.clk(clk),
		.top_pin(in_wire_7),
		.pin(input_to_grid_7)
	);

	io1in_pad in_pad_8(
		.clk(clk),
		.top_pin(in_wire_8),
		.pin(input_to_grid_8)
	);

	io1in_pad in_pad_9(
		.clk(clk),
		.top_pin(in_wire_9),
		.pin(input_to_grid_9)
	);

	io1in_pad in_pad_10(
		.clk(clk),
		.top_pin(in_wire_10),
		.pin(input_to_grid_10)
	);

	io1in_pad in_pad_11(
		.clk(clk),
		.top_pin(in_wire_11),
		.pin(input_to_grid_11)
	);

	io1in_pad in_pad_12(
		.clk(clk),
		.top_pin(in_wire_12),
		.pin(input_to_grid_12)
	);

	io1in_pad in_pad_13(
		.clk(clk),
		.top_pin(in_wire_13),
		.pin(input_to_grid_13)
	);

	io1in_pad in_pad_14(
		.clk(clk),
		.top_pin(in_wire_14),
		.pin(input_to_grid_14)
	);

	io1in_pad in_pad_15(
		.clk(clk),
		.top_pin(in_wire_15),
		.pin(input_to_grid_15)
	);

	io1in_pad in_pad_16(
		.clk(clk),
		.top_pin(in_wire_16),
		.pin(input_to_grid_16)
	);

	io1in_pad in_pad_17(
		.clk(clk),
		.top_pin(in_wire_17),
		.pin(input_to_grid_17)
	);

	io1in_pad in_pad_18(
		.clk(clk),
		.top_pin(in_wire_18),
		.pin(input_to_grid_18)
	);

	io1in_pad in_pad_19(
		.clk(clk),
		.top_pin(in_wire_19),
		.pin(input_to_grid_19)
	);

	io1in_pad in_pad_20(
		.clk(clk),
		.top_pin(in_wire_20),
		.pin(input_to_grid_20)
	);

	io1in_pad in_pad_21(
		.clk(clk),
		.top_pin(in_wire_21),
		.pin(input_to_grid_21)
	);

	io1in_pad in_pad_22(
		.clk(clk),
		.top_pin(in_wire_22),
		.pin(input_to_grid_22)
	);

	io1in_pad in_pad_23(
		.clk(clk),
		.top_pin(in_wire_23),
		.pin(input_to_grid_23)
	);

	io1in_pad in_pad_24(
		.clk(clk),
		.top_pin(in_wire_24),
		.pin(input_to_grid_24)
	);

	io1in_pad in_pad_25(
		.clk(clk),
		.top_pin(in_wire_25),
		.pin(input_to_grid_25)
	);

	io1in_pad in_pad_26(
		.clk(clk),
		.top_pin(in_wire_26),
		.pin(input_to_grid_26)
	);

	io1in_pad in_pad_27(
		.clk(clk),
		.top_pin(in_wire_27),
		.pin(input_to_grid_27)
	);

	io1in_pad in_pad_28(
		.clk(clk),
		.top_pin(in_wire_28),
		.pin(input_to_grid_28)
	);

	io1in_pad in_pad_29(
		.clk(clk),
		.top_pin(in_wire_29),
		.pin(input_to_grid_29)
	);

	io1in_pad in_pad_30(
		.clk(clk),
		.top_pin(in_wire_30),
		.pin(input_to_grid_30)
	);

	io1in_pad in_pad_31(
		.clk(clk),
		.top_pin(in_wire_31),
		.pin(input_to_grid_31)
	);

	// output pads
	io1out_pad out_pad_0(
		.clk(clk),
		.top_pin(out_wire_0),
		.pin(grid_to_output_0)
	);

	io1out_pad out_pad_1(
		.clk(clk),
		.top_pin(out_wire_1),
		.pin(grid_to_output_1)
	);

	io1out_pad out_pad_2(
		.clk(clk),
		.top_pin(out_wire_2),
		.pin(grid_to_output_2)
	);

	io1out_pad out_pad_3(
		.clk(clk),
		.top_pin(out_wire_3),
		.pin(grid_to_output_3)
	);

	io1out_pad out_pad_4(
		.clk(clk),
		.top_pin(out_wire_4),
		.pin(grid_to_output_4)
	);

	io1out_pad out_pad_5(
		.clk(clk),
		.top_pin(out_wire_5),
		.pin(grid_to_output_5)
	);

	io1out_pad out_pad_6(
		.clk(clk),
		.top_pin(out_wire_6),
		.pin(grid_to_output_6)
	);

	io1out_pad out_pad_7(
		.clk(clk),
		.top_pin(out_wire_7),
		.pin(grid_to_output_7)
	);

	io1out_pad out_pad_8(
		.clk(clk),
		.top_pin(out_wire_8),
		.pin(grid_to_output_8)
	);

	io1out_pad out_pad_9(
		.clk(clk),
		.top_pin(out_wire_9),
		.pin(grid_to_output_9)
	);

	io1out_pad out_pad_10(
		.clk(clk),
		.top_pin(out_wire_10),
		.pin(grid_to_output_10)
	);

	io1out_pad out_pad_11(
		.clk(clk),
		.top_pin(out_wire_11),
		.pin(grid_to_output_11)
	);

	io1out_pad out_pad_12(
		.clk(clk),
		.top_pin(out_wire_12),
		.pin(grid_to_output_12)
	);

	io1out_pad out_pad_13(
		.clk(clk),
		.top_pin(out_wire_13),
		.pin(grid_to_output_13)
	);

	io1out_pad out_pad_14(
		.clk(clk),
		.top_pin(out_wire_14),
		.pin(grid_to_output_14)
	);

	io1out_pad out_pad_15(
		.clk(clk),
		.top_pin(out_wire_15),
		.pin(grid_to_output_15)
	);

	io1out_pad out_pad_16(
		.clk(clk),
		.top_pin(out_wire_16),
		.pin(grid_to_output_16)
	);

	io1out_pad out_pad_17(
		.clk(clk),
		.top_pin(out_wire_17),
		.pin(grid_to_output_17)
	);

	io1out_pad out_pad_18(
		.clk(clk),
		.top_pin(out_wire_18),
		.pin(grid_to_output_18)
	);

	io1out_pad out_pad_19(
		.clk(clk),
		.top_pin(out_wire_19),
		.pin(grid_to_output_19)
	);

	io1out_pad out_pad_20(
		.clk(clk),
		.top_pin(out_wire_20),
		.pin(grid_to_output_20)
	);

	io1out_pad out_pad_21(
		.clk(clk),
		.top_pin(out_wire_21),
		.pin(grid_to_output_21)
	);

	io1out_pad out_pad_22(
		.clk(clk),
		.top_pin(out_wire_22),
		.pin(grid_to_output_22)
	);

	io1out_pad out_pad_23(
		.clk(clk),
		.top_pin(out_wire_23),
		.pin(grid_to_output_23)
	);

	io1out_pad out_pad_24(
		.clk(clk),
		.top_pin(out_wire_24),
		.pin(grid_to_output_24)
	);

	io1out_pad out_pad_25(
		.clk(clk),
		.top_pin(out_wire_25),
		.pin(grid_to_output_25)
	);

	io1out_pad out_pad_26(
		.clk(clk),
		.top_pin(out_wire_26),
		.pin(grid_to_output_26)
	);

	io1out_pad out_pad_27(
		.clk(clk),
		.top_pin(out_wire_27),
		.pin(grid_to_output_27)
	);

	io1out_pad out_pad_28(
		.clk(clk),
		.top_pin(out_wire_28),
		.pin(grid_to_output_28)
	);

	io1out_pad out_pad_29(
		.clk(clk),
		.top_pin(out_wire_29),
		.pin(grid_to_output_29)
	);

	io1out_pad out_pad_30(
		.clk(clk),
		.top_pin(out_wire_30),
		.pin(grid_to_output_30)
	);

	io1out_pad out_pad_31(
		.clk(clk),
		.top_pin(out_wire_31),
		.pin(grid_to_output_31)
	);

	// PE tile grid
	// Vertical wires
	wire vertical_tile_0_0_to_tile_1_0_0;
	wire vertical_tile_0_0_to_tile_1_0_1;
	wire vertical_tile_0_0_to_tile_1_0_2;
	wire vertical_tile_0_0_to_tile_1_0_3;
	wire vertical_tile_1_0_to_tile_0_0_0;
	wire vertical_tile_1_0_to_tile_0_0_1;
	wire vertical_tile_1_0_to_tile_0_0_2;
	wire vertical_tile_1_0_to_tile_0_0_3;

	wire vertical_tile_0_1_to_tile_1_1_0;
	wire vertical_tile_0_1_to_tile_1_1_1;
	wire vertical_tile_0_1_to_tile_1_1_2;
	wire vertical_tile_0_1_to_tile_1_1_3;
	wire vertical_tile_1_1_to_tile_0_1_0;
	wire vertical_tile_1_1_to_tile_0_1_1;
	wire vertical_tile_1_1_to_tile_0_1_2;
	wire vertical_tile_1_1_to_tile_0_1_3;

	wire vertical_tile_0_2_to_tile_1_2_0;
	wire vertical_tile_0_2_to_tile_1_2_1;
	wire vertical_tile_0_2_to_tile_1_2_2;
	wire vertical_tile_0_2_to_tile_1_2_3;
	wire vertical_tile_1_2_to_tile_0_2_0;
	wire vertical_tile_1_2_to_tile_0_2_1;
	wire vertical_tile_1_2_to_tile_0_2_2;
	wire vertical_tile_1_2_to_tile_0_2_3;

	wire vertical_tile_0_3_to_tile_1_3_0;
	wire vertical_tile_0_3_to_tile_1_3_1;
	wire vertical_tile_0_3_to_tile_1_3_2;
	wire vertical_tile_0_3_to_tile_1_3_3;
	wire vertical_tile_1_3_to_tile_0_3_0;
	wire vertical_tile_1_3_to_tile_0_3_1;
	wire vertical_tile_1_3_to_tile_0_3_2;
	wire vertical_tile_1_3_to_tile_0_3_3;

	wire vertical_tile_0_4_to_tile_1_4_0;
	wire vertical_tile_0_4_to_tile_1_4_1;
	wire vertical_tile_0_4_to_tile_1_4_2;
	wire vertical_tile_0_4_to_tile_1_4_3;
	wire vertical_tile_1_4_to_tile_0_4_0;
	wire vertical_tile_1_4_to_tile_0_4_1;
	wire vertical_tile_1_4_to_tile_0_4_2;
	wire vertical_tile_1_4_to_tile_0_4_3;

	wire vertical_tile_0_5_to_tile_1_5_0;
	wire vertical_tile_0_5_to_tile_1_5_1;
	wire vertical_tile_0_5_to_tile_1_5_2;
	wire vertical_tile_0_5_to_tile_1_5_3;
	wire vertical_tile_1_5_to_tile_0_5_0;
	wire vertical_tile_1_5_to_tile_0_5_1;
	wire vertical_tile_1_5_to_tile_0_5_2;
	wire vertical_tile_1_5_to_tile_0_5_3;

	wire vertical_tile_0_6_to_tile_1_6_0;
	wire vertical_tile_0_6_to_tile_1_6_1;
	wire vertical_tile_0_6_to_tile_1_6_2;
	wire vertical_tile_0_6_to_tile_1_6_3;
	wire vertical_tile_1_6_to_tile_0_6_0;
	wire vertical_tile_1_6_to_tile_0_6_1;
	wire vertical_tile_1_6_to_tile_0_6_2;
	wire vertical_tile_1_6_to_tile_0_6_3;

	wire vertical_tile_0_7_to_tile_1_7_0;
	wire vertical_tile_0_7_to_tile_1_7_1;
	wire vertical_tile_0_7_to_tile_1_7_2;
	wire vertical_tile_0_7_to_tile_1_7_3;
	wire vertical_tile_1_7_to_tile_0_7_0;
	wire vertical_tile_1_7_to_tile_0_7_1;
	wire vertical_tile_1_7_to_tile_0_7_2;
	wire vertical_tile_1_7_to_tile_0_7_3;

	wire vertical_tile_0_8_to_tile_1_8_0;
	wire vertical_tile_0_8_to_tile_1_8_1;
	wire vertical_tile_0_8_to_tile_1_8_2;
	wire vertical_tile_0_8_to_tile_1_8_3;
	wire vertical_tile_1_8_to_tile_0_8_0;
	wire vertical_tile_1_8_to_tile_0_8_1;
	wire vertical_tile_1_8_to_tile_0_8_2;
	wire vertical_tile_1_8_to_tile_0_8_3;

	wire vertical_tile_0_9_to_tile_1_9_0;
	wire vertical_tile_0_9_to_tile_1_9_1;
	wire vertical_tile_0_9_to_tile_1_9_2;
	wire vertical_tile_0_9_to_tile_1_9_3;
	wire vertical_tile_1_9_to_tile_0_9_0;
	wire vertical_tile_1_9_to_tile_0_9_1;
	wire vertical_tile_1_9_to_tile_0_9_2;
	wire vertical_tile_1_9_to_tile_0_9_3;

	wire vertical_tile_0_10_to_tile_1_10_0;
	wire vertical_tile_0_10_to_tile_1_10_1;
	wire vertical_tile_0_10_to_tile_1_10_2;
	wire vertical_tile_0_10_to_tile_1_10_3;
	wire vertical_tile_1_10_to_tile_0_10_0;
	wire vertical_tile_1_10_to_tile_0_10_1;
	wire vertical_tile_1_10_to_tile_0_10_2;
	wire vertical_tile_1_10_to_tile_0_10_3;

	wire vertical_tile_0_11_to_tile_1_11_0;
	wire vertical_tile_0_11_to_tile_1_11_1;
	wire vertical_tile_0_11_to_tile_1_11_2;
	wire vertical_tile_0_11_to_tile_1_11_3;
	wire vertical_tile_1_11_to_tile_0_11_0;
	wire vertical_tile_1_11_to_tile_0_11_1;
	wire vertical_tile_1_11_to_tile_0_11_2;
	wire vertical_tile_1_11_to_tile_0_11_3;

	wire vertical_tile_0_12_to_tile_1_12_0;
	wire vertical_tile_0_12_to_tile_1_12_1;
	wire vertical_tile_0_12_to_tile_1_12_2;
	wire vertical_tile_0_12_to_tile_1_12_3;
	wire vertical_tile_1_12_to_tile_0_12_0;
	wire vertical_tile_1_12_to_tile_0_12_1;
	wire vertical_tile_1_12_to_tile_0_12_2;
	wire vertical_tile_1_12_to_tile_0_12_3;

	wire vertical_tile_0_13_to_tile_1_13_0;
	wire vertical_tile_0_13_to_tile_1_13_1;
	wire vertical_tile_0_13_to_tile_1_13_2;
	wire vertical_tile_0_13_to_tile_1_13_3;
	wire vertical_tile_1_13_to_tile_0_13_0;
	wire vertical_tile_1_13_to_tile_0_13_1;
	wire vertical_tile_1_13_to_tile_0_13_2;
	wire vertical_tile_1_13_to_tile_0_13_3;

	wire vertical_tile_0_14_to_tile_1_14_0;
	wire vertical_tile_0_14_to_tile_1_14_1;
	wire vertical_tile_0_14_to_tile_1_14_2;
	wire vertical_tile_0_14_to_tile_1_14_3;
	wire vertical_tile_1_14_to_tile_0_14_0;
	wire vertical_tile_1_14_to_tile_0_14_1;
	wire vertical_tile_1_14_to_tile_0_14_2;
	wire vertical_tile_1_14_to_tile_0_14_3;

	wire vertical_tile_0_15_to_tile_1_15_0;
	wire vertical_tile_0_15_to_tile_1_15_1;
	wire vertical_tile_0_15_to_tile_1_15_2;
	wire vertical_tile_0_15_to_tile_1_15_3;
	wire vertical_tile_1_15_to_tile_0_15_0;
	wire vertical_tile_1_15_to_tile_0_15_1;
	wire vertical_tile_1_15_to_tile_0_15_2;
	wire vertical_tile_1_15_to_tile_0_15_3;

	wire vertical_tile_0_16_to_tile_1_16_0;
	wire vertical_tile_0_16_to_tile_1_16_1;
	wire vertical_tile_0_16_to_tile_1_16_2;
	wire vertical_tile_0_16_to_tile_1_16_3;
	wire vertical_tile_1_16_to_tile_0_16_0;
	wire vertical_tile_1_16_to_tile_0_16_1;
	wire vertical_tile_1_16_to_tile_0_16_2;
	wire vertical_tile_1_16_to_tile_0_16_3;

	wire vertical_tile_0_17_to_tile_1_17_0;
	wire vertical_tile_0_17_to_tile_1_17_1;
	wire vertical_tile_0_17_to_tile_1_17_2;
	wire vertical_tile_0_17_to_tile_1_17_3;
	wire vertical_tile_1_17_to_tile_0_17_0;
	wire vertical_tile_1_17_to_tile_0_17_1;
	wire vertical_tile_1_17_to_tile_0_17_2;
	wire vertical_tile_1_17_to_tile_0_17_3;

	wire vertical_tile_0_18_to_tile_1_18_0;
	wire vertical_tile_0_18_to_tile_1_18_1;
	wire vertical_tile_0_18_to_tile_1_18_2;
	wire vertical_tile_0_18_to_tile_1_18_3;
	wire vertical_tile_1_18_to_tile_0_18_0;
	wire vertical_tile_1_18_to_tile_0_18_1;
	wire vertical_tile_1_18_to_tile_0_18_2;
	wire vertical_tile_1_18_to_tile_0_18_3;

	wire vertical_tile_0_19_to_tile_1_19_0;
	wire vertical_tile_0_19_to_tile_1_19_1;
	wire vertical_tile_0_19_to_tile_1_19_2;
	wire vertical_tile_0_19_to_tile_1_19_3;
	wire vertical_tile_1_19_to_tile_0_19_0;
	wire vertical_tile_1_19_to_tile_0_19_1;
	wire vertical_tile_1_19_to_tile_0_19_2;
	wire vertical_tile_1_19_to_tile_0_19_3;

	wire vertical_tile_0_20_to_tile_1_20_0;
	wire vertical_tile_0_20_to_tile_1_20_1;
	wire vertical_tile_0_20_to_tile_1_20_2;
	wire vertical_tile_0_20_to_tile_1_20_3;
	wire vertical_tile_1_20_to_tile_0_20_0;
	wire vertical_tile_1_20_to_tile_0_20_1;
	wire vertical_tile_1_20_to_tile_0_20_2;
	wire vertical_tile_1_20_to_tile_0_20_3;

	wire vertical_tile_0_21_to_tile_1_21_0;
	wire vertical_tile_0_21_to_tile_1_21_1;
	wire vertical_tile_0_21_to_tile_1_21_2;
	wire vertical_tile_0_21_to_tile_1_21_3;
	wire vertical_tile_1_21_to_tile_0_21_0;
	wire vertical_tile_1_21_to_tile_0_21_1;
	wire vertical_tile_1_21_to_tile_0_21_2;
	wire vertical_tile_1_21_to_tile_0_21_3;

	wire vertical_tile_0_22_to_tile_1_22_0;
	wire vertical_tile_0_22_to_tile_1_22_1;
	wire vertical_tile_0_22_to_tile_1_22_2;
	wire vertical_tile_0_22_to_tile_1_22_3;
	wire vertical_tile_1_22_to_tile_0_22_0;
	wire vertical_tile_1_22_to_tile_0_22_1;
	wire vertical_tile_1_22_to_tile_0_22_2;
	wire vertical_tile_1_22_to_tile_0_22_3;

	wire vertical_tile_0_23_to_tile_1_23_0;
	wire vertical_tile_0_23_to_tile_1_23_1;
	wire vertical_tile_0_23_to_tile_1_23_2;
	wire vertical_tile_0_23_to_tile_1_23_3;
	wire vertical_tile_1_23_to_tile_0_23_0;
	wire vertical_tile_1_23_to_tile_0_23_1;
	wire vertical_tile_1_23_to_tile_0_23_2;
	wire vertical_tile_1_23_to_tile_0_23_3;

	wire vertical_tile_0_24_to_tile_1_24_0;
	wire vertical_tile_0_24_to_tile_1_24_1;
	wire vertical_tile_0_24_to_tile_1_24_2;
	wire vertical_tile_0_24_to_tile_1_24_3;
	wire vertical_tile_1_24_to_tile_0_24_0;
	wire vertical_tile_1_24_to_tile_0_24_1;
	wire vertical_tile_1_24_to_tile_0_24_2;
	wire vertical_tile_1_24_to_tile_0_24_3;

	wire vertical_tile_0_25_to_tile_1_25_0;
	wire vertical_tile_0_25_to_tile_1_25_1;
	wire vertical_tile_0_25_to_tile_1_25_2;
	wire vertical_tile_0_25_to_tile_1_25_3;
	wire vertical_tile_1_25_to_tile_0_25_0;
	wire vertical_tile_1_25_to_tile_0_25_1;
	wire vertical_tile_1_25_to_tile_0_25_2;
	wire vertical_tile_1_25_to_tile_0_25_3;

	wire vertical_tile_0_26_to_tile_1_26_0;
	wire vertical_tile_0_26_to_tile_1_26_1;
	wire vertical_tile_0_26_to_tile_1_26_2;
	wire vertical_tile_0_26_to_tile_1_26_3;
	wire vertical_tile_1_26_to_tile_0_26_0;
	wire vertical_tile_1_26_to_tile_0_26_1;
	wire vertical_tile_1_26_to_tile_0_26_2;
	wire vertical_tile_1_26_to_tile_0_26_3;

	wire vertical_tile_0_27_to_tile_1_27_0;
	wire vertical_tile_0_27_to_tile_1_27_1;
	wire vertical_tile_0_27_to_tile_1_27_2;
	wire vertical_tile_0_27_to_tile_1_27_3;
	wire vertical_tile_1_27_to_tile_0_27_0;
	wire vertical_tile_1_27_to_tile_0_27_1;
	wire vertical_tile_1_27_to_tile_0_27_2;
	wire vertical_tile_1_27_to_tile_0_27_3;

	wire vertical_tile_0_28_to_tile_1_28_0;
	wire vertical_tile_0_28_to_tile_1_28_1;
	wire vertical_tile_0_28_to_tile_1_28_2;
	wire vertical_tile_0_28_to_tile_1_28_3;
	wire vertical_tile_1_28_to_tile_0_28_0;
	wire vertical_tile_1_28_to_tile_0_28_1;
	wire vertical_tile_1_28_to_tile_0_28_2;
	wire vertical_tile_1_28_to_tile_0_28_3;

	wire vertical_tile_0_29_to_tile_1_29_0;
	wire vertical_tile_0_29_to_tile_1_29_1;
	wire vertical_tile_0_29_to_tile_1_29_2;
	wire vertical_tile_0_29_to_tile_1_29_3;
	wire vertical_tile_1_29_to_tile_0_29_0;
	wire vertical_tile_1_29_to_tile_0_29_1;
	wire vertical_tile_1_29_to_tile_0_29_2;
	wire vertical_tile_1_29_to_tile_0_29_3;

	wire vertical_tile_0_30_to_tile_1_30_0;
	wire vertical_tile_0_30_to_tile_1_30_1;
	wire vertical_tile_0_30_to_tile_1_30_2;
	wire vertical_tile_0_30_to_tile_1_30_3;
	wire vertical_tile_1_30_to_tile_0_30_0;
	wire vertical_tile_1_30_to_tile_0_30_1;
	wire vertical_tile_1_30_to_tile_0_30_2;
	wire vertical_tile_1_30_to_tile_0_30_3;

	wire vertical_tile_0_31_to_tile_1_31_0;
	wire vertical_tile_0_31_to_tile_1_31_1;
	wire vertical_tile_0_31_to_tile_1_31_2;
	wire vertical_tile_0_31_to_tile_1_31_3;
	wire vertical_tile_1_31_to_tile_0_31_0;
	wire vertical_tile_1_31_to_tile_0_31_1;
	wire vertical_tile_1_31_to_tile_0_31_2;
	wire vertical_tile_1_31_to_tile_0_31_3;

	wire vertical_tile_1_0_to_tile_2_0_0;
	wire vertical_tile_1_0_to_tile_2_0_1;
	wire vertical_tile_1_0_to_tile_2_0_2;
	wire vertical_tile_1_0_to_tile_2_0_3;
	wire vertical_tile_2_0_to_tile_1_0_0;
	wire vertical_tile_2_0_to_tile_1_0_1;
	wire vertical_tile_2_0_to_tile_1_0_2;
	wire vertical_tile_2_0_to_tile_1_0_3;

	wire vertical_tile_1_1_to_tile_2_1_0;
	wire vertical_tile_1_1_to_tile_2_1_1;
	wire vertical_tile_1_1_to_tile_2_1_2;
	wire vertical_tile_1_1_to_tile_2_1_3;
	wire vertical_tile_2_1_to_tile_1_1_0;
	wire vertical_tile_2_1_to_tile_1_1_1;
	wire vertical_tile_2_1_to_tile_1_1_2;
	wire vertical_tile_2_1_to_tile_1_1_3;

	wire vertical_tile_1_2_to_tile_2_2_0;
	wire vertical_tile_1_2_to_tile_2_2_1;
	wire vertical_tile_1_2_to_tile_2_2_2;
	wire vertical_tile_1_2_to_tile_2_2_3;
	wire vertical_tile_2_2_to_tile_1_2_0;
	wire vertical_tile_2_2_to_tile_1_2_1;
	wire vertical_tile_2_2_to_tile_1_2_2;
	wire vertical_tile_2_2_to_tile_1_2_3;

	wire vertical_tile_1_3_to_tile_2_3_0;
	wire vertical_tile_1_3_to_tile_2_3_1;
	wire vertical_tile_1_3_to_tile_2_3_2;
	wire vertical_tile_1_3_to_tile_2_3_3;
	wire vertical_tile_2_3_to_tile_1_3_0;
	wire vertical_tile_2_3_to_tile_1_3_1;
	wire vertical_tile_2_3_to_tile_1_3_2;
	wire vertical_tile_2_3_to_tile_1_3_3;

	wire vertical_tile_1_4_to_tile_2_4_0;
	wire vertical_tile_1_4_to_tile_2_4_1;
	wire vertical_tile_1_4_to_tile_2_4_2;
	wire vertical_tile_1_4_to_tile_2_4_3;
	wire vertical_tile_2_4_to_tile_1_4_0;
	wire vertical_tile_2_4_to_tile_1_4_1;
	wire vertical_tile_2_4_to_tile_1_4_2;
	wire vertical_tile_2_4_to_tile_1_4_3;

	wire vertical_tile_1_5_to_tile_2_5_0;
	wire vertical_tile_1_5_to_tile_2_5_1;
	wire vertical_tile_1_5_to_tile_2_5_2;
	wire vertical_tile_1_5_to_tile_2_5_3;
	wire vertical_tile_2_5_to_tile_1_5_0;
	wire vertical_tile_2_5_to_tile_1_5_1;
	wire vertical_tile_2_5_to_tile_1_5_2;
	wire vertical_tile_2_5_to_tile_1_5_3;

	wire vertical_tile_1_6_to_tile_2_6_0;
	wire vertical_tile_1_6_to_tile_2_6_1;
	wire vertical_tile_1_6_to_tile_2_6_2;
	wire vertical_tile_1_6_to_tile_2_6_3;
	wire vertical_tile_2_6_to_tile_1_6_0;
	wire vertical_tile_2_6_to_tile_1_6_1;
	wire vertical_tile_2_6_to_tile_1_6_2;
	wire vertical_tile_2_6_to_tile_1_6_3;

	wire vertical_tile_1_7_to_tile_2_7_0;
	wire vertical_tile_1_7_to_tile_2_7_1;
	wire vertical_tile_1_7_to_tile_2_7_2;
	wire vertical_tile_1_7_to_tile_2_7_3;
	wire vertical_tile_2_7_to_tile_1_7_0;
	wire vertical_tile_2_7_to_tile_1_7_1;
	wire vertical_tile_2_7_to_tile_1_7_2;
	wire vertical_tile_2_7_to_tile_1_7_3;

	wire vertical_tile_1_8_to_tile_2_8_0;
	wire vertical_tile_1_8_to_tile_2_8_1;
	wire vertical_tile_1_8_to_tile_2_8_2;
	wire vertical_tile_1_8_to_tile_2_8_3;
	wire vertical_tile_2_8_to_tile_1_8_0;
	wire vertical_tile_2_8_to_tile_1_8_1;
	wire vertical_tile_2_8_to_tile_1_8_2;
	wire vertical_tile_2_8_to_tile_1_8_3;

	wire vertical_tile_1_9_to_tile_2_9_0;
	wire vertical_tile_1_9_to_tile_2_9_1;
	wire vertical_tile_1_9_to_tile_2_9_2;
	wire vertical_tile_1_9_to_tile_2_9_3;
	wire vertical_tile_2_9_to_tile_1_9_0;
	wire vertical_tile_2_9_to_tile_1_9_1;
	wire vertical_tile_2_9_to_tile_1_9_2;
	wire vertical_tile_2_9_to_tile_1_9_3;

	wire vertical_tile_1_10_to_tile_2_10_0;
	wire vertical_tile_1_10_to_tile_2_10_1;
	wire vertical_tile_1_10_to_tile_2_10_2;
	wire vertical_tile_1_10_to_tile_2_10_3;
	wire vertical_tile_2_10_to_tile_1_10_0;
	wire vertical_tile_2_10_to_tile_1_10_1;
	wire vertical_tile_2_10_to_tile_1_10_2;
	wire vertical_tile_2_10_to_tile_1_10_3;

	wire vertical_tile_1_11_to_tile_2_11_0;
	wire vertical_tile_1_11_to_tile_2_11_1;
	wire vertical_tile_1_11_to_tile_2_11_2;
	wire vertical_tile_1_11_to_tile_2_11_3;
	wire vertical_tile_2_11_to_tile_1_11_0;
	wire vertical_tile_2_11_to_tile_1_11_1;
	wire vertical_tile_2_11_to_tile_1_11_2;
	wire vertical_tile_2_11_to_tile_1_11_3;

	wire vertical_tile_1_12_to_tile_2_12_0;
	wire vertical_tile_1_12_to_tile_2_12_1;
	wire vertical_tile_1_12_to_tile_2_12_2;
	wire vertical_tile_1_12_to_tile_2_12_3;
	wire vertical_tile_2_12_to_tile_1_12_0;
	wire vertical_tile_2_12_to_tile_1_12_1;
	wire vertical_tile_2_12_to_tile_1_12_2;
	wire vertical_tile_2_12_to_tile_1_12_3;

	wire vertical_tile_1_13_to_tile_2_13_0;
	wire vertical_tile_1_13_to_tile_2_13_1;
	wire vertical_tile_1_13_to_tile_2_13_2;
	wire vertical_tile_1_13_to_tile_2_13_3;
	wire vertical_tile_2_13_to_tile_1_13_0;
	wire vertical_tile_2_13_to_tile_1_13_1;
	wire vertical_tile_2_13_to_tile_1_13_2;
	wire vertical_tile_2_13_to_tile_1_13_3;

	wire vertical_tile_1_14_to_tile_2_14_0;
	wire vertical_tile_1_14_to_tile_2_14_1;
	wire vertical_tile_1_14_to_tile_2_14_2;
	wire vertical_tile_1_14_to_tile_2_14_3;
	wire vertical_tile_2_14_to_tile_1_14_0;
	wire vertical_tile_2_14_to_tile_1_14_1;
	wire vertical_tile_2_14_to_tile_1_14_2;
	wire vertical_tile_2_14_to_tile_1_14_3;

	wire vertical_tile_1_15_to_tile_2_15_0;
	wire vertical_tile_1_15_to_tile_2_15_1;
	wire vertical_tile_1_15_to_tile_2_15_2;
	wire vertical_tile_1_15_to_tile_2_15_3;
	wire vertical_tile_2_15_to_tile_1_15_0;
	wire vertical_tile_2_15_to_tile_1_15_1;
	wire vertical_tile_2_15_to_tile_1_15_2;
	wire vertical_tile_2_15_to_tile_1_15_3;

	wire vertical_tile_1_16_to_tile_2_16_0;
	wire vertical_tile_1_16_to_tile_2_16_1;
	wire vertical_tile_1_16_to_tile_2_16_2;
	wire vertical_tile_1_16_to_tile_2_16_3;
	wire vertical_tile_2_16_to_tile_1_16_0;
	wire vertical_tile_2_16_to_tile_1_16_1;
	wire vertical_tile_2_16_to_tile_1_16_2;
	wire vertical_tile_2_16_to_tile_1_16_3;

	wire vertical_tile_1_17_to_tile_2_17_0;
	wire vertical_tile_1_17_to_tile_2_17_1;
	wire vertical_tile_1_17_to_tile_2_17_2;
	wire vertical_tile_1_17_to_tile_2_17_3;
	wire vertical_tile_2_17_to_tile_1_17_0;
	wire vertical_tile_2_17_to_tile_1_17_1;
	wire vertical_tile_2_17_to_tile_1_17_2;
	wire vertical_tile_2_17_to_tile_1_17_3;

	wire vertical_tile_1_18_to_tile_2_18_0;
	wire vertical_tile_1_18_to_tile_2_18_1;
	wire vertical_tile_1_18_to_tile_2_18_2;
	wire vertical_tile_1_18_to_tile_2_18_3;
	wire vertical_tile_2_18_to_tile_1_18_0;
	wire vertical_tile_2_18_to_tile_1_18_1;
	wire vertical_tile_2_18_to_tile_1_18_2;
	wire vertical_tile_2_18_to_tile_1_18_3;

	wire vertical_tile_1_19_to_tile_2_19_0;
	wire vertical_tile_1_19_to_tile_2_19_1;
	wire vertical_tile_1_19_to_tile_2_19_2;
	wire vertical_tile_1_19_to_tile_2_19_3;
	wire vertical_tile_2_19_to_tile_1_19_0;
	wire vertical_tile_2_19_to_tile_1_19_1;
	wire vertical_tile_2_19_to_tile_1_19_2;
	wire vertical_tile_2_19_to_tile_1_19_3;

	wire vertical_tile_1_20_to_tile_2_20_0;
	wire vertical_tile_1_20_to_tile_2_20_1;
	wire vertical_tile_1_20_to_tile_2_20_2;
	wire vertical_tile_1_20_to_tile_2_20_3;
	wire vertical_tile_2_20_to_tile_1_20_0;
	wire vertical_tile_2_20_to_tile_1_20_1;
	wire vertical_tile_2_20_to_tile_1_20_2;
	wire vertical_tile_2_20_to_tile_1_20_3;

	wire vertical_tile_1_21_to_tile_2_21_0;
	wire vertical_tile_1_21_to_tile_2_21_1;
	wire vertical_tile_1_21_to_tile_2_21_2;
	wire vertical_tile_1_21_to_tile_2_21_3;
	wire vertical_tile_2_21_to_tile_1_21_0;
	wire vertical_tile_2_21_to_tile_1_21_1;
	wire vertical_tile_2_21_to_tile_1_21_2;
	wire vertical_tile_2_21_to_tile_1_21_3;

	wire vertical_tile_1_22_to_tile_2_22_0;
	wire vertical_tile_1_22_to_tile_2_22_1;
	wire vertical_tile_1_22_to_tile_2_22_2;
	wire vertical_tile_1_22_to_tile_2_22_3;
	wire vertical_tile_2_22_to_tile_1_22_0;
	wire vertical_tile_2_22_to_tile_1_22_1;
	wire vertical_tile_2_22_to_tile_1_22_2;
	wire vertical_tile_2_22_to_tile_1_22_3;

	wire vertical_tile_1_23_to_tile_2_23_0;
	wire vertical_tile_1_23_to_tile_2_23_1;
	wire vertical_tile_1_23_to_tile_2_23_2;
	wire vertical_tile_1_23_to_tile_2_23_3;
	wire vertical_tile_2_23_to_tile_1_23_0;
	wire vertical_tile_2_23_to_tile_1_23_1;
	wire vertical_tile_2_23_to_tile_1_23_2;
	wire vertical_tile_2_23_to_tile_1_23_3;

	wire vertical_tile_1_24_to_tile_2_24_0;
	wire vertical_tile_1_24_to_tile_2_24_1;
	wire vertical_tile_1_24_to_tile_2_24_2;
	wire vertical_tile_1_24_to_tile_2_24_3;
	wire vertical_tile_2_24_to_tile_1_24_0;
	wire vertical_tile_2_24_to_tile_1_24_1;
	wire vertical_tile_2_24_to_tile_1_24_2;
	wire vertical_tile_2_24_to_tile_1_24_3;

	wire vertical_tile_1_25_to_tile_2_25_0;
	wire vertical_tile_1_25_to_tile_2_25_1;
	wire vertical_tile_1_25_to_tile_2_25_2;
	wire vertical_tile_1_25_to_tile_2_25_3;
	wire vertical_tile_2_25_to_tile_1_25_0;
	wire vertical_tile_2_25_to_tile_1_25_1;
	wire vertical_tile_2_25_to_tile_1_25_2;
	wire vertical_tile_2_25_to_tile_1_25_3;

	wire vertical_tile_1_26_to_tile_2_26_0;
	wire vertical_tile_1_26_to_tile_2_26_1;
	wire vertical_tile_1_26_to_tile_2_26_2;
	wire vertical_tile_1_26_to_tile_2_26_3;
	wire vertical_tile_2_26_to_tile_1_26_0;
	wire vertical_tile_2_26_to_tile_1_26_1;
	wire vertical_tile_2_26_to_tile_1_26_2;
	wire vertical_tile_2_26_to_tile_1_26_3;

	wire vertical_tile_1_27_to_tile_2_27_0;
	wire vertical_tile_1_27_to_tile_2_27_1;
	wire vertical_tile_1_27_to_tile_2_27_2;
	wire vertical_tile_1_27_to_tile_2_27_3;
	wire vertical_tile_2_27_to_tile_1_27_0;
	wire vertical_tile_2_27_to_tile_1_27_1;
	wire vertical_tile_2_27_to_tile_1_27_2;
	wire vertical_tile_2_27_to_tile_1_27_3;

	wire vertical_tile_1_28_to_tile_2_28_0;
	wire vertical_tile_1_28_to_tile_2_28_1;
	wire vertical_tile_1_28_to_tile_2_28_2;
	wire vertical_tile_1_28_to_tile_2_28_3;
	wire vertical_tile_2_28_to_tile_1_28_0;
	wire vertical_tile_2_28_to_tile_1_28_1;
	wire vertical_tile_2_28_to_tile_1_28_2;
	wire vertical_tile_2_28_to_tile_1_28_3;

	wire vertical_tile_1_29_to_tile_2_29_0;
	wire vertical_tile_1_29_to_tile_2_29_1;
	wire vertical_tile_1_29_to_tile_2_29_2;
	wire vertical_tile_1_29_to_tile_2_29_3;
	wire vertical_tile_2_29_to_tile_1_29_0;
	wire vertical_tile_2_29_to_tile_1_29_1;
	wire vertical_tile_2_29_to_tile_1_29_2;
	wire vertical_tile_2_29_to_tile_1_29_3;

	wire vertical_tile_1_30_to_tile_2_30_0;
	wire vertical_tile_1_30_to_tile_2_30_1;
	wire vertical_tile_1_30_to_tile_2_30_2;
	wire vertical_tile_1_30_to_tile_2_30_3;
	wire vertical_tile_2_30_to_tile_1_30_0;
	wire vertical_tile_2_30_to_tile_1_30_1;
	wire vertical_tile_2_30_to_tile_1_30_2;
	wire vertical_tile_2_30_to_tile_1_30_3;

	wire vertical_tile_1_31_to_tile_2_31_0;
	wire vertical_tile_1_31_to_tile_2_31_1;
	wire vertical_tile_1_31_to_tile_2_31_2;
	wire vertical_tile_1_31_to_tile_2_31_3;
	wire vertical_tile_2_31_to_tile_1_31_0;
	wire vertical_tile_2_31_to_tile_1_31_1;
	wire vertical_tile_2_31_to_tile_1_31_2;
	wire vertical_tile_2_31_to_tile_1_31_3;

	wire vertical_tile_2_0_to_tile_3_0_0;
	wire vertical_tile_2_0_to_tile_3_0_1;
	wire vertical_tile_2_0_to_tile_3_0_2;
	wire vertical_tile_2_0_to_tile_3_0_3;
	wire vertical_tile_3_0_to_tile_2_0_0;
	wire vertical_tile_3_0_to_tile_2_0_1;
	wire vertical_tile_3_0_to_tile_2_0_2;
	wire vertical_tile_3_0_to_tile_2_0_3;

	wire vertical_tile_2_1_to_tile_3_1_0;
	wire vertical_tile_2_1_to_tile_3_1_1;
	wire vertical_tile_2_1_to_tile_3_1_2;
	wire vertical_tile_2_1_to_tile_3_1_3;
	wire vertical_tile_3_1_to_tile_2_1_0;
	wire vertical_tile_3_1_to_tile_2_1_1;
	wire vertical_tile_3_1_to_tile_2_1_2;
	wire vertical_tile_3_1_to_tile_2_1_3;

	wire vertical_tile_2_2_to_tile_3_2_0;
	wire vertical_tile_2_2_to_tile_3_2_1;
	wire vertical_tile_2_2_to_tile_3_2_2;
	wire vertical_tile_2_2_to_tile_3_2_3;
	wire vertical_tile_3_2_to_tile_2_2_0;
	wire vertical_tile_3_2_to_tile_2_2_1;
	wire vertical_tile_3_2_to_tile_2_2_2;
	wire vertical_tile_3_2_to_tile_2_2_3;

	wire vertical_tile_2_3_to_tile_3_3_0;
	wire vertical_tile_2_3_to_tile_3_3_1;
	wire vertical_tile_2_3_to_tile_3_3_2;
	wire vertical_tile_2_3_to_tile_3_3_3;
	wire vertical_tile_3_3_to_tile_2_3_0;
	wire vertical_tile_3_3_to_tile_2_3_1;
	wire vertical_tile_3_3_to_tile_2_3_2;
	wire vertical_tile_3_3_to_tile_2_3_3;

	wire vertical_tile_2_4_to_tile_3_4_0;
	wire vertical_tile_2_4_to_tile_3_4_1;
	wire vertical_tile_2_4_to_tile_3_4_2;
	wire vertical_tile_2_4_to_tile_3_4_3;
	wire vertical_tile_3_4_to_tile_2_4_0;
	wire vertical_tile_3_4_to_tile_2_4_1;
	wire vertical_tile_3_4_to_tile_2_4_2;
	wire vertical_tile_3_4_to_tile_2_4_3;

	wire vertical_tile_2_5_to_tile_3_5_0;
	wire vertical_tile_2_5_to_tile_3_5_1;
	wire vertical_tile_2_5_to_tile_3_5_2;
	wire vertical_tile_2_5_to_tile_3_5_3;
	wire vertical_tile_3_5_to_tile_2_5_0;
	wire vertical_tile_3_5_to_tile_2_5_1;
	wire vertical_tile_3_5_to_tile_2_5_2;
	wire vertical_tile_3_5_to_tile_2_5_3;

	wire vertical_tile_2_6_to_tile_3_6_0;
	wire vertical_tile_2_6_to_tile_3_6_1;
	wire vertical_tile_2_6_to_tile_3_6_2;
	wire vertical_tile_2_6_to_tile_3_6_3;
	wire vertical_tile_3_6_to_tile_2_6_0;
	wire vertical_tile_3_6_to_tile_2_6_1;
	wire vertical_tile_3_6_to_tile_2_6_2;
	wire vertical_tile_3_6_to_tile_2_6_3;

	wire vertical_tile_2_7_to_tile_3_7_0;
	wire vertical_tile_2_7_to_tile_3_7_1;
	wire vertical_tile_2_7_to_tile_3_7_2;
	wire vertical_tile_2_7_to_tile_3_7_3;
	wire vertical_tile_3_7_to_tile_2_7_0;
	wire vertical_tile_3_7_to_tile_2_7_1;
	wire vertical_tile_3_7_to_tile_2_7_2;
	wire vertical_tile_3_7_to_tile_2_7_3;

	wire vertical_tile_2_8_to_tile_3_8_0;
	wire vertical_tile_2_8_to_tile_3_8_1;
	wire vertical_tile_2_8_to_tile_3_8_2;
	wire vertical_tile_2_8_to_tile_3_8_3;
	wire vertical_tile_3_8_to_tile_2_8_0;
	wire vertical_tile_3_8_to_tile_2_8_1;
	wire vertical_tile_3_8_to_tile_2_8_2;
	wire vertical_tile_3_8_to_tile_2_8_3;

	wire vertical_tile_2_9_to_tile_3_9_0;
	wire vertical_tile_2_9_to_tile_3_9_1;
	wire vertical_tile_2_9_to_tile_3_9_2;
	wire vertical_tile_2_9_to_tile_3_9_3;
	wire vertical_tile_3_9_to_tile_2_9_0;
	wire vertical_tile_3_9_to_tile_2_9_1;
	wire vertical_tile_3_9_to_tile_2_9_2;
	wire vertical_tile_3_9_to_tile_2_9_3;

	wire vertical_tile_2_10_to_tile_3_10_0;
	wire vertical_tile_2_10_to_tile_3_10_1;
	wire vertical_tile_2_10_to_tile_3_10_2;
	wire vertical_tile_2_10_to_tile_3_10_3;
	wire vertical_tile_3_10_to_tile_2_10_0;
	wire vertical_tile_3_10_to_tile_2_10_1;
	wire vertical_tile_3_10_to_tile_2_10_2;
	wire vertical_tile_3_10_to_tile_2_10_3;

	wire vertical_tile_2_11_to_tile_3_11_0;
	wire vertical_tile_2_11_to_tile_3_11_1;
	wire vertical_tile_2_11_to_tile_3_11_2;
	wire vertical_tile_2_11_to_tile_3_11_3;
	wire vertical_tile_3_11_to_tile_2_11_0;
	wire vertical_tile_3_11_to_tile_2_11_1;
	wire vertical_tile_3_11_to_tile_2_11_2;
	wire vertical_tile_3_11_to_tile_2_11_3;

	wire vertical_tile_2_12_to_tile_3_12_0;
	wire vertical_tile_2_12_to_tile_3_12_1;
	wire vertical_tile_2_12_to_tile_3_12_2;
	wire vertical_tile_2_12_to_tile_3_12_3;
	wire vertical_tile_3_12_to_tile_2_12_0;
	wire vertical_tile_3_12_to_tile_2_12_1;
	wire vertical_tile_3_12_to_tile_2_12_2;
	wire vertical_tile_3_12_to_tile_2_12_3;

	wire vertical_tile_2_13_to_tile_3_13_0;
	wire vertical_tile_2_13_to_tile_3_13_1;
	wire vertical_tile_2_13_to_tile_3_13_2;
	wire vertical_tile_2_13_to_tile_3_13_3;
	wire vertical_tile_3_13_to_tile_2_13_0;
	wire vertical_tile_3_13_to_tile_2_13_1;
	wire vertical_tile_3_13_to_tile_2_13_2;
	wire vertical_tile_3_13_to_tile_2_13_3;

	wire vertical_tile_2_14_to_tile_3_14_0;
	wire vertical_tile_2_14_to_tile_3_14_1;
	wire vertical_tile_2_14_to_tile_3_14_2;
	wire vertical_tile_2_14_to_tile_3_14_3;
	wire vertical_tile_3_14_to_tile_2_14_0;
	wire vertical_tile_3_14_to_tile_2_14_1;
	wire vertical_tile_3_14_to_tile_2_14_2;
	wire vertical_tile_3_14_to_tile_2_14_3;

	wire vertical_tile_2_15_to_tile_3_15_0;
	wire vertical_tile_2_15_to_tile_3_15_1;
	wire vertical_tile_2_15_to_tile_3_15_2;
	wire vertical_tile_2_15_to_tile_3_15_3;
	wire vertical_tile_3_15_to_tile_2_15_0;
	wire vertical_tile_3_15_to_tile_2_15_1;
	wire vertical_tile_3_15_to_tile_2_15_2;
	wire vertical_tile_3_15_to_tile_2_15_3;

	wire vertical_tile_2_16_to_tile_3_16_0;
	wire vertical_tile_2_16_to_tile_3_16_1;
	wire vertical_tile_2_16_to_tile_3_16_2;
	wire vertical_tile_2_16_to_tile_3_16_3;
	wire vertical_tile_3_16_to_tile_2_16_0;
	wire vertical_tile_3_16_to_tile_2_16_1;
	wire vertical_tile_3_16_to_tile_2_16_2;
	wire vertical_tile_3_16_to_tile_2_16_3;

	wire vertical_tile_2_17_to_tile_3_17_0;
	wire vertical_tile_2_17_to_tile_3_17_1;
	wire vertical_tile_2_17_to_tile_3_17_2;
	wire vertical_tile_2_17_to_tile_3_17_3;
	wire vertical_tile_3_17_to_tile_2_17_0;
	wire vertical_tile_3_17_to_tile_2_17_1;
	wire vertical_tile_3_17_to_tile_2_17_2;
	wire vertical_tile_3_17_to_tile_2_17_3;

	wire vertical_tile_2_18_to_tile_3_18_0;
	wire vertical_tile_2_18_to_tile_3_18_1;
	wire vertical_tile_2_18_to_tile_3_18_2;
	wire vertical_tile_2_18_to_tile_3_18_3;
	wire vertical_tile_3_18_to_tile_2_18_0;
	wire vertical_tile_3_18_to_tile_2_18_1;
	wire vertical_tile_3_18_to_tile_2_18_2;
	wire vertical_tile_3_18_to_tile_2_18_3;

	wire vertical_tile_2_19_to_tile_3_19_0;
	wire vertical_tile_2_19_to_tile_3_19_1;
	wire vertical_tile_2_19_to_tile_3_19_2;
	wire vertical_tile_2_19_to_tile_3_19_3;
	wire vertical_tile_3_19_to_tile_2_19_0;
	wire vertical_tile_3_19_to_tile_2_19_1;
	wire vertical_tile_3_19_to_tile_2_19_2;
	wire vertical_tile_3_19_to_tile_2_19_3;

	wire vertical_tile_2_20_to_tile_3_20_0;
	wire vertical_tile_2_20_to_tile_3_20_1;
	wire vertical_tile_2_20_to_tile_3_20_2;
	wire vertical_tile_2_20_to_tile_3_20_3;
	wire vertical_tile_3_20_to_tile_2_20_0;
	wire vertical_tile_3_20_to_tile_2_20_1;
	wire vertical_tile_3_20_to_tile_2_20_2;
	wire vertical_tile_3_20_to_tile_2_20_3;

	wire vertical_tile_2_21_to_tile_3_21_0;
	wire vertical_tile_2_21_to_tile_3_21_1;
	wire vertical_tile_2_21_to_tile_3_21_2;
	wire vertical_tile_2_21_to_tile_3_21_3;
	wire vertical_tile_3_21_to_tile_2_21_0;
	wire vertical_tile_3_21_to_tile_2_21_1;
	wire vertical_tile_3_21_to_tile_2_21_2;
	wire vertical_tile_3_21_to_tile_2_21_3;

	wire vertical_tile_2_22_to_tile_3_22_0;
	wire vertical_tile_2_22_to_tile_3_22_1;
	wire vertical_tile_2_22_to_tile_3_22_2;
	wire vertical_tile_2_22_to_tile_3_22_3;
	wire vertical_tile_3_22_to_tile_2_22_0;
	wire vertical_tile_3_22_to_tile_2_22_1;
	wire vertical_tile_3_22_to_tile_2_22_2;
	wire vertical_tile_3_22_to_tile_2_22_3;

	wire vertical_tile_2_23_to_tile_3_23_0;
	wire vertical_tile_2_23_to_tile_3_23_1;
	wire vertical_tile_2_23_to_tile_3_23_2;
	wire vertical_tile_2_23_to_tile_3_23_3;
	wire vertical_tile_3_23_to_tile_2_23_0;
	wire vertical_tile_3_23_to_tile_2_23_1;
	wire vertical_tile_3_23_to_tile_2_23_2;
	wire vertical_tile_3_23_to_tile_2_23_3;

	wire vertical_tile_2_24_to_tile_3_24_0;
	wire vertical_tile_2_24_to_tile_3_24_1;
	wire vertical_tile_2_24_to_tile_3_24_2;
	wire vertical_tile_2_24_to_tile_3_24_3;
	wire vertical_tile_3_24_to_tile_2_24_0;
	wire vertical_tile_3_24_to_tile_2_24_1;
	wire vertical_tile_3_24_to_tile_2_24_2;
	wire vertical_tile_3_24_to_tile_2_24_3;

	wire vertical_tile_2_25_to_tile_3_25_0;
	wire vertical_tile_2_25_to_tile_3_25_1;
	wire vertical_tile_2_25_to_tile_3_25_2;
	wire vertical_tile_2_25_to_tile_3_25_3;
	wire vertical_tile_3_25_to_tile_2_25_0;
	wire vertical_tile_3_25_to_tile_2_25_1;
	wire vertical_tile_3_25_to_tile_2_25_2;
	wire vertical_tile_3_25_to_tile_2_25_3;

	wire vertical_tile_2_26_to_tile_3_26_0;
	wire vertical_tile_2_26_to_tile_3_26_1;
	wire vertical_tile_2_26_to_tile_3_26_2;
	wire vertical_tile_2_26_to_tile_3_26_3;
	wire vertical_tile_3_26_to_tile_2_26_0;
	wire vertical_tile_3_26_to_tile_2_26_1;
	wire vertical_tile_3_26_to_tile_2_26_2;
	wire vertical_tile_3_26_to_tile_2_26_3;

	wire vertical_tile_2_27_to_tile_3_27_0;
	wire vertical_tile_2_27_to_tile_3_27_1;
	wire vertical_tile_2_27_to_tile_3_27_2;
	wire vertical_tile_2_27_to_tile_3_27_3;
	wire vertical_tile_3_27_to_tile_2_27_0;
	wire vertical_tile_3_27_to_tile_2_27_1;
	wire vertical_tile_3_27_to_tile_2_27_2;
	wire vertical_tile_3_27_to_tile_2_27_3;

	wire vertical_tile_2_28_to_tile_3_28_0;
	wire vertical_tile_2_28_to_tile_3_28_1;
	wire vertical_tile_2_28_to_tile_3_28_2;
	wire vertical_tile_2_28_to_tile_3_28_3;
	wire vertical_tile_3_28_to_tile_2_28_0;
	wire vertical_tile_3_28_to_tile_2_28_1;
	wire vertical_tile_3_28_to_tile_2_28_2;
	wire vertical_tile_3_28_to_tile_2_28_3;

	wire vertical_tile_2_29_to_tile_3_29_0;
	wire vertical_tile_2_29_to_tile_3_29_1;
	wire vertical_tile_2_29_to_tile_3_29_2;
	wire vertical_tile_2_29_to_tile_3_29_3;
	wire vertical_tile_3_29_to_tile_2_29_0;
	wire vertical_tile_3_29_to_tile_2_29_1;
	wire vertical_tile_3_29_to_tile_2_29_2;
	wire vertical_tile_3_29_to_tile_2_29_3;

	wire vertical_tile_2_30_to_tile_3_30_0;
	wire vertical_tile_2_30_to_tile_3_30_1;
	wire vertical_tile_2_30_to_tile_3_30_2;
	wire vertical_tile_2_30_to_tile_3_30_3;
	wire vertical_tile_3_30_to_tile_2_30_0;
	wire vertical_tile_3_30_to_tile_2_30_1;
	wire vertical_tile_3_30_to_tile_2_30_2;
	wire vertical_tile_3_30_to_tile_2_30_3;

	wire vertical_tile_2_31_to_tile_3_31_0;
	wire vertical_tile_2_31_to_tile_3_31_1;
	wire vertical_tile_2_31_to_tile_3_31_2;
	wire vertical_tile_2_31_to_tile_3_31_3;
	wire vertical_tile_3_31_to_tile_2_31_0;
	wire vertical_tile_3_31_to_tile_2_31_1;
	wire vertical_tile_3_31_to_tile_2_31_2;
	wire vertical_tile_3_31_to_tile_2_31_3;

	wire vertical_tile_3_0_to_tile_4_0_0;
	wire vertical_tile_3_0_to_tile_4_0_1;
	wire vertical_tile_3_0_to_tile_4_0_2;
	wire vertical_tile_3_0_to_tile_4_0_3;
	wire vertical_tile_4_0_to_tile_3_0_0;
	wire vertical_tile_4_0_to_tile_3_0_1;
	wire vertical_tile_4_0_to_tile_3_0_2;
	wire vertical_tile_4_0_to_tile_3_0_3;

	wire vertical_tile_3_1_to_tile_4_1_0;
	wire vertical_tile_3_1_to_tile_4_1_1;
	wire vertical_tile_3_1_to_tile_4_1_2;
	wire vertical_tile_3_1_to_tile_4_1_3;
	wire vertical_tile_4_1_to_tile_3_1_0;
	wire vertical_tile_4_1_to_tile_3_1_1;
	wire vertical_tile_4_1_to_tile_3_1_2;
	wire vertical_tile_4_1_to_tile_3_1_3;

	wire vertical_tile_3_2_to_tile_4_2_0;
	wire vertical_tile_3_2_to_tile_4_2_1;
	wire vertical_tile_3_2_to_tile_4_2_2;
	wire vertical_tile_3_2_to_tile_4_2_3;
	wire vertical_tile_4_2_to_tile_3_2_0;
	wire vertical_tile_4_2_to_tile_3_2_1;
	wire vertical_tile_4_2_to_tile_3_2_2;
	wire vertical_tile_4_2_to_tile_3_2_3;

	wire vertical_tile_3_3_to_tile_4_3_0;
	wire vertical_tile_3_3_to_tile_4_3_1;
	wire vertical_tile_3_3_to_tile_4_3_2;
	wire vertical_tile_3_3_to_tile_4_3_3;
	wire vertical_tile_4_3_to_tile_3_3_0;
	wire vertical_tile_4_3_to_tile_3_3_1;
	wire vertical_tile_4_3_to_tile_3_3_2;
	wire vertical_tile_4_3_to_tile_3_3_3;

	wire vertical_tile_3_4_to_tile_4_4_0;
	wire vertical_tile_3_4_to_tile_4_4_1;
	wire vertical_tile_3_4_to_tile_4_4_2;
	wire vertical_tile_3_4_to_tile_4_4_3;
	wire vertical_tile_4_4_to_tile_3_4_0;
	wire vertical_tile_4_4_to_tile_3_4_1;
	wire vertical_tile_4_4_to_tile_3_4_2;
	wire vertical_tile_4_4_to_tile_3_4_3;

	wire vertical_tile_3_5_to_tile_4_5_0;
	wire vertical_tile_3_5_to_tile_4_5_1;
	wire vertical_tile_3_5_to_tile_4_5_2;
	wire vertical_tile_3_5_to_tile_4_5_3;
	wire vertical_tile_4_5_to_tile_3_5_0;
	wire vertical_tile_4_5_to_tile_3_5_1;
	wire vertical_tile_4_5_to_tile_3_5_2;
	wire vertical_tile_4_5_to_tile_3_5_3;

	wire vertical_tile_3_6_to_tile_4_6_0;
	wire vertical_tile_3_6_to_tile_4_6_1;
	wire vertical_tile_3_6_to_tile_4_6_2;
	wire vertical_tile_3_6_to_tile_4_6_3;
	wire vertical_tile_4_6_to_tile_3_6_0;
	wire vertical_tile_4_6_to_tile_3_6_1;
	wire vertical_tile_4_6_to_tile_3_6_2;
	wire vertical_tile_4_6_to_tile_3_6_3;

	wire vertical_tile_3_7_to_tile_4_7_0;
	wire vertical_tile_3_7_to_tile_4_7_1;
	wire vertical_tile_3_7_to_tile_4_7_2;
	wire vertical_tile_3_7_to_tile_4_7_3;
	wire vertical_tile_4_7_to_tile_3_7_0;
	wire vertical_tile_4_7_to_tile_3_7_1;
	wire vertical_tile_4_7_to_tile_3_7_2;
	wire vertical_tile_4_7_to_tile_3_7_3;

	wire vertical_tile_3_8_to_tile_4_8_0;
	wire vertical_tile_3_8_to_tile_4_8_1;
	wire vertical_tile_3_8_to_tile_4_8_2;
	wire vertical_tile_3_8_to_tile_4_8_3;
	wire vertical_tile_4_8_to_tile_3_8_0;
	wire vertical_tile_4_8_to_tile_3_8_1;
	wire vertical_tile_4_8_to_tile_3_8_2;
	wire vertical_tile_4_8_to_tile_3_8_3;

	wire vertical_tile_3_9_to_tile_4_9_0;
	wire vertical_tile_3_9_to_tile_4_9_1;
	wire vertical_tile_3_9_to_tile_4_9_2;
	wire vertical_tile_3_9_to_tile_4_9_3;
	wire vertical_tile_4_9_to_tile_3_9_0;
	wire vertical_tile_4_9_to_tile_3_9_1;
	wire vertical_tile_4_9_to_tile_3_9_2;
	wire vertical_tile_4_9_to_tile_3_9_3;

	wire vertical_tile_3_10_to_tile_4_10_0;
	wire vertical_tile_3_10_to_tile_4_10_1;
	wire vertical_tile_3_10_to_tile_4_10_2;
	wire vertical_tile_3_10_to_tile_4_10_3;
	wire vertical_tile_4_10_to_tile_3_10_0;
	wire vertical_tile_4_10_to_tile_3_10_1;
	wire vertical_tile_4_10_to_tile_3_10_2;
	wire vertical_tile_4_10_to_tile_3_10_3;

	wire vertical_tile_3_11_to_tile_4_11_0;
	wire vertical_tile_3_11_to_tile_4_11_1;
	wire vertical_tile_3_11_to_tile_4_11_2;
	wire vertical_tile_3_11_to_tile_4_11_3;
	wire vertical_tile_4_11_to_tile_3_11_0;
	wire vertical_tile_4_11_to_tile_3_11_1;
	wire vertical_tile_4_11_to_tile_3_11_2;
	wire vertical_tile_4_11_to_tile_3_11_3;

	wire vertical_tile_3_12_to_tile_4_12_0;
	wire vertical_tile_3_12_to_tile_4_12_1;
	wire vertical_tile_3_12_to_tile_4_12_2;
	wire vertical_tile_3_12_to_tile_4_12_3;
	wire vertical_tile_4_12_to_tile_3_12_0;
	wire vertical_tile_4_12_to_tile_3_12_1;
	wire vertical_tile_4_12_to_tile_3_12_2;
	wire vertical_tile_4_12_to_tile_3_12_3;

	wire vertical_tile_3_13_to_tile_4_13_0;
	wire vertical_tile_3_13_to_tile_4_13_1;
	wire vertical_tile_3_13_to_tile_4_13_2;
	wire vertical_tile_3_13_to_tile_4_13_3;
	wire vertical_tile_4_13_to_tile_3_13_0;
	wire vertical_tile_4_13_to_tile_3_13_1;
	wire vertical_tile_4_13_to_tile_3_13_2;
	wire vertical_tile_4_13_to_tile_3_13_3;

	wire vertical_tile_3_14_to_tile_4_14_0;
	wire vertical_tile_3_14_to_tile_4_14_1;
	wire vertical_tile_3_14_to_tile_4_14_2;
	wire vertical_tile_3_14_to_tile_4_14_3;
	wire vertical_tile_4_14_to_tile_3_14_0;
	wire vertical_tile_4_14_to_tile_3_14_1;
	wire vertical_tile_4_14_to_tile_3_14_2;
	wire vertical_tile_4_14_to_tile_3_14_3;

	wire vertical_tile_3_15_to_tile_4_15_0;
	wire vertical_tile_3_15_to_tile_4_15_1;
	wire vertical_tile_3_15_to_tile_4_15_2;
	wire vertical_tile_3_15_to_tile_4_15_3;
	wire vertical_tile_4_15_to_tile_3_15_0;
	wire vertical_tile_4_15_to_tile_3_15_1;
	wire vertical_tile_4_15_to_tile_3_15_2;
	wire vertical_tile_4_15_to_tile_3_15_3;

	wire vertical_tile_3_16_to_tile_4_16_0;
	wire vertical_tile_3_16_to_tile_4_16_1;
	wire vertical_tile_3_16_to_tile_4_16_2;
	wire vertical_tile_3_16_to_tile_4_16_3;
	wire vertical_tile_4_16_to_tile_3_16_0;
	wire vertical_tile_4_16_to_tile_3_16_1;
	wire vertical_tile_4_16_to_tile_3_16_2;
	wire vertical_tile_4_16_to_tile_3_16_3;

	wire vertical_tile_3_17_to_tile_4_17_0;
	wire vertical_tile_3_17_to_tile_4_17_1;
	wire vertical_tile_3_17_to_tile_4_17_2;
	wire vertical_tile_3_17_to_tile_4_17_3;
	wire vertical_tile_4_17_to_tile_3_17_0;
	wire vertical_tile_4_17_to_tile_3_17_1;
	wire vertical_tile_4_17_to_tile_3_17_2;
	wire vertical_tile_4_17_to_tile_3_17_3;

	wire vertical_tile_3_18_to_tile_4_18_0;
	wire vertical_tile_3_18_to_tile_4_18_1;
	wire vertical_tile_3_18_to_tile_4_18_2;
	wire vertical_tile_3_18_to_tile_4_18_3;
	wire vertical_tile_4_18_to_tile_3_18_0;
	wire vertical_tile_4_18_to_tile_3_18_1;
	wire vertical_tile_4_18_to_tile_3_18_2;
	wire vertical_tile_4_18_to_tile_3_18_3;

	wire vertical_tile_3_19_to_tile_4_19_0;
	wire vertical_tile_3_19_to_tile_4_19_1;
	wire vertical_tile_3_19_to_tile_4_19_2;
	wire vertical_tile_3_19_to_tile_4_19_3;
	wire vertical_tile_4_19_to_tile_3_19_0;
	wire vertical_tile_4_19_to_tile_3_19_1;
	wire vertical_tile_4_19_to_tile_3_19_2;
	wire vertical_tile_4_19_to_tile_3_19_3;

	wire vertical_tile_3_20_to_tile_4_20_0;
	wire vertical_tile_3_20_to_tile_4_20_1;
	wire vertical_tile_3_20_to_tile_4_20_2;
	wire vertical_tile_3_20_to_tile_4_20_3;
	wire vertical_tile_4_20_to_tile_3_20_0;
	wire vertical_tile_4_20_to_tile_3_20_1;
	wire vertical_tile_4_20_to_tile_3_20_2;
	wire vertical_tile_4_20_to_tile_3_20_3;

	wire vertical_tile_3_21_to_tile_4_21_0;
	wire vertical_tile_3_21_to_tile_4_21_1;
	wire vertical_tile_3_21_to_tile_4_21_2;
	wire vertical_tile_3_21_to_tile_4_21_3;
	wire vertical_tile_4_21_to_tile_3_21_0;
	wire vertical_tile_4_21_to_tile_3_21_1;
	wire vertical_tile_4_21_to_tile_3_21_2;
	wire vertical_tile_4_21_to_tile_3_21_3;

	wire vertical_tile_3_22_to_tile_4_22_0;
	wire vertical_tile_3_22_to_tile_4_22_1;
	wire vertical_tile_3_22_to_tile_4_22_2;
	wire vertical_tile_3_22_to_tile_4_22_3;
	wire vertical_tile_4_22_to_tile_3_22_0;
	wire vertical_tile_4_22_to_tile_3_22_1;
	wire vertical_tile_4_22_to_tile_3_22_2;
	wire vertical_tile_4_22_to_tile_3_22_3;

	wire vertical_tile_3_23_to_tile_4_23_0;
	wire vertical_tile_3_23_to_tile_4_23_1;
	wire vertical_tile_3_23_to_tile_4_23_2;
	wire vertical_tile_3_23_to_tile_4_23_3;
	wire vertical_tile_4_23_to_tile_3_23_0;
	wire vertical_tile_4_23_to_tile_3_23_1;
	wire vertical_tile_4_23_to_tile_3_23_2;
	wire vertical_tile_4_23_to_tile_3_23_3;

	wire vertical_tile_3_24_to_tile_4_24_0;
	wire vertical_tile_3_24_to_tile_4_24_1;
	wire vertical_tile_3_24_to_tile_4_24_2;
	wire vertical_tile_3_24_to_tile_4_24_3;
	wire vertical_tile_4_24_to_tile_3_24_0;
	wire vertical_tile_4_24_to_tile_3_24_1;
	wire vertical_tile_4_24_to_tile_3_24_2;
	wire vertical_tile_4_24_to_tile_3_24_3;

	wire vertical_tile_3_25_to_tile_4_25_0;
	wire vertical_tile_3_25_to_tile_4_25_1;
	wire vertical_tile_3_25_to_tile_4_25_2;
	wire vertical_tile_3_25_to_tile_4_25_3;
	wire vertical_tile_4_25_to_tile_3_25_0;
	wire vertical_tile_4_25_to_tile_3_25_1;
	wire vertical_tile_4_25_to_tile_3_25_2;
	wire vertical_tile_4_25_to_tile_3_25_3;

	wire vertical_tile_3_26_to_tile_4_26_0;
	wire vertical_tile_3_26_to_tile_4_26_1;
	wire vertical_tile_3_26_to_tile_4_26_2;
	wire vertical_tile_3_26_to_tile_4_26_3;
	wire vertical_tile_4_26_to_tile_3_26_0;
	wire vertical_tile_4_26_to_tile_3_26_1;
	wire vertical_tile_4_26_to_tile_3_26_2;
	wire vertical_tile_4_26_to_tile_3_26_3;

	wire vertical_tile_3_27_to_tile_4_27_0;
	wire vertical_tile_3_27_to_tile_4_27_1;
	wire vertical_tile_3_27_to_tile_4_27_2;
	wire vertical_tile_3_27_to_tile_4_27_3;
	wire vertical_tile_4_27_to_tile_3_27_0;
	wire vertical_tile_4_27_to_tile_3_27_1;
	wire vertical_tile_4_27_to_tile_3_27_2;
	wire vertical_tile_4_27_to_tile_3_27_3;

	wire vertical_tile_3_28_to_tile_4_28_0;
	wire vertical_tile_3_28_to_tile_4_28_1;
	wire vertical_tile_3_28_to_tile_4_28_2;
	wire vertical_tile_3_28_to_tile_4_28_3;
	wire vertical_tile_4_28_to_tile_3_28_0;
	wire vertical_tile_4_28_to_tile_3_28_1;
	wire vertical_tile_4_28_to_tile_3_28_2;
	wire vertical_tile_4_28_to_tile_3_28_3;

	wire vertical_tile_3_29_to_tile_4_29_0;
	wire vertical_tile_3_29_to_tile_4_29_1;
	wire vertical_tile_3_29_to_tile_4_29_2;
	wire vertical_tile_3_29_to_tile_4_29_3;
	wire vertical_tile_4_29_to_tile_3_29_0;
	wire vertical_tile_4_29_to_tile_3_29_1;
	wire vertical_tile_4_29_to_tile_3_29_2;
	wire vertical_tile_4_29_to_tile_3_29_3;

	wire vertical_tile_3_30_to_tile_4_30_0;
	wire vertical_tile_3_30_to_tile_4_30_1;
	wire vertical_tile_3_30_to_tile_4_30_2;
	wire vertical_tile_3_30_to_tile_4_30_3;
	wire vertical_tile_4_30_to_tile_3_30_0;
	wire vertical_tile_4_30_to_tile_3_30_1;
	wire vertical_tile_4_30_to_tile_3_30_2;
	wire vertical_tile_4_30_to_tile_3_30_3;

	wire vertical_tile_3_31_to_tile_4_31_0;
	wire vertical_tile_3_31_to_tile_4_31_1;
	wire vertical_tile_3_31_to_tile_4_31_2;
	wire vertical_tile_3_31_to_tile_4_31_3;
	wire vertical_tile_4_31_to_tile_3_31_0;
	wire vertical_tile_4_31_to_tile_3_31_1;
	wire vertical_tile_4_31_to_tile_3_31_2;
	wire vertical_tile_4_31_to_tile_3_31_3;

	wire vertical_tile_4_0_to_tile_5_0_0;
	wire vertical_tile_4_0_to_tile_5_0_1;
	wire vertical_tile_4_0_to_tile_5_0_2;
	wire vertical_tile_4_0_to_tile_5_0_3;
	wire vertical_tile_5_0_to_tile_4_0_0;
	wire vertical_tile_5_0_to_tile_4_0_1;
	wire vertical_tile_5_0_to_tile_4_0_2;
	wire vertical_tile_5_0_to_tile_4_0_3;

	wire vertical_tile_4_1_to_tile_5_1_0;
	wire vertical_tile_4_1_to_tile_5_1_1;
	wire vertical_tile_4_1_to_tile_5_1_2;
	wire vertical_tile_4_1_to_tile_5_1_3;
	wire vertical_tile_5_1_to_tile_4_1_0;
	wire vertical_tile_5_1_to_tile_4_1_1;
	wire vertical_tile_5_1_to_tile_4_1_2;
	wire vertical_tile_5_1_to_tile_4_1_3;

	wire vertical_tile_4_2_to_tile_5_2_0;
	wire vertical_tile_4_2_to_tile_5_2_1;
	wire vertical_tile_4_2_to_tile_5_2_2;
	wire vertical_tile_4_2_to_tile_5_2_3;
	wire vertical_tile_5_2_to_tile_4_2_0;
	wire vertical_tile_5_2_to_tile_4_2_1;
	wire vertical_tile_5_2_to_tile_4_2_2;
	wire vertical_tile_5_2_to_tile_4_2_3;

	wire vertical_tile_4_3_to_tile_5_3_0;
	wire vertical_tile_4_3_to_tile_5_3_1;
	wire vertical_tile_4_3_to_tile_5_3_2;
	wire vertical_tile_4_3_to_tile_5_3_3;
	wire vertical_tile_5_3_to_tile_4_3_0;
	wire vertical_tile_5_3_to_tile_4_3_1;
	wire vertical_tile_5_3_to_tile_4_3_2;
	wire vertical_tile_5_3_to_tile_4_3_3;

	wire vertical_tile_4_4_to_tile_5_4_0;
	wire vertical_tile_4_4_to_tile_5_4_1;
	wire vertical_tile_4_4_to_tile_5_4_2;
	wire vertical_tile_4_4_to_tile_5_4_3;
	wire vertical_tile_5_4_to_tile_4_4_0;
	wire vertical_tile_5_4_to_tile_4_4_1;
	wire vertical_tile_5_4_to_tile_4_4_2;
	wire vertical_tile_5_4_to_tile_4_4_3;

	wire vertical_tile_4_5_to_tile_5_5_0;
	wire vertical_tile_4_5_to_tile_5_5_1;
	wire vertical_tile_4_5_to_tile_5_5_2;
	wire vertical_tile_4_5_to_tile_5_5_3;
	wire vertical_tile_5_5_to_tile_4_5_0;
	wire vertical_tile_5_5_to_tile_4_5_1;
	wire vertical_tile_5_5_to_tile_4_5_2;
	wire vertical_tile_5_5_to_tile_4_5_3;

	wire vertical_tile_4_6_to_tile_5_6_0;
	wire vertical_tile_4_6_to_tile_5_6_1;
	wire vertical_tile_4_6_to_tile_5_6_2;
	wire vertical_tile_4_6_to_tile_5_6_3;
	wire vertical_tile_5_6_to_tile_4_6_0;
	wire vertical_tile_5_6_to_tile_4_6_1;
	wire vertical_tile_5_6_to_tile_4_6_2;
	wire vertical_tile_5_6_to_tile_4_6_3;

	wire vertical_tile_4_7_to_tile_5_7_0;
	wire vertical_tile_4_7_to_tile_5_7_1;
	wire vertical_tile_4_7_to_tile_5_7_2;
	wire vertical_tile_4_7_to_tile_5_7_3;
	wire vertical_tile_5_7_to_tile_4_7_0;
	wire vertical_tile_5_7_to_tile_4_7_1;
	wire vertical_tile_5_7_to_tile_4_7_2;
	wire vertical_tile_5_7_to_tile_4_7_3;

	wire vertical_tile_4_8_to_tile_5_8_0;
	wire vertical_tile_4_8_to_tile_5_8_1;
	wire vertical_tile_4_8_to_tile_5_8_2;
	wire vertical_tile_4_8_to_tile_5_8_3;
	wire vertical_tile_5_8_to_tile_4_8_0;
	wire vertical_tile_5_8_to_tile_4_8_1;
	wire vertical_tile_5_8_to_tile_4_8_2;
	wire vertical_tile_5_8_to_tile_4_8_3;

	wire vertical_tile_4_9_to_tile_5_9_0;
	wire vertical_tile_4_9_to_tile_5_9_1;
	wire vertical_tile_4_9_to_tile_5_9_2;
	wire vertical_tile_4_9_to_tile_5_9_3;
	wire vertical_tile_5_9_to_tile_4_9_0;
	wire vertical_tile_5_9_to_tile_4_9_1;
	wire vertical_tile_5_9_to_tile_4_9_2;
	wire vertical_tile_5_9_to_tile_4_9_3;

	wire vertical_tile_4_10_to_tile_5_10_0;
	wire vertical_tile_4_10_to_tile_5_10_1;
	wire vertical_tile_4_10_to_tile_5_10_2;
	wire vertical_tile_4_10_to_tile_5_10_3;
	wire vertical_tile_5_10_to_tile_4_10_0;
	wire vertical_tile_5_10_to_tile_4_10_1;
	wire vertical_tile_5_10_to_tile_4_10_2;
	wire vertical_tile_5_10_to_tile_4_10_3;

	wire vertical_tile_4_11_to_tile_5_11_0;
	wire vertical_tile_4_11_to_tile_5_11_1;
	wire vertical_tile_4_11_to_tile_5_11_2;
	wire vertical_tile_4_11_to_tile_5_11_3;
	wire vertical_tile_5_11_to_tile_4_11_0;
	wire vertical_tile_5_11_to_tile_4_11_1;
	wire vertical_tile_5_11_to_tile_4_11_2;
	wire vertical_tile_5_11_to_tile_4_11_3;

	wire vertical_tile_4_12_to_tile_5_12_0;
	wire vertical_tile_4_12_to_tile_5_12_1;
	wire vertical_tile_4_12_to_tile_5_12_2;
	wire vertical_tile_4_12_to_tile_5_12_3;
	wire vertical_tile_5_12_to_tile_4_12_0;
	wire vertical_tile_5_12_to_tile_4_12_1;
	wire vertical_tile_5_12_to_tile_4_12_2;
	wire vertical_tile_5_12_to_tile_4_12_3;

	wire vertical_tile_4_13_to_tile_5_13_0;
	wire vertical_tile_4_13_to_tile_5_13_1;
	wire vertical_tile_4_13_to_tile_5_13_2;
	wire vertical_tile_4_13_to_tile_5_13_3;
	wire vertical_tile_5_13_to_tile_4_13_0;
	wire vertical_tile_5_13_to_tile_4_13_1;
	wire vertical_tile_5_13_to_tile_4_13_2;
	wire vertical_tile_5_13_to_tile_4_13_3;

	wire vertical_tile_4_14_to_tile_5_14_0;
	wire vertical_tile_4_14_to_tile_5_14_1;
	wire vertical_tile_4_14_to_tile_5_14_2;
	wire vertical_tile_4_14_to_tile_5_14_3;
	wire vertical_tile_5_14_to_tile_4_14_0;
	wire vertical_tile_5_14_to_tile_4_14_1;
	wire vertical_tile_5_14_to_tile_4_14_2;
	wire vertical_tile_5_14_to_tile_4_14_3;

	wire vertical_tile_4_15_to_tile_5_15_0;
	wire vertical_tile_4_15_to_tile_5_15_1;
	wire vertical_tile_4_15_to_tile_5_15_2;
	wire vertical_tile_4_15_to_tile_5_15_3;
	wire vertical_tile_5_15_to_tile_4_15_0;
	wire vertical_tile_5_15_to_tile_4_15_1;
	wire vertical_tile_5_15_to_tile_4_15_2;
	wire vertical_tile_5_15_to_tile_4_15_3;

	wire vertical_tile_4_16_to_tile_5_16_0;
	wire vertical_tile_4_16_to_tile_5_16_1;
	wire vertical_tile_4_16_to_tile_5_16_2;
	wire vertical_tile_4_16_to_tile_5_16_3;
	wire vertical_tile_5_16_to_tile_4_16_0;
	wire vertical_tile_5_16_to_tile_4_16_1;
	wire vertical_tile_5_16_to_tile_4_16_2;
	wire vertical_tile_5_16_to_tile_4_16_3;

	wire vertical_tile_4_17_to_tile_5_17_0;
	wire vertical_tile_4_17_to_tile_5_17_1;
	wire vertical_tile_4_17_to_tile_5_17_2;
	wire vertical_tile_4_17_to_tile_5_17_3;
	wire vertical_tile_5_17_to_tile_4_17_0;
	wire vertical_tile_5_17_to_tile_4_17_1;
	wire vertical_tile_5_17_to_tile_4_17_2;
	wire vertical_tile_5_17_to_tile_4_17_3;

	wire vertical_tile_4_18_to_tile_5_18_0;
	wire vertical_tile_4_18_to_tile_5_18_1;
	wire vertical_tile_4_18_to_tile_5_18_2;
	wire vertical_tile_4_18_to_tile_5_18_3;
	wire vertical_tile_5_18_to_tile_4_18_0;
	wire vertical_tile_5_18_to_tile_4_18_1;
	wire vertical_tile_5_18_to_tile_4_18_2;
	wire vertical_tile_5_18_to_tile_4_18_3;

	wire vertical_tile_4_19_to_tile_5_19_0;
	wire vertical_tile_4_19_to_tile_5_19_1;
	wire vertical_tile_4_19_to_tile_5_19_2;
	wire vertical_tile_4_19_to_tile_5_19_3;
	wire vertical_tile_5_19_to_tile_4_19_0;
	wire vertical_tile_5_19_to_tile_4_19_1;
	wire vertical_tile_5_19_to_tile_4_19_2;
	wire vertical_tile_5_19_to_tile_4_19_3;

	wire vertical_tile_4_20_to_tile_5_20_0;
	wire vertical_tile_4_20_to_tile_5_20_1;
	wire vertical_tile_4_20_to_tile_5_20_2;
	wire vertical_tile_4_20_to_tile_5_20_3;
	wire vertical_tile_5_20_to_tile_4_20_0;
	wire vertical_tile_5_20_to_tile_4_20_1;
	wire vertical_tile_5_20_to_tile_4_20_2;
	wire vertical_tile_5_20_to_tile_4_20_3;

	wire vertical_tile_4_21_to_tile_5_21_0;
	wire vertical_tile_4_21_to_tile_5_21_1;
	wire vertical_tile_4_21_to_tile_5_21_2;
	wire vertical_tile_4_21_to_tile_5_21_3;
	wire vertical_tile_5_21_to_tile_4_21_0;
	wire vertical_tile_5_21_to_tile_4_21_1;
	wire vertical_tile_5_21_to_tile_4_21_2;
	wire vertical_tile_5_21_to_tile_4_21_3;

	wire vertical_tile_4_22_to_tile_5_22_0;
	wire vertical_tile_4_22_to_tile_5_22_1;
	wire vertical_tile_4_22_to_tile_5_22_2;
	wire vertical_tile_4_22_to_tile_5_22_3;
	wire vertical_tile_5_22_to_tile_4_22_0;
	wire vertical_tile_5_22_to_tile_4_22_1;
	wire vertical_tile_5_22_to_tile_4_22_2;
	wire vertical_tile_5_22_to_tile_4_22_3;

	wire vertical_tile_4_23_to_tile_5_23_0;
	wire vertical_tile_4_23_to_tile_5_23_1;
	wire vertical_tile_4_23_to_tile_5_23_2;
	wire vertical_tile_4_23_to_tile_5_23_3;
	wire vertical_tile_5_23_to_tile_4_23_0;
	wire vertical_tile_5_23_to_tile_4_23_1;
	wire vertical_tile_5_23_to_tile_4_23_2;
	wire vertical_tile_5_23_to_tile_4_23_3;

	wire vertical_tile_4_24_to_tile_5_24_0;
	wire vertical_tile_4_24_to_tile_5_24_1;
	wire vertical_tile_4_24_to_tile_5_24_2;
	wire vertical_tile_4_24_to_tile_5_24_3;
	wire vertical_tile_5_24_to_tile_4_24_0;
	wire vertical_tile_5_24_to_tile_4_24_1;
	wire vertical_tile_5_24_to_tile_4_24_2;
	wire vertical_tile_5_24_to_tile_4_24_3;

	wire vertical_tile_4_25_to_tile_5_25_0;
	wire vertical_tile_4_25_to_tile_5_25_1;
	wire vertical_tile_4_25_to_tile_5_25_2;
	wire vertical_tile_4_25_to_tile_5_25_3;
	wire vertical_tile_5_25_to_tile_4_25_0;
	wire vertical_tile_5_25_to_tile_4_25_1;
	wire vertical_tile_5_25_to_tile_4_25_2;
	wire vertical_tile_5_25_to_tile_4_25_3;

	wire vertical_tile_4_26_to_tile_5_26_0;
	wire vertical_tile_4_26_to_tile_5_26_1;
	wire vertical_tile_4_26_to_tile_5_26_2;
	wire vertical_tile_4_26_to_tile_5_26_3;
	wire vertical_tile_5_26_to_tile_4_26_0;
	wire vertical_tile_5_26_to_tile_4_26_1;
	wire vertical_tile_5_26_to_tile_4_26_2;
	wire vertical_tile_5_26_to_tile_4_26_3;

	wire vertical_tile_4_27_to_tile_5_27_0;
	wire vertical_tile_4_27_to_tile_5_27_1;
	wire vertical_tile_4_27_to_tile_5_27_2;
	wire vertical_tile_4_27_to_tile_5_27_3;
	wire vertical_tile_5_27_to_tile_4_27_0;
	wire vertical_tile_5_27_to_tile_4_27_1;
	wire vertical_tile_5_27_to_tile_4_27_2;
	wire vertical_tile_5_27_to_tile_4_27_3;

	wire vertical_tile_4_28_to_tile_5_28_0;
	wire vertical_tile_4_28_to_tile_5_28_1;
	wire vertical_tile_4_28_to_tile_5_28_2;
	wire vertical_tile_4_28_to_tile_5_28_3;
	wire vertical_tile_5_28_to_tile_4_28_0;
	wire vertical_tile_5_28_to_tile_4_28_1;
	wire vertical_tile_5_28_to_tile_4_28_2;
	wire vertical_tile_5_28_to_tile_4_28_3;

	wire vertical_tile_4_29_to_tile_5_29_0;
	wire vertical_tile_4_29_to_tile_5_29_1;
	wire vertical_tile_4_29_to_tile_5_29_2;
	wire vertical_tile_4_29_to_tile_5_29_3;
	wire vertical_tile_5_29_to_tile_4_29_0;
	wire vertical_tile_5_29_to_tile_4_29_1;
	wire vertical_tile_5_29_to_tile_4_29_2;
	wire vertical_tile_5_29_to_tile_4_29_3;

	wire vertical_tile_4_30_to_tile_5_30_0;
	wire vertical_tile_4_30_to_tile_5_30_1;
	wire vertical_tile_4_30_to_tile_5_30_2;
	wire vertical_tile_4_30_to_tile_5_30_3;
	wire vertical_tile_5_30_to_tile_4_30_0;
	wire vertical_tile_5_30_to_tile_4_30_1;
	wire vertical_tile_5_30_to_tile_4_30_2;
	wire vertical_tile_5_30_to_tile_4_30_3;

	wire vertical_tile_4_31_to_tile_5_31_0;
	wire vertical_tile_4_31_to_tile_5_31_1;
	wire vertical_tile_4_31_to_tile_5_31_2;
	wire vertical_tile_4_31_to_tile_5_31_3;
	wire vertical_tile_5_31_to_tile_4_31_0;
	wire vertical_tile_5_31_to_tile_4_31_1;
	wire vertical_tile_5_31_to_tile_4_31_2;
	wire vertical_tile_5_31_to_tile_4_31_3;

	wire vertical_tile_5_0_to_tile_6_0_0;
	wire vertical_tile_5_0_to_tile_6_0_1;
	wire vertical_tile_5_0_to_tile_6_0_2;
	wire vertical_tile_5_0_to_tile_6_0_3;
	wire vertical_tile_6_0_to_tile_5_0_0;
	wire vertical_tile_6_0_to_tile_5_0_1;
	wire vertical_tile_6_0_to_tile_5_0_2;
	wire vertical_tile_6_0_to_tile_5_0_3;

	wire vertical_tile_5_1_to_tile_6_1_0;
	wire vertical_tile_5_1_to_tile_6_1_1;
	wire vertical_tile_5_1_to_tile_6_1_2;
	wire vertical_tile_5_1_to_tile_6_1_3;
	wire vertical_tile_6_1_to_tile_5_1_0;
	wire vertical_tile_6_1_to_tile_5_1_1;
	wire vertical_tile_6_1_to_tile_5_1_2;
	wire vertical_tile_6_1_to_tile_5_1_3;

	wire vertical_tile_5_2_to_tile_6_2_0;
	wire vertical_tile_5_2_to_tile_6_2_1;
	wire vertical_tile_5_2_to_tile_6_2_2;
	wire vertical_tile_5_2_to_tile_6_2_3;
	wire vertical_tile_6_2_to_tile_5_2_0;
	wire vertical_tile_6_2_to_tile_5_2_1;
	wire vertical_tile_6_2_to_tile_5_2_2;
	wire vertical_tile_6_2_to_tile_5_2_3;

	wire vertical_tile_5_3_to_tile_6_3_0;
	wire vertical_tile_5_3_to_tile_6_3_1;
	wire vertical_tile_5_3_to_tile_6_3_2;
	wire vertical_tile_5_3_to_tile_6_3_3;
	wire vertical_tile_6_3_to_tile_5_3_0;
	wire vertical_tile_6_3_to_tile_5_3_1;
	wire vertical_tile_6_3_to_tile_5_3_2;
	wire vertical_tile_6_3_to_tile_5_3_3;

	wire vertical_tile_5_4_to_tile_6_4_0;
	wire vertical_tile_5_4_to_tile_6_4_1;
	wire vertical_tile_5_4_to_tile_6_4_2;
	wire vertical_tile_5_4_to_tile_6_4_3;
	wire vertical_tile_6_4_to_tile_5_4_0;
	wire vertical_tile_6_4_to_tile_5_4_1;
	wire vertical_tile_6_4_to_tile_5_4_2;
	wire vertical_tile_6_4_to_tile_5_4_3;

	wire vertical_tile_5_5_to_tile_6_5_0;
	wire vertical_tile_5_5_to_tile_6_5_1;
	wire vertical_tile_5_5_to_tile_6_5_2;
	wire vertical_tile_5_5_to_tile_6_5_3;
	wire vertical_tile_6_5_to_tile_5_5_0;
	wire vertical_tile_6_5_to_tile_5_5_1;
	wire vertical_tile_6_5_to_tile_5_5_2;
	wire vertical_tile_6_5_to_tile_5_5_3;

	wire vertical_tile_5_6_to_tile_6_6_0;
	wire vertical_tile_5_6_to_tile_6_6_1;
	wire vertical_tile_5_6_to_tile_6_6_2;
	wire vertical_tile_5_6_to_tile_6_6_3;
	wire vertical_tile_6_6_to_tile_5_6_0;
	wire vertical_tile_6_6_to_tile_5_6_1;
	wire vertical_tile_6_6_to_tile_5_6_2;
	wire vertical_tile_6_6_to_tile_5_6_3;

	wire vertical_tile_5_7_to_tile_6_7_0;
	wire vertical_tile_5_7_to_tile_6_7_1;
	wire vertical_tile_5_7_to_tile_6_7_2;
	wire vertical_tile_5_7_to_tile_6_7_3;
	wire vertical_tile_6_7_to_tile_5_7_0;
	wire vertical_tile_6_7_to_tile_5_7_1;
	wire vertical_tile_6_7_to_tile_5_7_2;
	wire vertical_tile_6_7_to_tile_5_7_3;

	wire vertical_tile_5_8_to_tile_6_8_0;
	wire vertical_tile_5_8_to_tile_6_8_1;
	wire vertical_tile_5_8_to_tile_6_8_2;
	wire vertical_tile_5_8_to_tile_6_8_3;
	wire vertical_tile_6_8_to_tile_5_8_0;
	wire vertical_tile_6_8_to_tile_5_8_1;
	wire vertical_tile_6_8_to_tile_5_8_2;
	wire vertical_tile_6_8_to_tile_5_8_3;

	wire vertical_tile_5_9_to_tile_6_9_0;
	wire vertical_tile_5_9_to_tile_6_9_1;
	wire vertical_tile_5_9_to_tile_6_9_2;
	wire vertical_tile_5_9_to_tile_6_9_3;
	wire vertical_tile_6_9_to_tile_5_9_0;
	wire vertical_tile_6_9_to_tile_5_9_1;
	wire vertical_tile_6_9_to_tile_5_9_2;
	wire vertical_tile_6_9_to_tile_5_9_3;

	wire vertical_tile_5_10_to_tile_6_10_0;
	wire vertical_tile_5_10_to_tile_6_10_1;
	wire vertical_tile_5_10_to_tile_6_10_2;
	wire vertical_tile_5_10_to_tile_6_10_3;
	wire vertical_tile_6_10_to_tile_5_10_0;
	wire vertical_tile_6_10_to_tile_5_10_1;
	wire vertical_tile_6_10_to_tile_5_10_2;
	wire vertical_tile_6_10_to_tile_5_10_3;

	wire vertical_tile_5_11_to_tile_6_11_0;
	wire vertical_tile_5_11_to_tile_6_11_1;
	wire vertical_tile_5_11_to_tile_6_11_2;
	wire vertical_tile_5_11_to_tile_6_11_3;
	wire vertical_tile_6_11_to_tile_5_11_0;
	wire vertical_tile_6_11_to_tile_5_11_1;
	wire vertical_tile_6_11_to_tile_5_11_2;
	wire vertical_tile_6_11_to_tile_5_11_3;

	wire vertical_tile_5_12_to_tile_6_12_0;
	wire vertical_tile_5_12_to_tile_6_12_1;
	wire vertical_tile_5_12_to_tile_6_12_2;
	wire vertical_tile_5_12_to_tile_6_12_3;
	wire vertical_tile_6_12_to_tile_5_12_0;
	wire vertical_tile_6_12_to_tile_5_12_1;
	wire vertical_tile_6_12_to_tile_5_12_2;
	wire vertical_tile_6_12_to_tile_5_12_3;

	wire vertical_tile_5_13_to_tile_6_13_0;
	wire vertical_tile_5_13_to_tile_6_13_1;
	wire vertical_tile_5_13_to_tile_6_13_2;
	wire vertical_tile_5_13_to_tile_6_13_3;
	wire vertical_tile_6_13_to_tile_5_13_0;
	wire vertical_tile_6_13_to_tile_5_13_1;
	wire vertical_tile_6_13_to_tile_5_13_2;
	wire vertical_tile_6_13_to_tile_5_13_3;

	wire vertical_tile_5_14_to_tile_6_14_0;
	wire vertical_tile_5_14_to_tile_6_14_1;
	wire vertical_tile_5_14_to_tile_6_14_2;
	wire vertical_tile_5_14_to_tile_6_14_3;
	wire vertical_tile_6_14_to_tile_5_14_0;
	wire vertical_tile_6_14_to_tile_5_14_1;
	wire vertical_tile_6_14_to_tile_5_14_2;
	wire vertical_tile_6_14_to_tile_5_14_3;

	wire vertical_tile_5_15_to_tile_6_15_0;
	wire vertical_tile_5_15_to_tile_6_15_1;
	wire vertical_tile_5_15_to_tile_6_15_2;
	wire vertical_tile_5_15_to_tile_6_15_3;
	wire vertical_tile_6_15_to_tile_5_15_0;
	wire vertical_tile_6_15_to_tile_5_15_1;
	wire vertical_tile_6_15_to_tile_5_15_2;
	wire vertical_tile_6_15_to_tile_5_15_3;

	wire vertical_tile_5_16_to_tile_6_16_0;
	wire vertical_tile_5_16_to_tile_6_16_1;
	wire vertical_tile_5_16_to_tile_6_16_2;
	wire vertical_tile_5_16_to_tile_6_16_3;
	wire vertical_tile_6_16_to_tile_5_16_0;
	wire vertical_tile_6_16_to_tile_5_16_1;
	wire vertical_tile_6_16_to_tile_5_16_2;
	wire vertical_tile_6_16_to_tile_5_16_3;

	wire vertical_tile_5_17_to_tile_6_17_0;
	wire vertical_tile_5_17_to_tile_6_17_1;
	wire vertical_tile_5_17_to_tile_6_17_2;
	wire vertical_tile_5_17_to_tile_6_17_3;
	wire vertical_tile_6_17_to_tile_5_17_0;
	wire vertical_tile_6_17_to_tile_5_17_1;
	wire vertical_tile_6_17_to_tile_5_17_2;
	wire vertical_tile_6_17_to_tile_5_17_3;

	wire vertical_tile_5_18_to_tile_6_18_0;
	wire vertical_tile_5_18_to_tile_6_18_1;
	wire vertical_tile_5_18_to_tile_6_18_2;
	wire vertical_tile_5_18_to_tile_6_18_3;
	wire vertical_tile_6_18_to_tile_5_18_0;
	wire vertical_tile_6_18_to_tile_5_18_1;
	wire vertical_tile_6_18_to_tile_5_18_2;
	wire vertical_tile_6_18_to_tile_5_18_3;

	wire vertical_tile_5_19_to_tile_6_19_0;
	wire vertical_tile_5_19_to_tile_6_19_1;
	wire vertical_tile_5_19_to_tile_6_19_2;
	wire vertical_tile_5_19_to_tile_6_19_3;
	wire vertical_tile_6_19_to_tile_5_19_0;
	wire vertical_tile_6_19_to_tile_5_19_1;
	wire vertical_tile_6_19_to_tile_5_19_2;
	wire vertical_tile_6_19_to_tile_5_19_3;

	wire vertical_tile_5_20_to_tile_6_20_0;
	wire vertical_tile_5_20_to_tile_6_20_1;
	wire vertical_tile_5_20_to_tile_6_20_2;
	wire vertical_tile_5_20_to_tile_6_20_3;
	wire vertical_tile_6_20_to_tile_5_20_0;
	wire vertical_tile_6_20_to_tile_5_20_1;
	wire vertical_tile_6_20_to_tile_5_20_2;
	wire vertical_tile_6_20_to_tile_5_20_3;

	wire vertical_tile_5_21_to_tile_6_21_0;
	wire vertical_tile_5_21_to_tile_6_21_1;
	wire vertical_tile_5_21_to_tile_6_21_2;
	wire vertical_tile_5_21_to_tile_6_21_3;
	wire vertical_tile_6_21_to_tile_5_21_0;
	wire vertical_tile_6_21_to_tile_5_21_1;
	wire vertical_tile_6_21_to_tile_5_21_2;
	wire vertical_tile_6_21_to_tile_5_21_3;

	wire vertical_tile_5_22_to_tile_6_22_0;
	wire vertical_tile_5_22_to_tile_6_22_1;
	wire vertical_tile_5_22_to_tile_6_22_2;
	wire vertical_tile_5_22_to_tile_6_22_3;
	wire vertical_tile_6_22_to_tile_5_22_0;
	wire vertical_tile_6_22_to_tile_5_22_1;
	wire vertical_tile_6_22_to_tile_5_22_2;
	wire vertical_tile_6_22_to_tile_5_22_3;

	wire vertical_tile_5_23_to_tile_6_23_0;
	wire vertical_tile_5_23_to_tile_6_23_1;
	wire vertical_tile_5_23_to_tile_6_23_2;
	wire vertical_tile_5_23_to_tile_6_23_3;
	wire vertical_tile_6_23_to_tile_5_23_0;
	wire vertical_tile_6_23_to_tile_5_23_1;
	wire vertical_tile_6_23_to_tile_5_23_2;
	wire vertical_tile_6_23_to_tile_5_23_3;

	wire vertical_tile_5_24_to_tile_6_24_0;
	wire vertical_tile_5_24_to_tile_6_24_1;
	wire vertical_tile_5_24_to_tile_6_24_2;
	wire vertical_tile_5_24_to_tile_6_24_3;
	wire vertical_tile_6_24_to_tile_5_24_0;
	wire vertical_tile_6_24_to_tile_5_24_1;
	wire vertical_tile_6_24_to_tile_5_24_2;
	wire vertical_tile_6_24_to_tile_5_24_3;

	wire vertical_tile_5_25_to_tile_6_25_0;
	wire vertical_tile_5_25_to_tile_6_25_1;
	wire vertical_tile_5_25_to_tile_6_25_2;
	wire vertical_tile_5_25_to_tile_6_25_3;
	wire vertical_tile_6_25_to_tile_5_25_0;
	wire vertical_tile_6_25_to_tile_5_25_1;
	wire vertical_tile_6_25_to_tile_5_25_2;
	wire vertical_tile_6_25_to_tile_5_25_3;

	wire vertical_tile_5_26_to_tile_6_26_0;
	wire vertical_tile_5_26_to_tile_6_26_1;
	wire vertical_tile_5_26_to_tile_6_26_2;
	wire vertical_tile_5_26_to_tile_6_26_3;
	wire vertical_tile_6_26_to_tile_5_26_0;
	wire vertical_tile_6_26_to_tile_5_26_1;
	wire vertical_tile_6_26_to_tile_5_26_2;
	wire vertical_tile_6_26_to_tile_5_26_3;

	wire vertical_tile_5_27_to_tile_6_27_0;
	wire vertical_tile_5_27_to_tile_6_27_1;
	wire vertical_tile_5_27_to_tile_6_27_2;
	wire vertical_tile_5_27_to_tile_6_27_3;
	wire vertical_tile_6_27_to_tile_5_27_0;
	wire vertical_tile_6_27_to_tile_5_27_1;
	wire vertical_tile_6_27_to_tile_5_27_2;
	wire vertical_tile_6_27_to_tile_5_27_3;

	wire vertical_tile_5_28_to_tile_6_28_0;
	wire vertical_tile_5_28_to_tile_6_28_1;
	wire vertical_tile_5_28_to_tile_6_28_2;
	wire vertical_tile_5_28_to_tile_6_28_3;
	wire vertical_tile_6_28_to_tile_5_28_0;
	wire vertical_tile_6_28_to_tile_5_28_1;
	wire vertical_tile_6_28_to_tile_5_28_2;
	wire vertical_tile_6_28_to_tile_5_28_3;

	wire vertical_tile_5_29_to_tile_6_29_0;
	wire vertical_tile_5_29_to_tile_6_29_1;
	wire vertical_tile_5_29_to_tile_6_29_2;
	wire vertical_tile_5_29_to_tile_6_29_3;
	wire vertical_tile_6_29_to_tile_5_29_0;
	wire vertical_tile_6_29_to_tile_5_29_1;
	wire vertical_tile_6_29_to_tile_5_29_2;
	wire vertical_tile_6_29_to_tile_5_29_3;

	wire vertical_tile_5_30_to_tile_6_30_0;
	wire vertical_tile_5_30_to_tile_6_30_1;
	wire vertical_tile_5_30_to_tile_6_30_2;
	wire vertical_tile_5_30_to_tile_6_30_3;
	wire vertical_tile_6_30_to_tile_5_30_0;
	wire vertical_tile_6_30_to_tile_5_30_1;
	wire vertical_tile_6_30_to_tile_5_30_2;
	wire vertical_tile_6_30_to_tile_5_30_3;

	wire vertical_tile_5_31_to_tile_6_31_0;
	wire vertical_tile_5_31_to_tile_6_31_1;
	wire vertical_tile_5_31_to_tile_6_31_2;
	wire vertical_tile_5_31_to_tile_6_31_3;
	wire vertical_tile_6_31_to_tile_5_31_0;
	wire vertical_tile_6_31_to_tile_5_31_1;
	wire vertical_tile_6_31_to_tile_5_31_2;
	wire vertical_tile_6_31_to_tile_5_31_3;

	wire vertical_tile_6_0_to_tile_7_0_0;
	wire vertical_tile_6_0_to_tile_7_0_1;
	wire vertical_tile_6_0_to_tile_7_0_2;
	wire vertical_tile_6_0_to_tile_7_0_3;
	wire vertical_tile_7_0_to_tile_6_0_0;
	wire vertical_tile_7_0_to_tile_6_0_1;
	wire vertical_tile_7_0_to_tile_6_0_2;
	wire vertical_tile_7_0_to_tile_6_0_3;

	wire vertical_tile_6_1_to_tile_7_1_0;
	wire vertical_tile_6_1_to_tile_7_1_1;
	wire vertical_tile_6_1_to_tile_7_1_2;
	wire vertical_tile_6_1_to_tile_7_1_3;
	wire vertical_tile_7_1_to_tile_6_1_0;
	wire vertical_tile_7_1_to_tile_6_1_1;
	wire vertical_tile_7_1_to_tile_6_1_2;
	wire vertical_tile_7_1_to_tile_6_1_3;

	wire vertical_tile_6_2_to_tile_7_2_0;
	wire vertical_tile_6_2_to_tile_7_2_1;
	wire vertical_tile_6_2_to_tile_7_2_2;
	wire vertical_tile_6_2_to_tile_7_2_3;
	wire vertical_tile_7_2_to_tile_6_2_0;
	wire vertical_tile_7_2_to_tile_6_2_1;
	wire vertical_tile_7_2_to_tile_6_2_2;
	wire vertical_tile_7_2_to_tile_6_2_3;

	wire vertical_tile_6_3_to_tile_7_3_0;
	wire vertical_tile_6_3_to_tile_7_3_1;
	wire vertical_tile_6_3_to_tile_7_3_2;
	wire vertical_tile_6_3_to_tile_7_3_3;
	wire vertical_tile_7_3_to_tile_6_3_0;
	wire vertical_tile_7_3_to_tile_6_3_1;
	wire vertical_tile_7_3_to_tile_6_3_2;
	wire vertical_tile_7_3_to_tile_6_3_3;

	wire vertical_tile_6_4_to_tile_7_4_0;
	wire vertical_tile_6_4_to_tile_7_4_1;
	wire vertical_tile_6_4_to_tile_7_4_2;
	wire vertical_tile_6_4_to_tile_7_4_3;
	wire vertical_tile_7_4_to_tile_6_4_0;
	wire vertical_tile_7_4_to_tile_6_4_1;
	wire vertical_tile_7_4_to_tile_6_4_2;
	wire vertical_tile_7_4_to_tile_6_4_3;

	wire vertical_tile_6_5_to_tile_7_5_0;
	wire vertical_tile_6_5_to_tile_7_5_1;
	wire vertical_tile_6_5_to_tile_7_5_2;
	wire vertical_tile_6_5_to_tile_7_5_3;
	wire vertical_tile_7_5_to_tile_6_5_0;
	wire vertical_tile_7_5_to_tile_6_5_1;
	wire vertical_tile_7_5_to_tile_6_5_2;
	wire vertical_tile_7_5_to_tile_6_5_3;

	wire vertical_tile_6_6_to_tile_7_6_0;
	wire vertical_tile_6_6_to_tile_7_6_1;
	wire vertical_tile_6_6_to_tile_7_6_2;
	wire vertical_tile_6_6_to_tile_7_6_3;
	wire vertical_tile_7_6_to_tile_6_6_0;
	wire vertical_tile_7_6_to_tile_6_6_1;
	wire vertical_tile_7_6_to_tile_6_6_2;
	wire vertical_tile_7_6_to_tile_6_6_3;

	wire vertical_tile_6_7_to_tile_7_7_0;
	wire vertical_tile_6_7_to_tile_7_7_1;
	wire vertical_tile_6_7_to_tile_7_7_2;
	wire vertical_tile_6_7_to_tile_7_7_3;
	wire vertical_tile_7_7_to_tile_6_7_0;
	wire vertical_tile_7_7_to_tile_6_7_1;
	wire vertical_tile_7_7_to_tile_6_7_2;
	wire vertical_tile_7_7_to_tile_6_7_3;

	wire vertical_tile_6_8_to_tile_7_8_0;
	wire vertical_tile_6_8_to_tile_7_8_1;
	wire vertical_tile_6_8_to_tile_7_8_2;
	wire vertical_tile_6_8_to_tile_7_8_3;
	wire vertical_tile_7_8_to_tile_6_8_0;
	wire vertical_tile_7_8_to_tile_6_8_1;
	wire vertical_tile_7_8_to_tile_6_8_2;
	wire vertical_tile_7_8_to_tile_6_8_3;

	wire vertical_tile_6_9_to_tile_7_9_0;
	wire vertical_tile_6_9_to_tile_7_9_1;
	wire vertical_tile_6_9_to_tile_7_9_2;
	wire vertical_tile_6_9_to_tile_7_9_3;
	wire vertical_tile_7_9_to_tile_6_9_0;
	wire vertical_tile_7_9_to_tile_6_9_1;
	wire vertical_tile_7_9_to_tile_6_9_2;
	wire vertical_tile_7_9_to_tile_6_9_3;

	wire vertical_tile_6_10_to_tile_7_10_0;
	wire vertical_tile_6_10_to_tile_7_10_1;
	wire vertical_tile_6_10_to_tile_7_10_2;
	wire vertical_tile_6_10_to_tile_7_10_3;
	wire vertical_tile_7_10_to_tile_6_10_0;
	wire vertical_tile_7_10_to_tile_6_10_1;
	wire vertical_tile_7_10_to_tile_6_10_2;
	wire vertical_tile_7_10_to_tile_6_10_3;

	wire vertical_tile_6_11_to_tile_7_11_0;
	wire vertical_tile_6_11_to_tile_7_11_1;
	wire vertical_tile_6_11_to_tile_7_11_2;
	wire vertical_tile_6_11_to_tile_7_11_3;
	wire vertical_tile_7_11_to_tile_6_11_0;
	wire vertical_tile_7_11_to_tile_6_11_1;
	wire vertical_tile_7_11_to_tile_6_11_2;
	wire vertical_tile_7_11_to_tile_6_11_3;

	wire vertical_tile_6_12_to_tile_7_12_0;
	wire vertical_tile_6_12_to_tile_7_12_1;
	wire vertical_tile_6_12_to_tile_7_12_2;
	wire vertical_tile_6_12_to_tile_7_12_3;
	wire vertical_tile_7_12_to_tile_6_12_0;
	wire vertical_tile_7_12_to_tile_6_12_1;
	wire vertical_tile_7_12_to_tile_6_12_2;
	wire vertical_tile_7_12_to_tile_6_12_3;

	wire vertical_tile_6_13_to_tile_7_13_0;
	wire vertical_tile_6_13_to_tile_7_13_1;
	wire vertical_tile_6_13_to_tile_7_13_2;
	wire vertical_tile_6_13_to_tile_7_13_3;
	wire vertical_tile_7_13_to_tile_6_13_0;
	wire vertical_tile_7_13_to_tile_6_13_1;
	wire vertical_tile_7_13_to_tile_6_13_2;
	wire vertical_tile_7_13_to_tile_6_13_3;

	wire vertical_tile_6_14_to_tile_7_14_0;
	wire vertical_tile_6_14_to_tile_7_14_1;
	wire vertical_tile_6_14_to_tile_7_14_2;
	wire vertical_tile_6_14_to_tile_7_14_3;
	wire vertical_tile_7_14_to_tile_6_14_0;
	wire vertical_tile_7_14_to_tile_6_14_1;
	wire vertical_tile_7_14_to_tile_6_14_2;
	wire vertical_tile_7_14_to_tile_6_14_3;

	wire vertical_tile_6_15_to_tile_7_15_0;
	wire vertical_tile_6_15_to_tile_7_15_1;
	wire vertical_tile_6_15_to_tile_7_15_2;
	wire vertical_tile_6_15_to_tile_7_15_3;
	wire vertical_tile_7_15_to_tile_6_15_0;
	wire vertical_tile_7_15_to_tile_6_15_1;
	wire vertical_tile_7_15_to_tile_6_15_2;
	wire vertical_tile_7_15_to_tile_6_15_3;

	wire vertical_tile_6_16_to_tile_7_16_0;
	wire vertical_tile_6_16_to_tile_7_16_1;
	wire vertical_tile_6_16_to_tile_7_16_2;
	wire vertical_tile_6_16_to_tile_7_16_3;
	wire vertical_tile_7_16_to_tile_6_16_0;
	wire vertical_tile_7_16_to_tile_6_16_1;
	wire vertical_tile_7_16_to_tile_6_16_2;
	wire vertical_tile_7_16_to_tile_6_16_3;

	wire vertical_tile_6_17_to_tile_7_17_0;
	wire vertical_tile_6_17_to_tile_7_17_1;
	wire vertical_tile_6_17_to_tile_7_17_2;
	wire vertical_tile_6_17_to_tile_7_17_3;
	wire vertical_tile_7_17_to_tile_6_17_0;
	wire vertical_tile_7_17_to_tile_6_17_1;
	wire vertical_tile_7_17_to_tile_6_17_2;
	wire vertical_tile_7_17_to_tile_6_17_3;

	wire vertical_tile_6_18_to_tile_7_18_0;
	wire vertical_tile_6_18_to_tile_7_18_1;
	wire vertical_tile_6_18_to_tile_7_18_2;
	wire vertical_tile_6_18_to_tile_7_18_3;
	wire vertical_tile_7_18_to_tile_6_18_0;
	wire vertical_tile_7_18_to_tile_6_18_1;
	wire vertical_tile_7_18_to_tile_6_18_2;
	wire vertical_tile_7_18_to_tile_6_18_3;

	wire vertical_tile_6_19_to_tile_7_19_0;
	wire vertical_tile_6_19_to_tile_7_19_1;
	wire vertical_tile_6_19_to_tile_7_19_2;
	wire vertical_tile_6_19_to_tile_7_19_3;
	wire vertical_tile_7_19_to_tile_6_19_0;
	wire vertical_tile_7_19_to_tile_6_19_1;
	wire vertical_tile_7_19_to_tile_6_19_2;
	wire vertical_tile_7_19_to_tile_6_19_3;

	wire vertical_tile_6_20_to_tile_7_20_0;
	wire vertical_tile_6_20_to_tile_7_20_1;
	wire vertical_tile_6_20_to_tile_7_20_2;
	wire vertical_tile_6_20_to_tile_7_20_3;
	wire vertical_tile_7_20_to_tile_6_20_0;
	wire vertical_tile_7_20_to_tile_6_20_1;
	wire vertical_tile_7_20_to_tile_6_20_2;
	wire vertical_tile_7_20_to_tile_6_20_3;

	wire vertical_tile_6_21_to_tile_7_21_0;
	wire vertical_tile_6_21_to_tile_7_21_1;
	wire vertical_tile_6_21_to_tile_7_21_2;
	wire vertical_tile_6_21_to_tile_7_21_3;
	wire vertical_tile_7_21_to_tile_6_21_0;
	wire vertical_tile_7_21_to_tile_6_21_1;
	wire vertical_tile_7_21_to_tile_6_21_2;
	wire vertical_tile_7_21_to_tile_6_21_3;

	wire vertical_tile_6_22_to_tile_7_22_0;
	wire vertical_tile_6_22_to_tile_7_22_1;
	wire vertical_tile_6_22_to_tile_7_22_2;
	wire vertical_tile_6_22_to_tile_7_22_3;
	wire vertical_tile_7_22_to_tile_6_22_0;
	wire vertical_tile_7_22_to_tile_6_22_1;
	wire vertical_tile_7_22_to_tile_6_22_2;
	wire vertical_tile_7_22_to_tile_6_22_3;

	wire vertical_tile_6_23_to_tile_7_23_0;
	wire vertical_tile_6_23_to_tile_7_23_1;
	wire vertical_tile_6_23_to_tile_7_23_2;
	wire vertical_tile_6_23_to_tile_7_23_3;
	wire vertical_tile_7_23_to_tile_6_23_0;
	wire vertical_tile_7_23_to_tile_6_23_1;
	wire vertical_tile_7_23_to_tile_6_23_2;
	wire vertical_tile_7_23_to_tile_6_23_3;

	wire vertical_tile_6_24_to_tile_7_24_0;
	wire vertical_tile_6_24_to_tile_7_24_1;
	wire vertical_tile_6_24_to_tile_7_24_2;
	wire vertical_tile_6_24_to_tile_7_24_3;
	wire vertical_tile_7_24_to_tile_6_24_0;
	wire vertical_tile_7_24_to_tile_6_24_1;
	wire vertical_tile_7_24_to_tile_6_24_2;
	wire vertical_tile_7_24_to_tile_6_24_3;

	wire vertical_tile_6_25_to_tile_7_25_0;
	wire vertical_tile_6_25_to_tile_7_25_1;
	wire vertical_tile_6_25_to_tile_7_25_2;
	wire vertical_tile_6_25_to_tile_7_25_3;
	wire vertical_tile_7_25_to_tile_6_25_0;
	wire vertical_tile_7_25_to_tile_6_25_1;
	wire vertical_tile_7_25_to_tile_6_25_2;
	wire vertical_tile_7_25_to_tile_6_25_3;

	wire vertical_tile_6_26_to_tile_7_26_0;
	wire vertical_tile_6_26_to_tile_7_26_1;
	wire vertical_tile_6_26_to_tile_7_26_2;
	wire vertical_tile_6_26_to_tile_7_26_3;
	wire vertical_tile_7_26_to_tile_6_26_0;
	wire vertical_tile_7_26_to_tile_6_26_1;
	wire vertical_tile_7_26_to_tile_6_26_2;
	wire vertical_tile_7_26_to_tile_6_26_3;

	wire vertical_tile_6_27_to_tile_7_27_0;
	wire vertical_tile_6_27_to_tile_7_27_1;
	wire vertical_tile_6_27_to_tile_7_27_2;
	wire vertical_tile_6_27_to_tile_7_27_3;
	wire vertical_tile_7_27_to_tile_6_27_0;
	wire vertical_tile_7_27_to_tile_6_27_1;
	wire vertical_tile_7_27_to_tile_6_27_2;
	wire vertical_tile_7_27_to_tile_6_27_3;

	wire vertical_tile_6_28_to_tile_7_28_0;
	wire vertical_tile_6_28_to_tile_7_28_1;
	wire vertical_tile_6_28_to_tile_7_28_2;
	wire vertical_tile_6_28_to_tile_7_28_3;
	wire vertical_tile_7_28_to_tile_6_28_0;
	wire vertical_tile_7_28_to_tile_6_28_1;
	wire vertical_tile_7_28_to_tile_6_28_2;
	wire vertical_tile_7_28_to_tile_6_28_3;

	wire vertical_tile_6_29_to_tile_7_29_0;
	wire vertical_tile_6_29_to_tile_7_29_1;
	wire vertical_tile_6_29_to_tile_7_29_2;
	wire vertical_tile_6_29_to_tile_7_29_3;
	wire vertical_tile_7_29_to_tile_6_29_0;
	wire vertical_tile_7_29_to_tile_6_29_1;
	wire vertical_tile_7_29_to_tile_6_29_2;
	wire vertical_tile_7_29_to_tile_6_29_3;

	wire vertical_tile_6_30_to_tile_7_30_0;
	wire vertical_tile_6_30_to_tile_7_30_1;
	wire vertical_tile_6_30_to_tile_7_30_2;
	wire vertical_tile_6_30_to_tile_7_30_3;
	wire vertical_tile_7_30_to_tile_6_30_0;
	wire vertical_tile_7_30_to_tile_6_30_1;
	wire vertical_tile_7_30_to_tile_6_30_2;
	wire vertical_tile_7_30_to_tile_6_30_3;

	wire vertical_tile_6_31_to_tile_7_31_0;
	wire vertical_tile_6_31_to_tile_7_31_1;
	wire vertical_tile_6_31_to_tile_7_31_2;
	wire vertical_tile_6_31_to_tile_7_31_3;
	wire vertical_tile_7_31_to_tile_6_31_0;
	wire vertical_tile_7_31_to_tile_6_31_1;
	wire vertical_tile_7_31_to_tile_6_31_2;
	wire vertical_tile_7_31_to_tile_6_31_3;

	wire vertical_tile_7_0_to_tile_8_0_0;
	wire vertical_tile_7_0_to_tile_8_0_1;
	wire vertical_tile_7_0_to_tile_8_0_2;
	wire vertical_tile_7_0_to_tile_8_0_3;
	wire vertical_tile_8_0_to_tile_7_0_0;
	wire vertical_tile_8_0_to_tile_7_0_1;
	wire vertical_tile_8_0_to_tile_7_0_2;
	wire vertical_tile_8_0_to_tile_7_0_3;

	wire vertical_tile_7_1_to_tile_8_1_0;
	wire vertical_tile_7_1_to_tile_8_1_1;
	wire vertical_tile_7_1_to_tile_8_1_2;
	wire vertical_tile_7_1_to_tile_8_1_3;
	wire vertical_tile_8_1_to_tile_7_1_0;
	wire vertical_tile_8_1_to_tile_7_1_1;
	wire vertical_tile_8_1_to_tile_7_1_2;
	wire vertical_tile_8_1_to_tile_7_1_3;

	wire vertical_tile_7_2_to_tile_8_2_0;
	wire vertical_tile_7_2_to_tile_8_2_1;
	wire vertical_tile_7_2_to_tile_8_2_2;
	wire vertical_tile_7_2_to_tile_8_2_3;
	wire vertical_tile_8_2_to_tile_7_2_0;
	wire vertical_tile_8_2_to_tile_7_2_1;
	wire vertical_tile_8_2_to_tile_7_2_2;
	wire vertical_tile_8_2_to_tile_7_2_3;

	wire vertical_tile_7_3_to_tile_8_3_0;
	wire vertical_tile_7_3_to_tile_8_3_1;
	wire vertical_tile_7_3_to_tile_8_3_2;
	wire vertical_tile_7_3_to_tile_8_3_3;
	wire vertical_tile_8_3_to_tile_7_3_0;
	wire vertical_tile_8_3_to_tile_7_3_1;
	wire vertical_tile_8_3_to_tile_7_3_2;
	wire vertical_tile_8_3_to_tile_7_3_3;

	wire vertical_tile_7_4_to_tile_8_4_0;
	wire vertical_tile_7_4_to_tile_8_4_1;
	wire vertical_tile_7_4_to_tile_8_4_2;
	wire vertical_tile_7_4_to_tile_8_4_3;
	wire vertical_tile_8_4_to_tile_7_4_0;
	wire vertical_tile_8_4_to_tile_7_4_1;
	wire vertical_tile_8_4_to_tile_7_4_2;
	wire vertical_tile_8_4_to_tile_7_4_3;

	wire vertical_tile_7_5_to_tile_8_5_0;
	wire vertical_tile_7_5_to_tile_8_5_1;
	wire vertical_tile_7_5_to_tile_8_5_2;
	wire vertical_tile_7_5_to_tile_8_5_3;
	wire vertical_tile_8_5_to_tile_7_5_0;
	wire vertical_tile_8_5_to_tile_7_5_1;
	wire vertical_tile_8_5_to_tile_7_5_2;
	wire vertical_tile_8_5_to_tile_7_5_3;

	wire vertical_tile_7_6_to_tile_8_6_0;
	wire vertical_tile_7_6_to_tile_8_6_1;
	wire vertical_tile_7_6_to_tile_8_6_2;
	wire vertical_tile_7_6_to_tile_8_6_3;
	wire vertical_tile_8_6_to_tile_7_6_0;
	wire vertical_tile_8_6_to_tile_7_6_1;
	wire vertical_tile_8_6_to_tile_7_6_2;
	wire vertical_tile_8_6_to_tile_7_6_3;

	wire vertical_tile_7_7_to_tile_8_7_0;
	wire vertical_tile_7_7_to_tile_8_7_1;
	wire vertical_tile_7_7_to_tile_8_7_2;
	wire vertical_tile_7_7_to_tile_8_7_3;
	wire vertical_tile_8_7_to_tile_7_7_0;
	wire vertical_tile_8_7_to_tile_7_7_1;
	wire vertical_tile_8_7_to_tile_7_7_2;
	wire vertical_tile_8_7_to_tile_7_7_3;

	wire vertical_tile_7_8_to_tile_8_8_0;
	wire vertical_tile_7_8_to_tile_8_8_1;
	wire vertical_tile_7_8_to_tile_8_8_2;
	wire vertical_tile_7_8_to_tile_8_8_3;
	wire vertical_tile_8_8_to_tile_7_8_0;
	wire vertical_tile_8_8_to_tile_7_8_1;
	wire vertical_tile_8_8_to_tile_7_8_2;
	wire vertical_tile_8_8_to_tile_7_8_3;

	wire vertical_tile_7_9_to_tile_8_9_0;
	wire vertical_tile_7_9_to_tile_8_9_1;
	wire vertical_tile_7_9_to_tile_8_9_2;
	wire vertical_tile_7_9_to_tile_8_9_3;
	wire vertical_tile_8_9_to_tile_7_9_0;
	wire vertical_tile_8_9_to_tile_7_9_1;
	wire vertical_tile_8_9_to_tile_7_9_2;
	wire vertical_tile_8_9_to_tile_7_9_3;

	wire vertical_tile_7_10_to_tile_8_10_0;
	wire vertical_tile_7_10_to_tile_8_10_1;
	wire vertical_tile_7_10_to_tile_8_10_2;
	wire vertical_tile_7_10_to_tile_8_10_3;
	wire vertical_tile_8_10_to_tile_7_10_0;
	wire vertical_tile_8_10_to_tile_7_10_1;
	wire vertical_tile_8_10_to_tile_7_10_2;
	wire vertical_tile_8_10_to_tile_7_10_3;

	wire vertical_tile_7_11_to_tile_8_11_0;
	wire vertical_tile_7_11_to_tile_8_11_1;
	wire vertical_tile_7_11_to_tile_8_11_2;
	wire vertical_tile_7_11_to_tile_8_11_3;
	wire vertical_tile_8_11_to_tile_7_11_0;
	wire vertical_tile_8_11_to_tile_7_11_1;
	wire vertical_tile_8_11_to_tile_7_11_2;
	wire vertical_tile_8_11_to_tile_7_11_3;

	wire vertical_tile_7_12_to_tile_8_12_0;
	wire vertical_tile_7_12_to_tile_8_12_1;
	wire vertical_tile_7_12_to_tile_8_12_2;
	wire vertical_tile_7_12_to_tile_8_12_3;
	wire vertical_tile_8_12_to_tile_7_12_0;
	wire vertical_tile_8_12_to_tile_7_12_1;
	wire vertical_tile_8_12_to_tile_7_12_2;
	wire vertical_tile_8_12_to_tile_7_12_3;

	wire vertical_tile_7_13_to_tile_8_13_0;
	wire vertical_tile_7_13_to_tile_8_13_1;
	wire vertical_tile_7_13_to_tile_8_13_2;
	wire vertical_tile_7_13_to_tile_8_13_3;
	wire vertical_tile_8_13_to_tile_7_13_0;
	wire vertical_tile_8_13_to_tile_7_13_1;
	wire vertical_tile_8_13_to_tile_7_13_2;
	wire vertical_tile_8_13_to_tile_7_13_3;

	wire vertical_tile_7_14_to_tile_8_14_0;
	wire vertical_tile_7_14_to_tile_8_14_1;
	wire vertical_tile_7_14_to_tile_8_14_2;
	wire vertical_tile_7_14_to_tile_8_14_3;
	wire vertical_tile_8_14_to_tile_7_14_0;
	wire vertical_tile_8_14_to_tile_7_14_1;
	wire vertical_tile_8_14_to_tile_7_14_2;
	wire vertical_tile_8_14_to_tile_7_14_3;

	wire vertical_tile_7_15_to_tile_8_15_0;
	wire vertical_tile_7_15_to_tile_8_15_1;
	wire vertical_tile_7_15_to_tile_8_15_2;
	wire vertical_tile_7_15_to_tile_8_15_3;
	wire vertical_tile_8_15_to_tile_7_15_0;
	wire vertical_tile_8_15_to_tile_7_15_1;
	wire vertical_tile_8_15_to_tile_7_15_2;
	wire vertical_tile_8_15_to_tile_7_15_3;

	wire vertical_tile_7_16_to_tile_8_16_0;
	wire vertical_tile_7_16_to_tile_8_16_1;
	wire vertical_tile_7_16_to_tile_8_16_2;
	wire vertical_tile_7_16_to_tile_8_16_3;
	wire vertical_tile_8_16_to_tile_7_16_0;
	wire vertical_tile_8_16_to_tile_7_16_1;
	wire vertical_tile_8_16_to_tile_7_16_2;
	wire vertical_tile_8_16_to_tile_7_16_3;

	wire vertical_tile_7_17_to_tile_8_17_0;
	wire vertical_tile_7_17_to_tile_8_17_1;
	wire vertical_tile_7_17_to_tile_8_17_2;
	wire vertical_tile_7_17_to_tile_8_17_3;
	wire vertical_tile_8_17_to_tile_7_17_0;
	wire vertical_tile_8_17_to_tile_7_17_1;
	wire vertical_tile_8_17_to_tile_7_17_2;
	wire vertical_tile_8_17_to_tile_7_17_3;

	wire vertical_tile_7_18_to_tile_8_18_0;
	wire vertical_tile_7_18_to_tile_8_18_1;
	wire vertical_tile_7_18_to_tile_8_18_2;
	wire vertical_tile_7_18_to_tile_8_18_3;
	wire vertical_tile_8_18_to_tile_7_18_0;
	wire vertical_tile_8_18_to_tile_7_18_1;
	wire vertical_tile_8_18_to_tile_7_18_2;
	wire vertical_tile_8_18_to_tile_7_18_3;

	wire vertical_tile_7_19_to_tile_8_19_0;
	wire vertical_tile_7_19_to_tile_8_19_1;
	wire vertical_tile_7_19_to_tile_8_19_2;
	wire vertical_tile_7_19_to_tile_8_19_3;
	wire vertical_tile_8_19_to_tile_7_19_0;
	wire vertical_tile_8_19_to_tile_7_19_1;
	wire vertical_tile_8_19_to_tile_7_19_2;
	wire vertical_tile_8_19_to_tile_7_19_3;

	wire vertical_tile_7_20_to_tile_8_20_0;
	wire vertical_tile_7_20_to_tile_8_20_1;
	wire vertical_tile_7_20_to_tile_8_20_2;
	wire vertical_tile_7_20_to_tile_8_20_3;
	wire vertical_tile_8_20_to_tile_7_20_0;
	wire vertical_tile_8_20_to_tile_7_20_1;
	wire vertical_tile_8_20_to_tile_7_20_2;
	wire vertical_tile_8_20_to_tile_7_20_3;

	wire vertical_tile_7_21_to_tile_8_21_0;
	wire vertical_tile_7_21_to_tile_8_21_1;
	wire vertical_tile_7_21_to_tile_8_21_2;
	wire vertical_tile_7_21_to_tile_8_21_3;
	wire vertical_tile_8_21_to_tile_7_21_0;
	wire vertical_tile_8_21_to_tile_7_21_1;
	wire vertical_tile_8_21_to_tile_7_21_2;
	wire vertical_tile_8_21_to_tile_7_21_3;

	wire vertical_tile_7_22_to_tile_8_22_0;
	wire vertical_tile_7_22_to_tile_8_22_1;
	wire vertical_tile_7_22_to_tile_8_22_2;
	wire vertical_tile_7_22_to_tile_8_22_3;
	wire vertical_tile_8_22_to_tile_7_22_0;
	wire vertical_tile_8_22_to_tile_7_22_1;
	wire vertical_tile_8_22_to_tile_7_22_2;
	wire vertical_tile_8_22_to_tile_7_22_3;

	wire vertical_tile_7_23_to_tile_8_23_0;
	wire vertical_tile_7_23_to_tile_8_23_1;
	wire vertical_tile_7_23_to_tile_8_23_2;
	wire vertical_tile_7_23_to_tile_8_23_3;
	wire vertical_tile_8_23_to_tile_7_23_0;
	wire vertical_tile_8_23_to_tile_7_23_1;
	wire vertical_tile_8_23_to_tile_7_23_2;
	wire vertical_tile_8_23_to_tile_7_23_3;

	wire vertical_tile_7_24_to_tile_8_24_0;
	wire vertical_tile_7_24_to_tile_8_24_1;
	wire vertical_tile_7_24_to_tile_8_24_2;
	wire vertical_tile_7_24_to_tile_8_24_3;
	wire vertical_tile_8_24_to_tile_7_24_0;
	wire vertical_tile_8_24_to_tile_7_24_1;
	wire vertical_tile_8_24_to_tile_7_24_2;
	wire vertical_tile_8_24_to_tile_7_24_3;

	wire vertical_tile_7_25_to_tile_8_25_0;
	wire vertical_tile_7_25_to_tile_8_25_1;
	wire vertical_tile_7_25_to_tile_8_25_2;
	wire vertical_tile_7_25_to_tile_8_25_3;
	wire vertical_tile_8_25_to_tile_7_25_0;
	wire vertical_tile_8_25_to_tile_7_25_1;
	wire vertical_tile_8_25_to_tile_7_25_2;
	wire vertical_tile_8_25_to_tile_7_25_3;

	wire vertical_tile_7_26_to_tile_8_26_0;
	wire vertical_tile_7_26_to_tile_8_26_1;
	wire vertical_tile_7_26_to_tile_8_26_2;
	wire vertical_tile_7_26_to_tile_8_26_3;
	wire vertical_tile_8_26_to_tile_7_26_0;
	wire vertical_tile_8_26_to_tile_7_26_1;
	wire vertical_tile_8_26_to_tile_7_26_2;
	wire vertical_tile_8_26_to_tile_7_26_3;

	wire vertical_tile_7_27_to_tile_8_27_0;
	wire vertical_tile_7_27_to_tile_8_27_1;
	wire vertical_tile_7_27_to_tile_8_27_2;
	wire vertical_tile_7_27_to_tile_8_27_3;
	wire vertical_tile_8_27_to_tile_7_27_0;
	wire vertical_tile_8_27_to_tile_7_27_1;
	wire vertical_tile_8_27_to_tile_7_27_2;
	wire vertical_tile_8_27_to_tile_7_27_3;

	wire vertical_tile_7_28_to_tile_8_28_0;
	wire vertical_tile_7_28_to_tile_8_28_1;
	wire vertical_tile_7_28_to_tile_8_28_2;
	wire vertical_tile_7_28_to_tile_8_28_3;
	wire vertical_tile_8_28_to_tile_7_28_0;
	wire vertical_tile_8_28_to_tile_7_28_1;
	wire vertical_tile_8_28_to_tile_7_28_2;
	wire vertical_tile_8_28_to_tile_7_28_3;

	wire vertical_tile_7_29_to_tile_8_29_0;
	wire vertical_tile_7_29_to_tile_8_29_1;
	wire vertical_tile_7_29_to_tile_8_29_2;
	wire vertical_tile_7_29_to_tile_8_29_3;
	wire vertical_tile_8_29_to_tile_7_29_0;
	wire vertical_tile_8_29_to_tile_7_29_1;
	wire vertical_tile_8_29_to_tile_7_29_2;
	wire vertical_tile_8_29_to_tile_7_29_3;

	wire vertical_tile_7_30_to_tile_8_30_0;
	wire vertical_tile_7_30_to_tile_8_30_1;
	wire vertical_tile_7_30_to_tile_8_30_2;
	wire vertical_tile_7_30_to_tile_8_30_3;
	wire vertical_tile_8_30_to_tile_7_30_0;
	wire vertical_tile_8_30_to_tile_7_30_1;
	wire vertical_tile_8_30_to_tile_7_30_2;
	wire vertical_tile_8_30_to_tile_7_30_3;

	wire vertical_tile_7_31_to_tile_8_31_0;
	wire vertical_tile_7_31_to_tile_8_31_1;
	wire vertical_tile_7_31_to_tile_8_31_2;
	wire vertical_tile_7_31_to_tile_8_31_3;
	wire vertical_tile_8_31_to_tile_7_31_0;
	wire vertical_tile_8_31_to_tile_7_31_1;
	wire vertical_tile_8_31_to_tile_7_31_2;
	wire vertical_tile_8_31_to_tile_7_31_3;

	wire vertical_tile_8_0_to_tile_9_0_0;
	wire vertical_tile_8_0_to_tile_9_0_1;
	wire vertical_tile_8_0_to_tile_9_0_2;
	wire vertical_tile_8_0_to_tile_9_0_3;
	wire vertical_tile_9_0_to_tile_8_0_0;
	wire vertical_tile_9_0_to_tile_8_0_1;
	wire vertical_tile_9_0_to_tile_8_0_2;
	wire vertical_tile_9_0_to_tile_8_0_3;

	wire vertical_tile_8_1_to_tile_9_1_0;
	wire vertical_tile_8_1_to_tile_9_1_1;
	wire vertical_tile_8_1_to_tile_9_1_2;
	wire vertical_tile_8_1_to_tile_9_1_3;
	wire vertical_tile_9_1_to_tile_8_1_0;
	wire vertical_tile_9_1_to_tile_8_1_1;
	wire vertical_tile_9_1_to_tile_8_1_2;
	wire vertical_tile_9_1_to_tile_8_1_3;

	wire vertical_tile_8_2_to_tile_9_2_0;
	wire vertical_tile_8_2_to_tile_9_2_1;
	wire vertical_tile_8_2_to_tile_9_2_2;
	wire vertical_tile_8_2_to_tile_9_2_3;
	wire vertical_tile_9_2_to_tile_8_2_0;
	wire vertical_tile_9_2_to_tile_8_2_1;
	wire vertical_tile_9_2_to_tile_8_2_2;
	wire vertical_tile_9_2_to_tile_8_2_3;

	wire vertical_tile_8_3_to_tile_9_3_0;
	wire vertical_tile_8_3_to_tile_9_3_1;
	wire vertical_tile_8_3_to_tile_9_3_2;
	wire vertical_tile_8_3_to_tile_9_3_3;
	wire vertical_tile_9_3_to_tile_8_3_0;
	wire vertical_tile_9_3_to_tile_8_3_1;
	wire vertical_tile_9_3_to_tile_8_3_2;
	wire vertical_tile_9_3_to_tile_8_3_3;

	wire vertical_tile_8_4_to_tile_9_4_0;
	wire vertical_tile_8_4_to_tile_9_4_1;
	wire vertical_tile_8_4_to_tile_9_4_2;
	wire vertical_tile_8_4_to_tile_9_4_3;
	wire vertical_tile_9_4_to_tile_8_4_0;
	wire vertical_tile_9_4_to_tile_8_4_1;
	wire vertical_tile_9_4_to_tile_8_4_2;
	wire vertical_tile_9_4_to_tile_8_4_3;

	wire vertical_tile_8_5_to_tile_9_5_0;
	wire vertical_tile_8_5_to_tile_9_5_1;
	wire vertical_tile_8_5_to_tile_9_5_2;
	wire vertical_tile_8_5_to_tile_9_5_3;
	wire vertical_tile_9_5_to_tile_8_5_0;
	wire vertical_tile_9_5_to_tile_8_5_1;
	wire vertical_tile_9_5_to_tile_8_5_2;
	wire vertical_tile_9_5_to_tile_8_5_3;

	wire vertical_tile_8_6_to_tile_9_6_0;
	wire vertical_tile_8_6_to_tile_9_6_1;
	wire vertical_tile_8_6_to_tile_9_6_2;
	wire vertical_tile_8_6_to_tile_9_6_3;
	wire vertical_tile_9_6_to_tile_8_6_0;
	wire vertical_tile_9_6_to_tile_8_6_1;
	wire vertical_tile_9_6_to_tile_8_6_2;
	wire vertical_tile_9_6_to_tile_8_6_3;

	wire vertical_tile_8_7_to_tile_9_7_0;
	wire vertical_tile_8_7_to_tile_9_7_1;
	wire vertical_tile_8_7_to_tile_9_7_2;
	wire vertical_tile_8_7_to_tile_9_7_3;
	wire vertical_tile_9_7_to_tile_8_7_0;
	wire vertical_tile_9_7_to_tile_8_7_1;
	wire vertical_tile_9_7_to_tile_8_7_2;
	wire vertical_tile_9_7_to_tile_8_7_3;

	wire vertical_tile_8_8_to_tile_9_8_0;
	wire vertical_tile_8_8_to_tile_9_8_1;
	wire vertical_tile_8_8_to_tile_9_8_2;
	wire vertical_tile_8_8_to_tile_9_8_3;
	wire vertical_tile_9_8_to_tile_8_8_0;
	wire vertical_tile_9_8_to_tile_8_8_1;
	wire vertical_tile_9_8_to_tile_8_8_2;
	wire vertical_tile_9_8_to_tile_8_8_3;

	wire vertical_tile_8_9_to_tile_9_9_0;
	wire vertical_tile_8_9_to_tile_9_9_1;
	wire vertical_tile_8_9_to_tile_9_9_2;
	wire vertical_tile_8_9_to_tile_9_9_3;
	wire vertical_tile_9_9_to_tile_8_9_0;
	wire vertical_tile_9_9_to_tile_8_9_1;
	wire vertical_tile_9_9_to_tile_8_9_2;
	wire vertical_tile_9_9_to_tile_8_9_3;

	wire vertical_tile_8_10_to_tile_9_10_0;
	wire vertical_tile_8_10_to_tile_9_10_1;
	wire vertical_tile_8_10_to_tile_9_10_2;
	wire vertical_tile_8_10_to_tile_9_10_3;
	wire vertical_tile_9_10_to_tile_8_10_0;
	wire vertical_tile_9_10_to_tile_8_10_1;
	wire vertical_tile_9_10_to_tile_8_10_2;
	wire vertical_tile_9_10_to_tile_8_10_3;

	wire vertical_tile_8_11_to_tile_9_11_0;
	wire vertical_tile_8_11_to_tile_9_11_1;
	wire vertical_tile_8_11_to_tile_9_11_2;
	wire vertical_tile_8_11_to_tile_9_11_3;
	wire vertical_tile_9_11_to_tile_8_11_0;
	wire vertical_tile_9_11_to_tile_8_11_1;
	wire vertical_tile_9_11_to_tile_8_11_2;
	wire vertical_tile_9_11_to_tile_8_11_3;

	wire vertical_tile_8_12_to_tile_9_12_0;
	wire vertical_tile_8_12_to_tile_9_12_1;
	wire vertical_tile_8_12_to_tile_9_12_2;
	wire vertical_tile_8_12_to_tile_9_12_3;
	wire vertical_tile_9_12_to_tile_8_12_0;
	wire vertical_tile_9_12_to_tile_8_12_1;
	wire vertical_tile_9_12_to_tile_8_12_2;
	wire vertical_tile_9_12_to_tile_8_12_3;

	wire vertical_tile_8_13_to_tile_9_13_0;
	wire vertical_tile_8_13_to_tile_9_13_1;
	wire vertical_tile_8_13_to_tile_9_13_2;
	wire vertical_tile_8_13_to_tile_9_13_3;
	wire vertical_tile_9_13_to_tile_8_13_0;
	wire vertical_tile_9_13_to_tile_8_13_1;
	wire vertical_tile_9_13_to_tile_8_13_2;
	wire vertical_tile_9_13_to_tile_8_13_3;

	wire vertical_tile_8_14_to_tile_9_14_0;
	wire vertical_tile_8_14_to_tile_9_14_1;
	wire vertical_tile_8_14_to_tile_9_14_2;
	wire vertical_tile_8_14_to_tile_9_14_3;
	wire vertical_tile_9_14_to_tile_8_14_0;
	wire vertical_tile_9_14_to_tile_8_14_1;
	wire vertical_tile_9_14_to_tile_8_14_2;
	wire vertical_tile_9_14_to_tile_8_14_3;

	wire vertical_tile_8_15_to_tile_9_15_0;
	wire vertical_tile_8_15_to_tile_9_15_1;
	wire vertical_tile_8_15_to_tile_9_15_2;
	wire vertical_tile_8_15_to_tile_9_15_3;
	wire vertical_tile_9_15_to_tile_8_15_0;
	wire vertical_tile_9_15_to_tile_8_15_1;
	wire vertical_tile_9_15_to_tile_8_15_2;
	wire vertical_tile_9_15_to_tile_8_15_3;

	wire vertical_tile_8_16_to_tile_9_16_0;
	wire vertical_tile_8_16_to_tile_9_16_1;
	wire vertical_tile_8_16_to_tile_9_16_2;
	wire vertical_tile_8_16_to_tile_9_16_3;
	wire vertical_tile_9_16_to_tile_8_16_0;
	wire vertical_tile_9_16_to_tile_8_16_1;
	wire vertical_tile_9_16_to_tile_8_16_2;
	wire vertical_tile_9_16_to_tile_8_16_3;

	wire vertical_tile_8_17_to_tile_9_17_0;
	wire vertical_tile_8_17_to_tile_9_17_1;
	wire vertical_tile_8_17_to_tile_9_17_2;
	wire vertical_tile_8_17_to_tile_9_17_3;
	wire vertical_tile_9_17_to_tile_8_17_0;
	wire vertical_tile_9_17_to_tile_8_17_1;
	wire vertical_tile_9_17_to_tile_8_17_2;
	wire vertical_tile_9_17_to_tile_8_17_3;

	wire vertical_tile_8_18_to_tile_9_18_0;
	wire vertical_tile_8_18_to_tile_9_18_1;
	wire vertical_tile_8_18_to_tile_9_18_2;
	wire vertical_tile_8_18_to_tile_9_18_3;
	wire vertical_tile_9_18_to_tile_8_18_0;
	wire vertical_tile_9_18_to_tile_8_18_1;
	wire vertical_tile_9_18_to_tile_8_18_2;
	wire vertical_tile_9_18_to_tile_8_18_3;

	wire vertical_tile_8_19_to_tile_9_19_0;
	wire vertical_tile_8_19_to_tile_9_19_1;
	wire vertical_tile_8_19_to_tile_9_19_2;
	wire vertical_tile_8_19_to_tile_9_19_3;
	wire vertical_tile_9_19_to_tile_8_19_0;
	wire vertical_tile_9_19_to_tile_8_19_1;
	wire vertical_tile_9_19_to_tile_8_19_2;
	wire vertical_tile_9_19_to_tile_8_19_3;

	wire vertical_tile_8_20_to_tile_9_20_0;
	wire vertical_tile_8_20_to_tile_9_20_1;
	wire vertical_tile_8_20_to_tile_9_20_2;
	wire vertical_tile_8_20_to_tile_9_20_3;
	wire vertical_tile_9_20_to_tile_8_20_0;
	wire vertical_tile_9_20_to_tile_8_20_1;
	wire vertical_tile_9_20_to_tile_8_20_2;
	wire vertical_tile_9_20_to_tile_8_20_3;

	wire vertical_tile_8_21_to_tile_9_21_0;
	wire vertical_tile_8_21_to_tile_9_21_1;
	wire vertical_tile_8_21_to_tile_9_21_2;
	wire vertical_tile_8_21_to_tile_9_21_3;
	wire vertical_tile_9_21_to_tile_8_21_0;
	wire vertical_tile_9_21_to_tile_8_21_1;
	wire vertical_tile_9_21_to_tile_8_21_2;
	wire vertical_tile_9_21_to_tile_8_21_3;

	wire vertical_tile_8_22_to_tile_9_22_0;
	wire vertical_tile_8_22_to_tile_9_22_1;
	wire vertical_tile_8_22_to_tile_9_22_2;
	wire vertical_tile_8_22_to_tile_9_22_3;
	wire vertical_tile_9_22_to_tile_8_22_0;
	wire vertical_tile_9_22_to_tile_8_22_1;
	wire vertical_tile_9_22_to_tile_8_22_2;
	wire vertical_tile_9_22_to_tile_8_22_3;

	wire vertical_tile_8_23_to_tile_9_23_0;
	wire vertical_tile_8_23_to_tile_9_23_1;
	wire vertical_tile_8_23_to_tile_9_23_2;
	wire vertical_tile_8_23_to_tile_9_23_3;
	wire vertical_tile_9_23_to_tile_8_23_0;
	wire vertical_tile_9_23_to_tile_8_23_1;
	wire vertical_tile_9_23_to_tile_8_23_2;
	wire vertical_tile_9_23_to_tile_8_23_3;

	wire vertical_tile_8_24_to_tile_9_24_0;
	wire vertical_tile_8_24_to_tile_9_24_1;
	wire vertical_tile_8_24_to_tile_9_24_2;
	wire vertical_tile_8_24_to_tile_9_24_3;
	wire vertical_tile_9_24_to_tile_8_24_0;
	wire vertical_tile_9_24_to_tile_8_24_1;
	wire vertical_tile_9_24_to_tile_8_24_2;
	wire vertical_tile_9_24_to_tile_8_24_3;

	wire vertical_tile_8_25_to_tile_9_25_0;
	wire vertical_tile_8_25_to_tile_9_25_1;
	wire vertical_tile_8_25_to_tile_9_25_2;
	wire vertical_tile_8_25_to_tile_9_25_3;
	wire vertical_tile_9_25_to_tile_8_25_0;
	wire vertical_tile_9_25_to_tile_8_25_1;
	wire vertical_tile_9_25_to_tile_8_25_2;
	wire vertical_tile_9_25_to_tile_8_25_3;

	wire vertical_tile_8_26_to_tile_9_26_0;
	wire vertical_tile_8_26_to_tile_9_26_1;
	wire vertical_tile_8_26_to_tile_9_26_2;
	wire vertical_tile_8_26_to_tile_9_26_3;
	wire vertical_tile_9_26_to_tile_8_26_0;
	wire vertical_tile_9_26_to_tile_8_26_1;
	wire vertical_tile_9_26_to_tile_8_26_2;
	wire vertical_tile_9_26_to_tile_8_26_3;

	wire vertical_tile_8_27_to_tile_9_27_0;
	wire vertical_tile_8_27_to_tile_9_27_1;
	wire vertical_tile_8_27_to_tile_9_27_2;
	wire vertical_tile_8_27_to_tile_9_27_3;
	wire vertical_tile_9_27_to_tile_8_27_0;
	wire vertical_tile_9_27_to_tile_8_27_1;
	wire vertical_tile_9_27_to_tile_8_27_2;
	wire vertical_tile_9_27_to_tile_8_27_3;

	wire vertical_tile_8_28_to_tile_9_28_0;
	wire vertical_tile_8_28_to_tile_9_28_1;
	wire vertical_tile_8_28_to_tile_9_28_2;
	wire vertical_tile_8_28_to_tile_9_28_3;
	wire vertical_tile_9_28_to_tile_8_28_0;
	wire vertical_tile_9_28_to_tile_8_28_1;
	wire vertical_tile_9_28_to_tile_8_28_2;
	wire vertical_tile_9_28_to_tile_8_28_3;

	wire vertical_tile_8_29_to_tile_9_29_0;
	wire vertical_tile_8_29_to_tile_9_29_1;
	wire vertical_tile_8_29_to_tile_9_29_2;
	wire vertical_tile_8_29_to_tile_9_29_3;
	wire vertical_tile_9_29_to_tile_8_29_0;
	wire vertical_tile_9_29_to_tile_8_29_1;
	wire vertical_tile_9_29_to_tile_8_29_2;
	wire vertical_tile_9_29_to_tile_8_29_3;

	wire vertical_tile_8_30_to_tile_9_30_0;
	wire vertical_tile_8_30_to_tile_9_30_1;
	wire vertical_tile_8_30_to_tile_9_30_2;
	wire vertical_tile_8_30_to_tile_9_30_3;
	wire vertical_tile_9_30_to_tile_8_30_0;
	wire vertical_tile_9_30_to_tile_8_30_1;
	wire vertical_tile_9_30_to_tile_8_30_2;
	wire vertical_tile_9_30_to_tile_8_30_3;

	wire vertical_tile_8_31_to_tile_9_31_0;
	wire vertical_tile_8_31_to_tile_9_31_1;
	wire vertical_tile_8_31_to_tile_9_31_2;
	wire vertical_tile_8_31_to_tile_9_31_3;
	wire vertical_tile_9_31_to_tile_8_31_0;
	wire vertical_tile_9_31_to_tile_8_31_1;
	wire vertical_tile_9_31_to_tile_8_31_2;
	wire vertical_tile_9_31_to_tile_8_31_3;

	wire vertical_tile_9_0_to_tile_10_0_0;
	wire vertical_tile_9_0_to_tile_10_0_1;
	wire vertical_tile_9_0_to_tile_10_0_2;
	wire vertical_tile_9_0_to_tile_10_0_3;
	wire vertical_tile_10_0_to_tile_9_0_0;
	wire vertical_tile_10_0_to_tile_9_0_1;
	wire vertical_tile_10_0_to_tile_9_0_2;
	wire vertical_tile_10_0_to_tile_9_0_3;

	wire vertical_tile_9_1_to_tile_10_1_0;
	wire vertical_tile_9_1_to_tile_10_1_1;
	wire vertical_tile_9_1_to_tile_10_1_2;
	wire vertical_tile_9_1_to_tile_10_1_3;
	wire vertical_tile_10_1_to_tile_9_1_0;
	wire vertical_tile_10_1_to_tile_9_1_1;
	wire vertical_tile_10_1_to_tile_9_1_2;
	wire vertical_tile_10_1_to_tile_9_1_3;

	wire vertical_tile_9_2_to_tile_10_2_0;
	wire vertical_tile_9_2_to_tile_10_2_1;
	wire vertical_tile_9_2_to_tile_10_2_2;
	wire vertical_tile_9_2_to_tile_10_2_3;
	wire vertical_tile_10_2_to_tile_9_2_0;
	wire vertical_tile_10_2_to_tile_9_2_1;
	wire vertical_tile_10_2_to_tile_9_2_2;
	wire vertical_tile_10_2_to_tile_9_2_3;

	wire vertical_tile_9_3_to_tile_10_3_0;
	wire vertical_tile_9_3_to_tile_10_3_1;
	wire vertical_tile_9_3_to_tile_10_3_2;
	wire vertical_tile_9_3_to_tile_10_3_3;
	wire vertical_tile_10_3_to_tile_9_3_0;
	wire vertical_tile_10_3_to_tile_9_3_1;
	wire vertical_tile_10_3_to_tile_9_3_2;
	wire vertical_tile_10_3_to_tile_9_3_3;

	wire vertical_tile_9_4_to_tile_10_4_0;
	wire vertical_tile_9_4_to_tile_10_4_1;
	wire vertical_tile_9_4_to_tile_10_4_2;
	wire vertical_tile_9_4_to_tile_10_4_3;
	wire vertical_tile_10_4_to_tile_9_4_0;
	wire vertical_tile_10_4_to_tile_9_4_1;
	wire vertical_tile_10_4_to_tile_9_4_2;
	wire vertical_tile_10_4_to_tile_9_4_3;

	wire vertical_tile_9_5_to_tile_10_5_0;
	wire vertical_tile_9_5_to_tile_10_5_1;
	wire vertical_tile_9_5_to_tile_10_5_2;
	wire vertical_tile_9_5_to_tile_10_5_3;
	wire vertical_tile_10_5_to_tile_9_5_0;
	wire vertical_tile_10_5_to_tile_9_5_1;
	wire vertical_tile_10_5_to_tile_9_5_2;
	wire vertical_tile_10_5_to_tile_9_5_3;

	wire vertical_tile_9_6_to_tile_10_6_0;
	wire vertical_tile_9_6_to_tile_10_6_1;
	wire vertical_tile_9_6_to_tile_10_6_2;
	wire vertical_tile_9_6_to_tile_10_6_3;
	wire vertical_tile_10_6_to_tile_9_6_0;
	wire vertical_tile_10_6_to_tile_9_6_1;
	wire vertical_tile_10_6_to_tile_9_6_2;
	wire vertical_tile_10_6_to_tile_9_6_3;

	wire vertical_tile_9_7_to_tile_10_7_0;
	wire vertical_tile_9_7_to_tile_10_7_1;
	wire vertical_tile_9_7_to_tile_10_7_2;
	wire vertical_tile_9_7_to_tile_10_7_3;
	wire vertical_tile_10_7_to_tile_9_7_0;
	wire vertical_tile_10_7_to_tile_9_7_1;
	wire vertical_tile_10_7_to_tile_9_7_2;
	wire vertical_tile_10_7_to_tile_9_7_3;

	wire vertical_tile_9_8_to_tile_10_8_0;
	wire vertical_tile_9_8_to_tile_10_8_1;
	wire vertical_tile_9_8_to_tile_10_8_2;
	wire vertical_tile_9_8_to_tile_10_8_3;
	wire vertical_tile_10_8_to_tile_9_8_0;
	wire vertical_tile_10_8_to_tile_9_8_1;
	wire vertical_tile_10_8_to_tile_9_8_2;
	wire vertical_tile_10_8_to_tile_9_8_3;

	wire vertical_tile_9_9_to_tile_10_9_0;
	wire vertical_tile_9_9_to_tile_10_9_1;
	wire vertical_tile_9_9_to_tile_10_9_2;
	wire vertical_tile_9_9_to_tile_10_9_3;
	wire vertical_tile_10_9_to_tile_9_9_0;
	wire vertical_tile_10_9_to_tile_9_9_1;
	wire vertical_tile_10_9_to_tile_9_9_2;
	wire vertical_tile_10_9_to_tile_9_9_3;

	wire vertical_tile_9_10_to_tile_10_10_0;
	wire vertical_tile_9_10_to_tile_10_10_1;
	wire vertical_tile_9_10_to_tile_10_10_2;
	wire vertical_tile_9_10_to_tile_10_10_3;
	wire vertical_tile_10_10_to_tile_9_10_0;
	wire vertical_tile_10_10_to_tile_9_10_1;
	wire vertical_tile_10_10_to_tile_9_10_2;
	wire vertical_tile_10_10_to_tile_9_10_3;

	wire vertical_tile_9_11_to_tile_10_11_0;
	wire vertical_tile_9_11_to_tile_10_11_1;
	wire vertical_tile_9_11_to_tile_10_11_2;
	wire vertical_tile_9_11_to_tile_10_11_3;
	wire vertical_tile_10_11_to_tile_9_11_0;
	wire vertical_tile_10_11_to_tile_9_11_1;
	wire vertical_tile_10_11_to_tile_9_11_2;
	wire vertical_tile_10_11_to_tile_9_11_3;

	wire vertical_tile_9_12_to_tile_10_12_0;
	wire vertical_tile_9_12_to_tile_10_12_1;
	wire vertical_tile_9_12_to_tile_10_12_2;
	wire vertical_tile_9_12_to_tile_10_12_3;
	wire vertical_tile_10_12_to_tile_9_12_0;
	wire vertical_tile_10_12_to_tile_9_12_1;
	wire vertical_tile_10_12_to_tile_9_12_2;
	wire vertical_tile_10_12_to_tile_9_12_3;

	wire vertical_tile_9_13_to_tile_10_13_0;
	wire vertical_tile_9_13_to_tile_10_13_1;
	wire vertical_tile_9_13_to_tile_10_13_2;
	wire vertical_tile_9_13_to_tile_10_13_3;
	wire vertical_tile_10_13_to_tile_9_13_0;
	wire vertical_tile_10_13_to_tile_9_13_1;
	wire vertical_tile_10_13_to_tile_9_13_2;
	wire vertical_tile_10_13_to_tile_9_13_3;

	wire vertical_tile_9_14_to_tile_10_14_0;
	wire vertical_tile_9_14_to_tile_10_14_1;
	wire vertical_tile_9_14_to_tile_10_14_2;
	wire vertical_tile_9_14_to_tile_10_14_3;
	wire vertical_tile_10_14_to_tile_9_14_0;
	wire vertical_tile_10_14_to_tile_9_14_1;
	wire vertical_tile_10_14_to_tile_9_14_2;
	wire vertical_tile_10_14_to_tile_9_14_3;

	wire vertical_tile_9_15_to_tile_10_15_0;
	wire vertical_tile_9_15_to_tile_10_15_1;
	wire vertical_tile_9_15_to_tile_10_15_2;
	wire vertical_tile_9_15_to_tile_10_15_3;
	wire vertical_tile_10_15_to_tile_9_15_0;
	wire vertical_tile_10_15_to_tile_9_15_1;
	wire vertical_tile_10_15_to_tile_9_15_2;
	wire vertical_tile_10_15_to_tile_9_15_3;

	wire vertical_tile_9_16_to_tile_10_16_0;
	wire vertical_tile_9_16_to_tile_10_16_1;
	wire vertical_tile_9_16_to_tile_10_16_2;
	wire vertical_tile_9_16_to_tile_10_16_3;
	wire vertical_tile_10_16_to_tile_9_16_0;
	wire vertical_tile_10_16_to_tile_9_16_1;
	wire vertical_tile_10_16_to_tile_9_16_2;
	wire vertical_tile_10_16_to_tile_9_16_3;

	wire vertical_tile_9_17_to_tile_10_17_0;
	wire vertical_tile_9_17_to_tile_10_17_1;
	wire vertical_tile_9_17_to_tile_10_17_2;
	wire vertical_tile_9_17_to_tile_10_17_3;
	wire vertical_tile_10_17_to_tile_9_17_0;
	wire vertical_tile_10_17_to_tile_9_17_1;
	wire vertical_tile_10_17_to_tile_9_17_2;
	wire vertical_tile_10_17_to_tile_9_17_3;

	wire vertical_tile_9_18_to_tile_10_18_0;
	wire vertical_tile_9_18_to_tile_10_18_1;
	wire vertical_tile_9_18_to_tile_10_18_2;
	wire vertical_tile_9_18_to_tile_10_18_3;
	wire vertical_tile_10_18_to_tile_9_18_0;
	wire vertical_tile_10_18_to_tile_9_18_1;
	wire vertical_tile_10_18_to_tile_9_18_2;
	wire vertical_tile_10_18_to_tile_9_18_3;

	wire vertical_tile_9_19_to_tile_10_19_0;
	wire vertical_tile_9_19_to_tile_10_19_1;
	wire vertical_tile_9_19_to_tile_10_19_2;
	wire vertical_tile_9_19_to_tile_10_19_3;
	wire vertical_tile_10_19_to_tile_9_19_0;
	wire vertical_tile_10_19_to_tile_9_19_1;
	wire vertical_tile_10_19_to_tile_9_19_2;
	wire vertical_tile_10_19_to_tile_9_19_3;

	wire vertical_tile_9_20_to_tile_10_20_0;
	wire vertical_tile_9_20_to_tile_10_20_1;
	wire vertical_tile_9_20_to_tile_10_20_2;
	wire vertical_tile_9_20_to_tile_10_20_3;
	wire vertical_tile_10_20_to_tile_9_20_0;
	wire vertical_tile_10_20_to_tile_9_20_1;
	wire vertical_tile_10_20_to_tile_9_20_2;
	wire vertical_tile_10_20_to_tile_9_20_3;

	wire vertical_tile_9_21_to_tile_10_21_0;
	wire vertical_tile_9_21_to_tile_10_21_1;
	wire vertical_tile_9_21_to_tile_10_21_2;
	wire vertical_tile_9_21_to_tile_10_21_3;
	wire vertical_tile_10_21_to_tile_9_21_0;
	wire vertical_tile_10_21_to_tile_9_21_1;
	wire vertical_tile_10_21_to_tile_9_21_2;
	wire vertical_tile_10_21_to_tile_9_21_3;

	wire vertical_tile_9_22_to_tile_10_22_0;
	wire vertical_tile_9_22_to_tile_10_22_1;
	wire vertical_tile_9_22_to_tile_10_22_2;
	wire vertical_tile_9_22_to_tile_10_22_3;
	wire vertical_tile_10_22_to_tile_9_22_0;
	wire vertical_tile_10_22_to_tile_9_22_1;
	wire vertical_tile_10_22_to_tile_9_22_2;
	wire vertical_tile_10_22_to_tile_9_22_3;

	wire vertical_tile_9_23_to_tile_10_23_0;
	wire vertical_tile_9_23_to_tile_10_23_1;
	wire vertical_tile_9_23_to_tile_10_23_2;
	wire vertical_tile_9_23_to_tile_10_23_3;
	wire vertical_tile_10_23_to_tile_9_23_0;
	wire vertical_tile_10_23_to_tile_9_23_1;
	wire vertical_tile_10_23_to_tile_9_23_2;
	wire vertical_tile_10_23_to_tile_9_23_3;

	wire vertical_tile_9_24_to_tile_10_24_0;
	wire vertical_tile_9_24_to_tile_10_24_1;
	wire vertical_tile_9_24_to_tile_10_24_2;
	wire vertical_tile_9_24_to_tile_10_24_3;
	wire vertical_tile_10_24_to_tile_9_24_0;
	wire vertical_tile_10_24_to_tile_9_24_1;
	wire vertical_tile_10_24_to_tile_9_24_2;
	wire vertical_tile_10_24_to_tile_9_24_3;

	wire vertical_tile_9_25_to_tile_10_25_0;
	wire vertical_tile_9_25_to_tile_10_25_1;
	wire vertical_tile_9_25_to_tile_10_25_2;
	wire vertical_tile_9_25_to_tile_10_25_3;
	wire vertical_tile_10_25_to_tile_9_25_0;
	wire vertical_tile_10_25_to_tile_9_25_1;
	wire vertical_tile_10_25_to_tile_9_25_2;
	wire vertical_tile_10_25_to_tile_9_25_3;

	wire vertical_tile_9_26_to_tile_10_26_0;
	wire vertical_tile_9_26_to_tile_10_26_1;
	wire vertical_tile_9_26_to_tile_10_26_2;
	wire vertical_tile_9_26_to_tile_10_26_3;
	wire vertical_tile_10_26_to_tile_9_26_0;
	wire vertical_tile_10_26_to_tile_9_26_1;
	wire vertical_tile_10_26_to_tile_9_26_2;
	wire vertical_tile_10_26_to_tile_9_26_3;

	wire vertical_tile_9_27_to_tile_10_27_0;
	wire vertical_tile_9_27_to_tile_10_27_1;
	wire vertical_tile_9_27_to_tile_10_27_2;
	wire vertical_tile_9_27_to_tile_10_27_3;
	wire vertical_tile_10_27_to_tile_9_27_0;
	wire vertical_tile_10_27_to_tile_9_27_1;
	wire vertical_tile_10_27_to_tile_9_27_2;
	wire vertical_tile_10_27_to_tile_9_27_3;

	wire vertical_tile_9_28_to_tile_10_28_0;
	wire vertical_tile_9_28_to_tile_10_28_1;
	wire vertical_tile_9_28_to_tile_10_28_2;
	wire vertical_tile_9_28_to_tile_10_28_3;
	wire vertical_tile_10_28_to_tile_9_28_0;
	wire vertical_tile_10_28_to_tile_9_28_1;
	wire vertical_tile_10_28_to_tile_9_28_2;
	wire vertical_tile_10_28_to_tile_9_28_3;

	wire vertical_tile_9_29_to_tile_10_29_0;
	wire vertical_tile_9_29_to_tile_10_29_1;
	wire vertical_tile_9_29_to_tile_10_29_2;
	wire vertical_tile_9_29_to_tile_10_29_3;
	wire vertical_tile_10_29_to_tile_9_29_0;
	wire vertical_tile_10_29_to_tile_9_29_1;
	wire vertical_tile_10_29_to_tile_9_29_2;
	wire vertical_tile_10_29_to_tile_9_29_3;

	wire vertical_tile_9_30_to_tile_10_30_0;
	wire vertical_tile_9_30_to_tile_10_30_1;
	wire vertical_tile_9_30_to_tile_10_30_2;
	wire vertical_tile_9_30_to_tile_10_30_3;
	wire vertical_tile_10_30_to_tile_9_30_0;
	wire vertical_tile_10_30_to_tile_9_30_1;
	wire vertical_tile_10_30_to_tile_9_30_2;
	wire vertical_tile_10_30_to_tile_9_30_3;

	wire vertical_tile_9_31_to_tile_10_31_0;
	wire vertical_tile_9_31_to_tile_10_31_1;
	wire vertical_tile_9_31_to_tile_10_31_2;
	wire vertical_tile_9_31_to_tile_10_31_3;
	wire vertical_tile_10_31_to_tile_9_31_0;
	wire vertical_tile_10_31_to_tile_9_31_1;
	wire vertical_tile_10_31_to_tile_9_31_2;
	wire vertical_tile_10_31_to_tile_9_31_3;

	wire vertical_tile_10_0_to_tile_11_0_0;
	wire vertical_tile_10_0_to_tile_11_0_1;
	wire vertical_tile_10_0_to_tile_11_0_2;
	wire vertical_tile_10_0_to_tile_11_0_3;
	wire vertical_tile_11_0_to_tile_10_0_0;
	wire vertical_tile_11_0_to_tile_10_0_1;
	wire vertical_tile_11_0_to_tile_10_0_2;
	wire vertical_tile_11_0_to_tile_10_0_3;

	wire vertical_tile_10_1_to_tile_11_1_0;
	wire vertical_tile_10_1_to_tile_11_1_1;
	wire vertical_tile_10_1_to_tile_11_1_2;
	wire vertical_tile_10_1_to_tile_11_1_3;
	wire vertical_tile_11_1_to_tile_10_1_0;
	wire vertical_tile_11_1_to_tile_10_1_1;
	wire vertical_tile_11_1_to_tile_10_1_2;
	wire vertical_tile_11_1_to_tile_10_1_3;

	wire vertical_tile_10_2_to_tile_11_2_0;
	wire vertical_tile_10_2_to_tile_11_2_1;
	wire vertical_tile_10_2_to_tile_11_2_2;
	wire vertical_tile_10_2_to_tile_11_2_3;
	wire vertical_tile_11_2_to_tile_10_2_0;
	wire vertical_tile_11_2_to_tile_10_2_1;
	wire vertical_tile_11_2_to_tile_10_2_2;
	wire vertical_tile_11_2_to_tile_10_2_3;

	wire vertical_tile_10_3_to_tile_11_3_0;
	wire vertical_tile_10_3_to_tile_11_3_1;
	wire vertical_tile_10_3_to_tile_11_3_2;
	wire vertical_tile_10_3_to_tile_11_3_3;
	wire vertical_tile_11_3_to_tile_10_3_0;
	wire vertical_tile_11_3_to_tile_10_3_1;
	wire vertical_tile_11_3_to_tile_10_3_2;
	wire vertical_tile_11_3_to_tile_10_3_3;

	wire vertical_tile_10_4_to_tile_11_4_0;
	wire vertical_tile_10_4_to_tile_11_4_1;
	wire vertical_tile_10_4_to_tile_11_4_2;
	wire vertical_tile_10_4_to_tile_11_4_3;
	wire vertical_tile_11_4_to_tile_10_4_0;
	wire vertical_tile_11_4_to_tile_10_4_1;
	wire vertical_tile_11_4_to_tile_10_4_2;
	wire vertical_tile_11_4_to_tile_10_4_3;

	wire vertical_tile_10_5_to_tile_11_5_0;
	wire vertical_tile_10_5_to_tile_11_5_1;
	wire vertical_tile_10_5_to_tile_11_5_2;
	wire vertical_tile_10_5_to_tile_11_5_3;
	wire vertical_tile_11_5_to_tile_10_5_0;
	wire vertical_tile_11_5_to_tile_10_5_1;
	wire vertical_tile_11_5_to_tile_10_5_2;
	wire vertical_tile_11_5_to_tile_10_5_3;

	wire vertical_tile_10_6_to_tile_11_6_0;
	wire vertical_tile_10_6_to_tile_11_6_1;
	wire vertical_tile_10_6_to_tile_11_6_2;
	wire vertical_tile_10_6_to_tile_11_6_3;
	wire vertical_tile_11_6_to_tile_10_6_0;
	wire vertical_tile_11_6_to_tile_10_6_1;
	wire vertical_tile_11_6_to_tile_10_6_2;
	wire vertical_tile_11_6_to_tile_10_6_3;

	wire vertical_tile_10_7_to_tile_11_7_0;
	wire vertical_tile_10_7_to_tile_11_7_1;
	wire vertical_tile_10_7_to_tile_11_7_2;
	wire vertical_tile_10_7_to_tile_11_7_3;
	wire vertical_tile_11_7_to_tile_10_7_0;
	wire vertical_tile_11_7_to_tile_10_7_1;
	wire vertical_tile_11_7_to_tile_10_7_2;
	wire vertical_tile_11_7_to_tile_10_7_3;

	wire vertical_tile_10_8_to_tile_11_8_0;
	wire vertical_tile_10_8_to_tile_11_8_1;
	wire vertical_tile_10_8_to_tile_11_8_2;
	wire vertical_tile_10_8_to_tile_11_8_3;
	wire vertical_tile_11_8_to_tile_10_8_0;
	wire vertical_tile_11_8_to_tile_10_8_1;
	wire vertical_tile_11_8_to_tile_10_8_2;
	wire vertical_tile_11_8_to_tile_10_8_3;

	wire vertical_tile_10_9_to_tile_11_9_0;
	wire vertical_tile_10_9_to_tile_11_9_1;
	wire vertical_tile_10_9_to_tile_11_9_2;
	wire vertical_tile_10_9_to_tile_11_9_3;
	wire vertical_tile_11_9_to_tile_10_9_0;
	wire vertical_tile_11_9_to_tile_10_9_1;
	wire vertical_tile_11_9_to_tile_10_9_2;
	wire vertical_tile_11_9_to_tile_10_9_3;

	wire vertical_tile_10_10_to_tile_11_10_0;
	wire vertical_tile_10_10_to_tile_11_10_1;
	wire vertical_tile_10_10_to_tile_11_10_2;
	wire vertical_tile_10_10_to_tile_11_10_3;
	wire vertical_tile_11_10_to_tile_10_10_0;
	wire vertical_tile_11_10_to_tile_10_10_1;
	wire vertical_tile_11_10_to_tile_10_10_2;
	wire vertical_tile_11_10_to_tile_10_10_3;

	wire vertical_tile_10_11_to_tile_11_11_0;
	wire vertical_tile_10_11_to_tile_11_11_1;
	wire vertical_tile_10_11_to_tile_11_11_2;
	wire vertical_tile_10_11_to_tile_11_11_3;
	wire vertical_tile_11_11_to_tile_10_11_0;
	wire vertical_tile_11_11_to_tile_10_11_1;
	wire vertical_tile_11_11_to_tile_10_11_2;
	wire vertical_tile_11_11_to_tile_10_11_3;

	wire vertical_tile_10_12_to_tile_11_12_0;
	wire vertical_tile_10_12_to_tile_11_12_1;
	wire vertical_tile_10_12_to_tile_11_12_2;
	wire vertical_tile_10_12_to_tile_11_12_3;
	wire vertical_tile_11_12_to_tile_10_12_0;
	wire vertical_tile_11_12_to_tile_10_12_1;
	wire vertical_tile_11_12_to_tile_10_12_2;
	wire vertical_tile_11_12_to_tile_10_12_3;

	wire vertical_tile_10_13_to_tile_11_13_0;
	wire vertical_tile_10_13_to_tile_11_13_1;
	wire vertical_tile_10_13_to_tile_11_13_2;
	wire vertical_tile_10_13_to_tile_11_13_3;
	wire vertical_tile_11_13_to_tile_10_13_0;
	wire vertical_tile_11_13_to_tile_10_13_1;
	wire vertical_tile_11_13_to_tile_10_13_2;
	wire vertical_tile_11_13_to_tile_10_13_3;

	wire vertical_tile_10_14_to_tile_11_14_0;
	wire vertical_tile_10_14_to_tile_11_14_1;
	wire vertical_tile_10_14_to_tile_11_14_2;
	wire vertical_tile_10_14_to_tile_11_14_3;
	wire vertical_tile_11_14_to_tile_10_14_0;
	wire vertical_tile_11_14_to_tile_10_14_1;
	wire vertical_tile_11_14_to_tile_10_14_2;
	wire vertical_tile_11_14_to_tile_10_14_3;

	wire vertical_tile_10_15_to_tile_11_15_0;
	wire vertical_tile_10_15_to_tile_11_15_1;
	wire vertical_tile_10_15_to_tile_11_15_2;
	wire vertical_tile_10_15_to_tile_11_15_3;
	wire vertical_tile_11_15_to_tile_10_15_0;
	wire vertical_tile_11_15_to_tile_10_15_1;
	wire vertical_tile_11_15_to_tile_10_15_2;
	wire vertical_tile_11_15_to_tile_10_15_3;

	wire vertical_tile_10_16_to_tile_11_16_0;
	wire vertical_tile_10_16_to_tile_11_16_1;
	wire vertical_tile_10_16_to_tile_11_16_2;
	wire vertical_tile_10_16_to_tile_11_16_3;
	wire vertical_tile_11_16_to_tile_10_16_0;
	wire vertical_tile_11_16_to_tile_10_16_1;
	wire vertical_tile_11_16_to_tile_10_16_2;
	wire vertical_tile_11_16_to_tile_10_16_3;

	wire vertical_tile_10_17_to_tile_11_17_0;
	wire vertical_tile_10_17_to_tile_11_17_1;
	wire vertical_tile_10_17_to_tile_11_17_2;
	wire vertical_tile_10_17_to_tile_11_17_3;
	wire vertical_tile_11_17_to_tile_10_17_0;
	wire vertical_tile_11_17_to_tile_10_17_1;
	wire vertical_tile_11_17_to_tile_10_17_2;
	wire vertical_tile_11_17_to_tile_10_17_3;

	wire vertical_tile_10_18_to_tile_11_18_0;
	wire vertical_tile_10_18_to_tile_11_18_1;
	wire vertical_tile_10_18_to_tile_11_18_2;
	wire vertical_tile_10_18_to_tile_11_18_3;
	wire vertical_tile_11_18_to_tile_10_18_0;
	wire vertical_tile_11_18_to_tile_10_18_1;
	wire vertical_tile_11_18_to_tile_10_18_2;
	wire vertical_tile_11_18_to_tile_10_18_3;

	wire vertical_tile_10_19_to_tile_11_19_0;
	wire vertical_tile_10_19_to_tile_11_19_1;
	wire vertical_tile_10_19_to_tile_11_19_2;
	wire vertical_tile_10_19_to_tile_11_19_3;
	wire vertical_tile_11_19_to_tile_10_19_0;
	wire vertical_tile_11_19_to_tile_10_19_1;
	wire vertical_tile_11_19_to_tile_10_19_2;
	wire vertical_tile_11_19_to_tile_10_19_3;

	wire vertical_tile_10_20_to_tile_11_20_0;
	wire vertical_tile_10_20_to_tile_11_20_1;
	wire vertical_tile_10_20_to_tile_11_20_2;
	wire vertical_tile_10_20_to_tile_11_20_3;
	wire vertical_tile_11_20_to_tile_10_20_0;
	wire vertical_tile_11_20_to_tile_10_20_1;
	wire vertical_tile_11_20_to_tile_10_20_2;
	wire vertical_tile_11_20_to_tile_10_20_3;

	wire vertical_tile_10_21_to_tile_11_21_0;
	wire vertical_tile_10_21_to_tile_11_21_1;
	wire vertical_tile_10_21_to_tile_11_21_2;
	wire vertical_tile_10_21_to_tile_11_21_3;
	wire vertical_tile_11_21_to_tile_10_21_0;
	wire vertical_tile_11_21_to_tile_10_21_1;
	wire vertical_tile_11_21_to_tile_10_21_2;
	wire vertical_tile_11_21_to_tile_10_21_3;

	wire vertical_tile_10_22_to_tile_11_22_0;
	wire vertical_tile_10_22_to_tile_11_22_1;
	wire vertical_tile_10_22_to_tile_11_22_2;
	wire vertical_tile_10_22_to_tile_11_22_3;
	wire vertical_tile_11_22_to_tile_10_22_0;
	wire vertical_tile_11_22_to_tile_10_22_1;
	wire vertical_tile_11_22_to_tile_10_22_2;
	wire vertical_tile_11_22_to_tile_10_22_3;

	wire vertical_tile_10_23_to_tile_11_23_0;
	wire vertical_tile_10_23_to_tile_11_23_1;
	wire vertical_tile_10_23_to_tile_11_23_2;
	wire vertical_tile_10_23_to_tile_11_23_3;
	wire vertical_tile_11_23_to_tile_10_23_0;
	wire vertical_tile_11_23_to_tile_10_23_1;
	wire vertical_tile_11_23_to_tile_10_23_2;
	wire vertical_tile_11_23_to_tile_10_23_3;

	wire vertical_tile_10_24_to_tile_11_24_0;
	wire vertical_tile_10_24_to_tile_11_24_1;
	wire vertical_tile_10_24_to_tile_11_24_2;
	wire vertical_tile_10_24_to_tile_11_24_3;
	wire vertical_tile_11_24_to_tile_10_24_0;
	wire vertical_tile_11_24_to_tile_10_24_1;
	wire vertical_tile_11_24_to_tile_10_24_2;
	wire vertical_tile_11_24_to_tile_10_24_3;

	wire vertical_tile_10_25_to_tile_11_25_0;
	wire vertical_tile_10_25_to_tile_11_25_1;
	wire vertical_tile_10_25_to_tile_11_25_2;
	wire vertical_tile_10_25_to_tile_11_25_3;
	wire vertical_tile_11_25_to_tile_10_25_0;
	wire vertical_tile_11_25_to_tile_10_25_1;
	wire vertical_tile_11_25_to_tile_10_25_2;
	wire vertical_tile_11_25_to_tile_10_25_3;

	wire vertical_tile_10_26_to_tile_11_26_0;
	wire vertical_tile_10_26_to_tile_11_26_1;
	wire vertical_tile_10_26_to_tile_11_26_2;
	wire vertical_tile_10_26_to_tile_11_26_3;
	wire vertical_tile_11_26_to_tile_10_26_0;
	wire vertical_tile_11_26_to_tile_10_26_1;
	wire vertical_tile_11_26_to_tile_10_26_2;
	wire vertical_tile_11_26_to_tile_10_26_3;

	wire vertical_tile_10_27_to_tile_11_27_0;
	wire vertical_tile_10_27_to_tile_11_27_1;
	wire vertical_tile_10_27_to_tile_11_27_2;
	wire vertical_tile_10_27_to_tile_11_27_3;
	wire vertical_tile_11_27_to_tile_10_27_0;
	wire vertical_tile_11_27_to_tile_10_27_1;
	wire vertical_tile_11_27_to_tile_10_27_2;
	wire vertical_tile_11_27_to_tile_10_27_3;

	wire vertical_tile_10_28_to_tile_11_28_0;
	wire vertical_tile_10_28_to_tile_11_28_1;
	wire vertical_tile_10_28_to_tile_11_28_2;
	wire vertical_tile_10_28_to_tile_11_28_3;
	wire vertical_tile_11_28_to_tile_10_28_0;
	wire vertical_tile_11_28_to_tile_10_28_1;
	wire vertical_tile_11_28_to_tile_10_28_2;
	wire vertical_tile_11_28_to_tile_10_28_3;

	wire vertical_tile_10_29_to_tile_11_29_0;
	wire vertical_tile_10_29_to_tile_11_29_1;
	wire vertical_tile_10_29_to_tile_11_29_2;
	wire vertical_tile_10_29_to_tile_11_29_3;
	wire vertical_tile_11_29_to_tile_10_29_0;
	wire vertical_tile_11_29_to_tile_10_29_1;
	wire vertical_tile_11_29_to_tile_10_29_2;
	wire vertical_tile_11_29_to_tile_10_29_3;

	wire vertical_tile_10_30_to_tile_11_30_0;
	wire vertical_tile_10_30_to_tile_11_30_1;
	wire vertical_tile_10_30_to_tile_11_30_2;
	wire vertical_tile_10_30_to_tile_11_30_3;
	wire vertical_tile_11_30_to_tile_10_30_0;
	wire vertical_tile_11_30_to_tile_10_30_1;
	wire vertical_tile_11_30_to_tile_10_30_2;
	wire vertical_tile_11_30_to_tile_10_30_3;

	wire vertical_tile_10_31_to_tile_11_31_0;
	wire vertical_tile_10_31_to_tile_11_31_1;
	wire vertical_tile_10_31_to_tile_11_31_2;
	wire vertical_tile_10_31_to_tile_11_31_3;
	wire vertical_tile_11_31_to_tile_10_31_0;
	wire vertical_tile_11_31_to_tile_10_31_1;
	wire vertical_tile_11_31_to_tile_10_31_2;
	wire vertical_tile_11_31_to_tile_10_31_3;

	wire vertical_tile_11_0_to_tile_12_0_0;
	wire vertical_tile_11_0_to_tile_12_0_1;
	wire vertical_tile_11_0_to_tile_12_0_2;
	wire vertical_tile_11_0_to_tile_12_0_3;
	wire vertical_tile_12_0_to_tile_11_0_0;
	wire vertical_tile_12_0_to_tile_11_0_1;
	wire vertical_tile_12_0_to_tile_11_0_2;
	wire vertical_tile_12_0_to_tile_11_0_3;

	wire vertical_tile_11_1_to_tile_12_1_0;
	wire vertical_tile_11_1_to_tile_12_1_1;
	wire vertical_tile_11_1_to_tile_12_1_2;
	wire vertical_tile_11_1_to_tile_12_1_3;
	wire vertical_tile_12_1_to_tile_11_1_0;
	wire vertical_tile_12_1_to_tile_11_1_1;
	wire vertical_tile_12_1_to_tile_11_1_2;
	wire vertical_tile_12_1_to_tile_11_1_3;

	wire vertical_tile_11_2_to_tile_12_2_0;
	wire vertical_tile_11_2_to_tile_12_2_1;
	wire vertical_tile_11_2_to_tile_12_2_2;
	wire vertical_tile_11_2_to_tile_12_2_3;
	wire vertical_tile_12_2_to_tile_11_2_0;
	wire vertical_tile_12_2_to_tile_11_2_1;
	wire vertical_tile_12_2_to_tile_11_2_2;
	wire vertical_tile_12_2_to_tile_11_2_3;

	wire vertical_tile_11_3_to_tile_12_3_0;
	wire vertical_tile_11_3_to_tile_12_3_1;
	wire vertical_tile_11_3_to_tile_12_3_2;
	wire vertical_tile_11_3_to_tile_12_3_3;
	wire vertical_tile_12_3_to_tile_11_3_0;
	wire vertical_tile_12_3_to_tile_11_3_1;
	wire vertical_tile_12_3_to_tile_11_3_2;
	wire vertical_tile_12_3_to_tile_11_3_3;

	wire vertical_tile_11_4_to_tile_12_4_0;
	wire vertical_tile_11_4_to_tile_12_4_1;
	wire vertical_tile_11_4_to_tile_12_4_2;
	wire vertical_tile_11_4_to_tile_12_4_3;
	wire vertical_tile_12_4_to_tile_11_4_0;
	wire vertical_tile_12_4_to_tile_11_4_1;
	wire vertical_tile_12_4_to_tile_11_4_2;
	wire vertical_tile_12_4_to_tile_11_4_3;

	wire vertical_tile_11_5_to_tile_12_5_0;
	wire vertical_tile_11_5_to_tile_12_5_1;
	wire vertical_tile_11_5_to_tile_12_5_2;
	wire vertical_tile_11_5_to_tile_12_5_3;
	wire vertical_tile_12_5_to_tile_11_5_0;
	wire vertical_tile_12_5_to_tile_11_5_1;
	wire vertical_tile_12_5_to_tile_11_5_2;
	wire vertical_tile_12_5_to_tile_11_5_3;

	wire vertical_tile_11_6_to_tile_12_6_0;
	wire vertical_tile_11_6_to_tile_12_6_1;
	wire vertical_tile_11_6_to_tile_12_6_2;
	wire vertical_tile_11_6_to_tile_12_6_3;
	wire vertical_tile_12_6_to_tile_11_6_0;
	wire vertical_tile_12_6_to_tile_11_6_1;
	wire vertical_tile_12_6_to_tile_11_6_2;
	wire vertical_tile_12_6_to_tile_11_6_3;

	wire vertical_tile_11_7_to_tile_12_7_0;
	wire vertical_tile_11_7_to_tile_12_7_1;
	wire vertical_tile_11_7_to_tile_12_7_2;
	wire vertical_tile_11_7_to_tile_12_7_3;
	wire vertical_tile_12_7_to_tile_11_7_0;
	wire vertical_tile_12_7_to_tile_11_7_1;
	wire vertical_tile_12_7_to_tile_11_7_2;
	wire vertical_tile_12_7_to_tile_11_7_3;

	wire vertical_tile_11_8_to_tile_12_8_0;
	wire vertical_tile_11_8_to_tile_12_8_1;
	wire vertical_tile_11_8_to_tile_12_8_2;
	wire vertical_tile_11_8_to_tile_12_8_3;
	wire vertical_tile_12_8_to_tile_11_8_0;
	wire vertical_tile_12_8_to_tile_11_8_1;
	wire vertical_tile_12_8_to_tile_11_8_2;
	wire vertical_tile_12_8_to_tile_11_8_3;

	wire vertical_tile_11_9_to_tile_12_9_0;
	wire vertical_tile_11_9_to_tile_12_9_1;
	wire vertical_tile_11_9_to_tile_12_9_2;
	wire vertical_tile_11_9_to_tile_12_9_3;
	wire vertical_tile_12_9_to_tile_11_9_0;
	wire vertical_tile_12_9_to_tile_11_9_1;
	wire vertical_tile_12_9_to_tile_11_9_2;
	wire vertical_tile_12_9_to_tile_11_9_3;

	wire vertical_tile_11_10_to_tile_12_10_0;
	wire vertical_tile_11_10_to_tile_12_10_1;
	wire vertical_tile_11_10_to_tile_12_10_2;
	wire vertical_tile_11_10_to_tile_12_10_3;
	wire vertical_tile_12_10_to_tile_11_10_0;
	wire vertical_tile_12_10_to_tile_11_10_1;
	wire vertical_tile_12_10_to_tile_11_10_2;
	wire vertical_tile_12_10_to_tile_11_10_3;

	wire vertical_tile_11_11_to_tile_12_11_0;
	wire vertical_tile_11_11_to_tile_12_11_1;
	wire vertical_tile_11_11_to_tile_12_11_2;
	wire vertical_tile_11_11_to_tile_12_11_3;
	wire vertical_tile_12_11_to_tile_11_11_0;
	wire vertical_tile_12_11_to_tile_11_11_1;
	wire vertical_tile_12_11_to_tile_11_11_2;
	wire vertical_tile_12_11_to_tile_11_11_3;

	wire vertical_tile_11_12_to_tile_12_12_0;
	wire vertical_tile_11_12_to_tile_12_12_1;
	wire vertical_tile_11_12_to_tile_12_12_2;
	wire vertical_tile_11_12_to_tile_12_12_3;
	wire vertical_tile_12_12_to_tile_11_12_0;
	wire vertical_tile_12_12_to_tile_11_12_1;
	wire vertical_tile_12_12_to_tile_11_12_2;
	wire vertical_tile_12_12_to_tile_11_12_3;

	wire vertical_tile_11_13_to_tile_12_13_0;
	wire vertical_tile_11_13_to_tile_12_13_1;
	wire vertical_tile_11_13_to_tile_12_13_2;
	wire vertical_tile_11_13_to_tile_12_13_3;
	wire vertical_tile_12_13_to_tile_11_13_0;
	wire vertical_tile_12_13_to_tile_11_13_1;
	wire vertical_tile_12_13_to_tile_11_13_2;
	wire vertical_tile_12_13_to_tile_11_13_3;

	wire vertical_tile_11_14_to_tile_12_14_0;
	wire vertical_tile_11_14_to_tile_12_14_1;
	wire vertical_tile_11_14_to_tile_12_14_2;
	wire vertical_tile_11_14_to_tile_12_14_3;
	wire vertical_tile_12_14_to_tile_11_14_0;
	wire vertical_tile_12_14_to_tile_11_14_1;
	wire vertical_tile_12_14_to_tile_11_14_2;
	wire vertical_tile_12_14_to_tile_11_14_3;

	wire vertical_tile_11_15_to_tile_12_15_0;
	wire vertical_tile_11_15_to_tile_12_15_1;
	wire vertical_tile_11_15_to_tile_12_15_2;
	wire vertical_tile_11_15_to_tile_12_15_3;
	wire vertical_tile_12_15_to_tile_11_15_0;
	wire vertical_tile_12_15_to_tile_11_15_1;
	wire vertical_tile_12_15_to_tile_11_15_2;
	wire vertical_tile_12_15_to_tile_11_15_3;

	wire vertical_tile_11_16_to_tile_12_16_0;
	wire vertical_tile_11_16_to_tile_12_16_1;
	wire vertical_tile_11_16_to_tile_12_16_2;
	wire vertical_tile_11_16_to_tile_12_16_3;
	wire vertical_tile_12_16_to_tile_11_16_0;
	wire vertical_tile_12_16_to_tile_11_16_1;
	wire vertical_tile_12_16_to_tile_11_16_2;
	wire vertical_tile_12_16_to_tile_11_16_3;

	wire vertical_tile_11_17_to_tile_12_17_0;
	wire vertical_tile_11_17_to_tile_12_17_1;
	wire vertical_tile_11_17_to_tile_12_17_2;
	wire vertical_tile_11_17_to_tile_12_17_3;
	wire vertical_tile_12_17_to_tile_11_17_0;
	wire vertical_tile_12_17_to_tile_11_17_1;
	wire vertical_tile_12_17_to_tile_11_17_2;
	wire vertical_tile_12_17_to_tile_11_17_3;

	wire vertical_tile_11_18_to_tile_12_18_0;
	wire vertical_tile_11_18_to_tile_12_18_1;
	wire vertical_tile_11_18_to_tile_12_18_2;
	wire vertical_tile_11_18_to_tile_12_18_3;
	wire vertical_tile_12_18_to_tile_11_18_0;
	wire vertical_tile_12_18_to_tile_11_18_1;
	wire vertical_tile_12_18_to_tile_11_18_2;
	wire vertical_tile_12_18_to_tile_11_18_3;

	wire vertical_tile_11_19_to_tile_12_19_0;
	wire vertical_tile_11_19_to_tile_12_19_1;
	wire vertical_tile_11_19_to_tile_12_19_2;
	wire vertical_tile_11_19_to_tile_12_19_3;
	wire vertical_tile_12_19_to_tile_11_19_0;
	wire vertical_tile_12_19_to_tile_11_19_1;
	wire vertical_tile_12_19_to_tile_11_19_2;
	wire vertical_tile_12_19_to_tile_11_19_3;

	wire vertical_tile_11_20_to_tile_12_20_0;
	wire vertical_tile_11_20_to_tile_12_20_1;
	wire vertical_tile_11_20_to_tile_12_20_2;
	wire vertical_tile_11_20_to_tile_12_20_3;
	wire vertical_tile_12_20_to_tile_11_20_0;
	wire vertical_tile_12_20_to_tile_11_20_1;
	wire vertical_tile_12_20_to_tile_11_20_2;
	wire vertical_tile_12_20_to_tile_11_20_3;

	wire vertical_tile_11_21_to_tile_12_21_0;
	wire vertical_tile_11_21_to_tile_12_21_1;
	wire vertical_tile_11_21_to_tile_12_21_2;
	wire vertical_tile_11_21_to_tile_12_21_3;
	wire vertical_tile_12_21_to_tile_11_21_0;
	wire vertical_tile_12_21_to_tile_11_21_1;
	wire vertical_tile_12_21_to_tile_11_21_2;
	wire vertical_tile_12_21_to_tile_11_21_3;

	wire vertical_tile_11_22_to_tile_12_22_0;
	wire vertical_tile_11_22_to_tile_12_22_1;
	wire vertical_tile_11_22_to_tile_12_22_2;
	wire vertical_tile_11_22_to_tile_12_22_3;
	wire vertical_tile_12_22_to_tile_11_22_0;
	wire vertical_tile_12_22_to_tile_11_22_1;
	wire vertical_tile_12_22_to_tile_11_22_2;
	wire vertical_tile_12_22_to_tile_11_22_3;

	wire vertical_tile_11_23_to_tile_12_23_0;
	wire vertical_tile_11_23_to_tile_12_23_1;
	wire vertical_tile_11_23_to_tile_12_23_2;
	wire vertical_tile_11_23_to_tile_12_23_3;
	wire vertical_tile_12_23_to_tile_11_23_0;
	wire vertical_tile_12_23_to_tile_11_23_1;
	wire vertical_tile_12_23_to_tile_11_23_2;
	wire vertical_tile_12_23_to_tile_11_23_3;

	wire vertical_tile_11_24_to_tile_12_24_0;
	wire vertical_tile_11_24_to_tile_12_24_1;
	wire vertical_tile_11_24_to_tile_12_24_2;
	wire vertical_tile_11_24_to_tile_12_24_3;
	wire vertical_tile_12_24_to_tile_11_24_0;
	wire vertical_tile_12_24_to_tile_11_24_1;
	wire vertical_tile_12_24_to_tile_11_24_2;
	wire vertical_tile_12_24_to_tile_11_24_3;

	wire vertical_tile_11_25_to_tile_12_25_0;
	wire vertical_tile_11_25_to_tile_12_25_1;
	wire vertical_tile_11_25_to_tile_12_25_2;
	wire vertical_tile_11_25_to_tile_12_25_3;
	wire vertical_tile_12_25_to_tile_11_25_0;
	wire vertical_tile_12_25_to_tile_11_25_1;
	wire vertical_tile_12_25_to_tile_11_25_2;
	wire vertical_tile_12_25_to_tile_11_25_3;

	wire vertical_tile_11_26_to_tile_12_26_0;
	wire vertical_tile_11_26_to_tile_12_26_1;
	wire vertical_tile_11_26_to_tile_12_26_2;
	wire vertical_tile_11_26_to_tile_12_26_3;
	wire vertical_tile_12_26_to_tile_11_26_0;
	wire vertical_tile_12_26_to_tile_11_26_1;
	wire vertical_tile_12_26_to_tile_11_26_2;
	wire vertical_tile_12_26_to_tile_11_26_3;

	wire vertical_tile_11_27_to_tile_12_27_0;
	wire vertical_tile_11_27_to_tile_12_27_1;
	wire vertical_tile_11_27_to_tile_12_27_2;
	wire vertical_tile_11_27_to_tile_12_27_3;
	wire vertical_tile_12_27_to_tile_11_27_0;
	wire vertical_tile_12_27_to_tile_11_27_1;
	wire vertical_tile_12_27_to_tile_11_27_2;
	wire vertical_tile_12_27_to_tile_11_27_3;

	wire vertical_tile_11_28_to_tile_12_28_0;
	wire vertical_tile_11_28_to_tile_12_28_1;
	wire vertical_tile_11_28_to_tile_12_28_2;
	wire vertical_tile_11_28_to_tile_12_28_3;
	wire vertical_tile_12_28_to_tile_11_28_0;
	wire vertical_tile_12_28_to_tile_11_28_1;
	wire vertical_tile_12_28_to_tile_11_28_2;
	wire vertical_tile_12_28_to_tile_11_28_3;

	wire vertical_tile_11_29_to_tile_12_29_0;
	wire vertical_tile_11_29_to_tile_12_29_1;
	wire vertical_tile_11_29_to_tile_12_29_2;
	wire vertical_tile_11_29_to_tile_12_29_3;
	wire vertical_tile_12_29_to_tile_11_29_0;
	wire vertical_tile_12_29_to_tile_11_29_1;
	wire vertical_tile_12_29_to_tile_11_29_2;
	wire vertical_tile_12_29_to_tile_11_29_3;

	wire vertical_tile_11_30_to_tile_12_30_0;
	wire vertical_tile_11_30_to_tile_12_30_1;
	wire vertical_tile_11_30_to_tile_12_30_2;
	wire vertical_tile_11_30_to_tile_12_30_3;
	wire vertical_tile_12_30_to_tile_11_30_0;
	wire vertical_tile_12_30_to_tile_11_30_1;
	wire vertical_tile_12_30_to_tile_11_30_2;
	wire vertical_tile_12_30_to_tile_11_30_3;

	wire vertical_tile_11_31_to_tile_12_31_0;
	wire vertical_tile_11_31_to_tile_12_31_1;
	wire vertical_tile_11_31_to_tile_12_31_2;
	wire vertical_tile_11_31_to_tile_12_31_3;
	wire vertical_tile_12_31_to_tile_11_31_0;
	wire vertical_tile_12_31_to_tile_11_31_1;
	wire vertical_tile_12_31_to_tile_11_31_2;
	wire vertical_tile_12_31_to_tile_11_31_3;

	wire vertical_tile_12_0_to_tile_13_0_0;
	wire vertical_tile_12_0_to_tile_13_0_1;
	wire vertical_tile_12_0_to_tile_13_0_2;
	wire vertical_tile_12_0_to_tile_13_0_3;
	wire vertical_tile_13_0_to_tile_12_0_0;
	wire vertical_tile_13_0_to_tile_12_0_1;
	wire vertical_tile_13_0_to_tile_12_0_2;
	wire vertical_tile_13_0_to_tile_12_0_3;

	wire vertical_tile_12_1_to_tile_13_1_0;
	wire vertical_tile_12_1_to_tile_13_1_1;
	wire vertical_tile_12_1_to_tile_13_1_2;
	wire vertical_tile_12_1_to_tile_13_1_3;
	wire vertical_tile_13_1_to_tile_12_1_0;
	wire vertical_tile_13_1_to_tile_12_1_1;
	wire vertical_tile_13_1_to_tile_12_1_2;
	wire vertical_tile_13_1_to_tile_12_1_3;

	wire vertical_tile_12_2_to_tile_13_2_0;
	wire vertical_tile_12_2_to_tile_13_2_1;
	wire vertical_tile_12_2_to_tile_13_2_2;
	wire vertical_tile_12_2_to_tile_13_2_3;
	wire vertical_tile_13_2_to_tile_12_2_0;
	wire vertical_tile_13_2_to_tile_12_2_1;
	wire vertical_tile_13_2_to_tile_12_2_2;
	wire vertical_tile_13_2_to_tile_12_2_3;

	wire vertical_tile_12_3_to_tile_13_3_0;
	wire vertical_tile_12_3_to_tile_13_3_1;
	wire vertical_tile_12_3_to_tile_13_3_2;
	wire vertical_tile_12_3_to_tile_13_3_3;
	wire vertical_tile_13_3_to_tile_12_3_0;
	wire vertical_tile_13_3_to_tile_12_3_1;
	wire vertical_tile_13_3_to_tile_12_3_2;
	wire vertical_tile_13_3_to_tile_12_3_3;

	wire vertical_tile_12_4_to_tile_13_4_0;
	wire vertical_tile_12_4_to_tile_13_4_1;
	wire vertical_tile_12_4_to_tile_13_4_2;
	wire vertical_tile_12_4_to_tile_13_4_3;
	wire vertical_tile_13_4_to_tile_12_4_0;
	wire vertical_tile_13_4_to_tile_12_4_1;
	wire vertical_tile_13_4_to_tile_12_4_2;
	wire vertical_tile_13_4_to_tile_12_4_3;

	wire vertical_tile_12_5_to_tile_13_5_0;
	wire vertical_tile_12_5_to_tile_13_5_1;
	wire vertical_tile_12_5_to_tile_13_5_2;
	wire vertical_tile_12_5_to_tile_13_5_3;
	wire vertical_tile_13_5_to_tile_12_5_0;
	wire vertical_tile_13_5_to_tile_12_5_1;
	wire vertical_tile_13_5_to_tile_12_5_2;
	wire vertical_tile_13_5_to_tile_12_5_3;

	wire vertical_tile_12_6_to_tile_13_6_0;
	wire vertical_tile_12_6_to_tile_13_6_1;
	wire vertical_tile_12_6_to_tile_13_6_2;
	wire vertical_tile_12_6_to_tile_13_6_3;
	wire vertical_tile_13_6_to_tile_12_6_0;
	wire vertical_tile_13_6_to_tile_12_6_1;
	wire vertical_tile_13_6_to_tile_12_6_2;
	wire vertical_tile_13_6_to_tile_12_6_3;

	wire vertical_tile_12_7_to_tile_13_7_0;
	wire vertical_tile_12_7_to_tile_13_7_1;
	wire vertical_tile_12_7_to_tile_13_7_2;
	wire vertical_tile_12_7_to_tile_13_7_3;
	wire vertical_tile_13_7_to_tile_12_7_0;
	wire vertical_tile_13_7_to_tile_12_7_1;
	wire vertical_tile_13_7_to_tile_12_7_2;
	wire vertical_tile_13_7_to_tile_12_7_3;

	wire vertical_tile_12_8_to_tile_13_8_0;
	wire vertical_tile_12_8_to_tile_13_8_1;
	wire vertical_tile_12_8_to_tile_13_8_2;
	wire vertical_tile_12_8_to_tile_13_8_3;
	wire vertical_tile_13_8_to_tile_12_8_0;
	wire vertical_tile_13_8_to_tile_12_8_1;
	wire vertical_tile_13_8_to_tile_12_8_2;
	wire vertical_tile_13_8_to_tile_12_8_3;

	wire vertical_tile_12_9_to_tile_13_9_0;
	wire vertical_tile_12_9_to_tile_13_9_1;
	wire vertical_tile_12_9_to_tile_13_9_2;
	wire vertical_tile_12_9_to_tile_13_9_3;
	wire vertical_tile_13_9_to_tile_12_9_0;
	wire vertical_tile_13_9_to_tile_12_9_1;
	wire vertical_tile_13_9_to_tile_12_9_2;
	wire vertical_tile_13_9_to_tile_12_9_3;

	wire vertical_tile_12_10_to_tile_13_10_0;
	wire vertical_tile_12_10_to_tile_13_10_1;
	wire vertical_tile_12_10_to_tile_13_10_2;
	wire vertical_tile_12_10_to_tile_13_10_3;
	wire vertical_tile_13_10_to_tile_12_10_0;
	wire vertical_tile_13_10_to_tile_12_10_1;
	wire vertical_tile_13_10_to_tile_12_10_2;
	wire vertical_tile_13_10_to_tile_12_10_3;

	wire vertical_tile_12_11_to_tile_13_11_0;
	wire vertical_tile_12_11_to_tile_13_11_1;
	wire vertical_tile_12_11_to_tile_13_11_2;
	wire vertical_tile_12_11_to_tile_13_11_3;
	wire vertical_tile_13_11_to_tile_12_11_0;
	wire vertical_tile_13_11_to_tile_12_11_1;
	wire vertical_tile_13_11_to_tile_12_11_2;
	wire vertical_tile_13_11_to_tile_12_11_3;

	wire vertical_tile_12_12_to_tile_13_12_0;
	wire vertical_tile_12_12_to_tile_13_12_1;
	wire vertical_tile_12_12_to_tile_13_12_2;
	wire vertical_tile_12_12_to_tile_13_12_3;
	wire vertical_tile_13_12_to_tile_12_12_0;
	wire vertical_tile_13_12_to_tile_12_12_1;
	wire vertical_tile_13_12_to_tile_12_12_2;
	wire vertical_tile_13_12_to_tile_12_12_3;

	wire vertical_tile_12_13_to_tile_13_13_0;
	wire vertical_tile_12_13_to_tile_13_13_1;
	wire vertical_tile_12_13_to_tile_13_13_2;
	wire vertical_tile_12_13_to_tile_13_13_3;
	wire vertical_tile_13_13_to_tile_12_13_0;
	wire vertical_tile_13_13_to_tile_12_13_1;
	wire vertical_tile_13_13_to_tile_12_13_2;
	wire vertical_tile_13_13_to_tile_12_13_3;

	wire vertical_tile_12_14_to_tile_13_14_0;
	wire vertical_tile_12_14_to_tile_13_14_1;
	wire vertical_tile_12_14_to_tile_13_14_2;
	wire vertical_tile_12_14_to_tile_13_14_3;
	wire vertical_tile_13_14_to_tile_12_14_0;
	wire vertical_tile_13_14_to_tile_12_14_1;
	wire vertical_tile_13_14_to_tile_12_14_2;
	wire vertical_tile_13_14_to_tile_12_14_3;

	wire vertical_tile_12_15_to_tile_13_15_0;
	wire vertical_tile_12_15_to_tile_13_15_1;
	wire vertical_tile_12_15_to_tile_13_15_2;
	wire vertical_tile_12_15_to_tile_13_15_3;
	wire vertical_tile_13_15_to_tile_12_15_0;
	wire vertical_tile_13_15_to_tile_12_15_1;
	wire vertical_tile_13_15_to_tile_12_15_2;
	wire vertical_tile_13_15_to_tile_12_15_3;

	wire vertical_tile_12_16_to_tile_13_16_0;
	wire vertical_tile_12_16_to_tile_13_16_1;
	wire vertical_tile_12_16_to_tile_13_16_2;
	wire vertical_tile_12_16_to_tile_13_16_3;
	wire vertical_tile_13_16_to_tile_12_16_0;
	wire vertical_tile_13_16_to_tile_12_16_1;
	wire vertical_tile_13_16_to_tile_12_16_2;
	wire vertical_tile_13_16_to_tile_12_16_3;

	wire vertical_tile_12_17_to_tile_13_17_0;
	wire vertical_tile_12_17_to_tile_13_17_1;
	wire vertical_tile_12_17_to_tile_13_17_2;
	wire vertical_tile_12_17_to_tile_13_17_3;
	wire vertical_tile_13_17_to_tile_12_17_0;
	wire vertical_tile_13_17_to_tile_12_17_1;
	wire vertical_tile_13_17_to_tile_12_17_2;
	wire vertical_tile_13_17_to_tile_12_17_3;

	wire vertical_tile_12_18_to_tile_13_18_0;
	wire vertical_tile_12_18_to_tile_13_18_1;
	wire vertical_tile_12_18_to_tile_13_18_2;
	wire vertical_tile_12_18_to_tile_13_18_3;
	wire vertical_tile_13_18_to_tile_12_18_0;
	wire vertical_tile_13_18_to_tile_12_18_1;
	wire vertical_tile_13_18_to_tile_12_18_2;
	wire vertical_tile_13_18_to_tile_12_18_3;

	wire vertical_tile_12_19_to_tile_13_19_0;
	wire vertical_tile_12_19_to_tile_13_19_1;
	wire vertical_tile_12_19_to_tile_13_19_2;
	wire vertical_tile_12_19_to_tile_13_19_3;
	wire vertical_tile_13_19_to_tile_12_19_0;
	wire vertical_tile_13_19_to_tile_12_19_1;
	wire vertical_tile_13_19_to_tile_12_19_2;
	wire vertical_tile_13_19_to_tile_12_19_3;

	wire vertical_tile_12_20_to_tile_13_20_0;
	wire vertical_tile_12_20_to_tile_13_20_1;
	wire vertical_tile_12_20_to_tile_13_20_2;
	wire vertical_tile_12_20_to_tile_13_20_3;
	wire vertical_tile_13_20_to_tile_12_20_0;
	wire vertical_tile_13_20_to_tile_12_20_1;
	wire vertical_tile_13_20_to_tile_12_20_2;
	wire vertical_tile_13_20_to_tile_12_20_3;

	wire vertical_tile_12_21_to_tile_13_21_0;
	wire vertical_tile_12_21_to_tile_13_21_1;
	wire vertical_tile_12_21_to_tile_13_21_2;
	wire vertical_tile_12_21_to_tile_13_21_3;
	wire vertical_tile_13_21_to_tile_12_21_0;
	wire vertical_tile_13_21_to_tile_12_21_1;
	wire vertical_tile_13_21_to_tile_12_21_2;
	wire vertical_tile_13_21_to_tile_12_21_3;

	wire vertical_tile_12_22_to_tile_13_22_0;
	wire vertical_tile_12_22_to_tile_13_22_1;
	wire vertical_tile_12_22_to_tile_13_22_2;
	wire vertical_tile_12_22_to_tile_13_22_3;
	wire vertical_tile_13_22_to_tile_12_22_0;
	wire vertical_tile_13_22_to_tile_12_22_1;
	wire vertical_tile_13_22_to_tile_12_22_2;
	wire vertical_tile_13_22_to_tile_12_22_3;

	wire vertical_tile_12_23_to_tile_13_23_0;
	wire vertical_tile_12_23_to_tile_13_23_1;
	wire vertical_tile_12_23_to_tile_13_23_2;
	wire vertical_tile_12_23_to_tile_13_23_3;
	wire vertical_tile_13_23_to_tile_12_23_0;
	wire vertical_tile_13_23_to_tile_12_23_1;
	wire vertical_tile_13_23_to_tile_12_23_2;
	wire vertical_tile_13_23_to_tile_12_23_3;

	wire vertical_tile_12_24_to_tile_13_24_0;
	wire vertical_tile_12_24_to_tile_13_24_1;
	wire vertical_tile_12_24_to_tile_13_24_2;
	wire vertical_tile_12_24_to_tile_13_24_3;
	wire vertical_tile_13_24_to_tile_12_24_0;
	wire vertical_tile_13_24_to_tile_12_24_1;
	wire vertical_tile_13_24_to_tile_12_24_2;
	wire vertical_tile_13_24_to_tile_12_24_3;

	wire vertical_tile_12_25_to_tile_13_25_0;
	wire vertical_tile_12_25_to_tile_13_25_1;
	wire vertical_tile_12_25_to_tile_13_25_2;
	wire vertical_tile_12_25_to_tile_13_25_3;
	wire vertical_tile_13_25_to_tile_12_25_0;
	wire vertical_tile_13_25_to_tile_12_25_1;
	wire vertical_tile_13_25_to_tile_12_25_2;
	wire vertical_tile_13_25_to_tile_12_25_3;

	wire vertical_tile_12_26_to_tile_13_26_0;
	wire vertical_tile_12_26_to_tile_13_26_1;
	wire vertical_tile_12_26_to_tile_13_26_2;
	wire vertical_tile_12_26_to_tile_13_26_3;
	wire vertical_tile_13_26_to_tile_12_26_0;
	wire vertical_tile_13_26_to_tile_12_26_1;
	wire vertical_tile_13_26_to_tile_12_26_2;
	wire vertical_tile_13_26_to_tile_12_26_3;

	wire vertical_tile_12_27_to_tile_13_27_0;
	wire vertical_tile_12_27_to_tile_13_27_1;
	wire vertical_tile_12_27_to_tile_13_27_2;
	wire vertical_tile_12_27_to_tile_13_27_3;
	wire vertical_tile_13_27_to_tile_12_27_0;
	wire vertical_tile_13_27_to_tile_12_27_1;
	wire vertical_tile_13_27_to_tile_12_27_2;
	wire vertical_tile_13_27_to_tile_12_27_3;

	wire vertical_tile_12_28_to_tile_13_28_0;
	wire vertical_tile_12_28_to_tile_13_28_1;
	wire vertical_tile_12_28_to_tile_13_28_2;
	wire vertical_tile_12_28_to_tile_13_28_3;
	wire vertical_tile_13_28_to_tile_12_28_0;
	wire vertical_tile_13_28_to_tile_12_28_1;
	wire vertical_tile_13_28_to_tile_12_28_2;
	wire vertical_tile_13_28_to_tile_12_28_3;

	wire vertical_tile_12_29_to_tile_13_29_0;
	wire vertical_tile_12_29_to_tile_13_29_1;
	wire vertical_tile_12_29_to_tile_13_29_2;
	wire vertical_tile_12_29_to_tile_13_29_3;
	wire vertical_tile_13_29_to_tile_12_29_0;
	wire vertical_tile_13_29_to_tile_12_29_1;
	wire vertical_tile_13_29_to_tile_12_29_2;
	wire vertical_tile_13_29_to_tile_12_29_3;

	wire vertical_tile_12_30_to_tile_13_30_0;
	wire vertical_tile_12_30_to_tile_13_30_1;
	wire vertical_tile_12_30_to_tile_13_30_2;
	wire vertical_tile_12_30_to_tile_13_30_3;
	wire vertical_tile_13_30_to_tile_12_30_0;
	wire vertical_tile_13_30_to_tile_12_30_1;
	wire vertical_tile_13_30_to_tile_12_30_2;
	wire vertical_tile_13_30_to_tile_12_30_3;

	wire vertical_tile_12_31_to_tile_13_31_0;
	wire vertical_tile_12_31_to_tile_13_31_1;
	wire vertical_tile_12_31_to_tile_13_31_2;
	wire vertical_tile_12_31_to_tile_13_31_3;
	wire vertical_tile_13_31_to_tile_12_31_0;
	wire vertical_tile_13_31_to_tile_12_31_1;
	wire vertical_tile_13_31_to_tile_12_31_2;
	wire vertical_tile_13_31_to_tile_12_31_3;

	wire vertical_tile_13_0_to_tile_14_0_0;
	wire vertical_tile_13_0_to_tile_14_0_1;
	wire vertical_tile_13_0_to_tile_14_0_2;
	wire vertical_tile_13_0_to_tile_14_0_3;
	wire vertical_tile_14_0_to_tile_13_0_0;
	wire vertical_tile_14_0_to_tile_13_0_1;
	wire vertical_tile_14_0_to_tile_13_0_2;
	wire vertical_tile_14_0_to_tile_13_0_3;

	wire vertical_tile_13_1_to_tile_14_1_0;
	wire vertical_tile_13_1_to_tile_14_1_1;
	wire vertical_tile_13_1_to_tile_14_1_2;
	wire vertical_tile_13_1_to_tile_14_1_3;
	wire vertical_tile_14_1_to_tile_13_1_0;
	wire vertical_tile_14_1_to_tile_13_1_1;
	wire vertical_tile_14_1_to_tile_13_1_2;
	wire vertical_tile_14_1_to_tile_13_1_3;

	wire vertical_tile_13_2_to_tile_14_2_0;
	wire vertical_tile_13_2_to_tile_14_2_1;
	wire vertical_tile_13_2_to_tile_14_2_2;
	wire vertical_tile_13_2_to_tile_14_2_3;
	wire vertical_tile_14_2_to_tile_13_2_0;
	wire vertical_tile_14_2_to_tile_13_2_1;
	wire vertical_tile_14_2_to_tile_13_2_2;
	wire vertical_tile_14_2_to_tile_13_2_3;

	wire vertical_tile_13_3_to_tile_14_3_0;
	wire vertical_tile_13_3_to_tile_14_3_1;
	wire vertical_tile_13_3_to_tile_14_3_2;
	wire vertical_tile_13_3_to_tile_14_3_3;
	wire vertical_tile_14_3_to_tile_13_3_0;
	wire vertical_tile_14_3_to_tile_13_3_1;
	wire vertical_tile_14_3_to_tile_13_3_2;
	wire vertical_tile_14_3_to_tile_13_3_3;

	wire vertical_tile_13_4_to_tile_14_4_0;
	wire vertical_tile_13_4_to_tile_14_4_1;
	wire vertical_tile_13_4_to_tile_14_4_2;
	wire vertical_tile_13_4_to_tile_14_4_3;
	wire vertical_tile_14_4_to_tile_13_4_0;
	wire vertical_tile_14_4_to_tile_13_4_1;
	wire vertical_tile_14_4_to_tile_13_4_2;
	wire vertical_tile_14_4_to_tile_13_4_3;

	wire vertical_tile_13_5_to_tile_14_5_0;
	wire vertical_tile_13_5_to_tile_14_5_1;
	wire vertical_tile_13_5_to_tile_14_5_2;
	wire vertical_tile_13_5_to_tile_14_5_3;
	wire vertical_tile_14_5_to_tile_13_5_0;
	wire vertical_tile_14_5_to_tile_13_5_1;
	wire vertical_tile_14_5_to_tile_13_5_2;
	wire vertical_tile_14_5_to_tile_13_5_3;

	wire vertical_tile_13_6_to_tile_14_6_0;
	wire vertical_tile_13_6_to_tile_14_6_1;
	wire vertical_tile_13_6_to_tile_14_6_2;
	wire vertical_tile_13_6_to_tile_14_6_3;
	wire vertical_tile_14_6_to_tile_13_6_0;
	wire vertical_tile_14_6_to_tile_13_6_1;
	wire vertical_tile_14_6_to_tile_13_6_2;
	wire vertical_tile_14_6_to_tile_13_6_3;

	wire vertical_tile_13_7_to_tile_14_7_0;
	wire vertical_tile_13_7_to_tile_14_7_1;
	wire vertical_tile_13_7_to_tile_14_7_2;
	wire vertical_tile_13_7_to_tile_14_7_3;
	wire vertical_tile_14_7_to_tile_13_7_0;
	wire vertical_tile_14_7_to_tile_13_7_1;
	wire vertical_tile_14_7_to_tile_13_7_2;
	wire vertical_tile_14_7_to_tile_13_7_3;

	wire vertical_tile_13_8_to_tile_14_8_0;
	wire vertical_tile_13_8_to_tile_14_8_1;
	wire vertical_tile_13_8_to_tile_14_8_2;
	wire vertical_tile_13_8_to_tile_14_8_3;
	wire vertical_tile_14_8_to_tile_13_8_0;
	wire vertical_tile_14_8_to_tile_13_8_1;
	wire vertical_tile_14_8_to_tile_13_8_2;
	wire vertical_tile_14_8_to_tile_13_8_3;

	wire vertical_tile_13_9_to_tile_14_9_0;
	wire vertical_tile_13_9_to_tile_14_9_1;
	wire vertical_tile_13_9_to_tile_14_9_2;
	wire vertical_tile_13_9_to_tile_14_9_3;
	wire vertical_tile_14_9_to_tile_13_9_0;
	wire vertical_tile_14_9_to_tile_13_9_1;
	wire vertical_tile_14_9_to_tile_13_9_2;
	wire vertical_tile_14_9_to_tile_13_9_3;

	wire vertical_tile_13_10_to_tile_14_10_0;
	wire vertical_tile_13_10_to_tile_14_10_1;
	wire vertical_tile_13_10_to_tile_14_10_2;
	wire vertical_tile_13_10_to_tile_14_10_3;
	wire vertical_tile_14_10_to_tile_13_10_0;
	wire vertical_tile_14_10_to_tile_13_10_1;
	wire vertical_tile_14_10_to_tile_13_10_2;
	wire vertical_tile_14_10_to_tile_13_10_3;

	wire vertical_tile_13_11_to_tile_14_11_0;
	wire vertical_tile_13_11_to_tile_14_11_1;
	wire vertical_tile_13_11_to_tile_14_11_2;
	wire vertical_tile_13_11_to_tile_14_11_3;
	wire vertical_tile_14_11_to_tile_13_11_0;
	wire vertical_tile_14_11_to_tile_13_11_1;
	wire vertical_tile_14_11_to_tile_13_11_2;
	wire vertical_tile_14_11_to_tile_13_11_3;

	wire vertical_tile_13_12_to_tile_14_12_0;
	wire vertical_tile_13_12_to_tile_14_12_1;
	wire vertical_tile_13_12_to_tile_14_12_2;
	wire vertical_tile_13_12_to_tile_14_12_3;
	wire vertical_tile_14_12_to_tile_13_12_0;
	wire vertical_tile_14_12_to_tile_13_12_1;
	wire vertical_tile_14_12_to_tile_13_12_2;
	wire vertical_tile_14_12_to_tile_13_12_3;

	wire vertical_tile_13_13_to_tile_14_13_0;
	wire vertical_tile_13_13_to_tile_14_13_1;
	wire vertical_tile_13_13_to_tile_14_13_2;
	wire vertical_tile_13_13_to_tile_14_13_3;
	wire vertical_tile_14_13_to_tile_13_13_0;
	wire vertical_tile_14_13_to_tile_13_13_1;
	wire vertical_tile_14_13_to_tile_13_13_2;
	wire vertical_tile_14_13_to_tile_13_13_3;

	wire vertical_tile_13_14_to_tile_14_14_0;
	wire vertical_tile_13_14_to_tile_14_14_1;
	wire vertical_tile_13_14_to_tile_14_14_2;
	wire vertical_tile_13_14_to_tile_14_14_3;
	wire vertical_tile_14_14_to_tile_13_14_0;
	wire vertical_tile_14_14_to_tile_13_14_1;
	wire vertical_tile_14_14_to_tile_13_14_2;
	wire vertical_tile_14_14_to_tile_13_14_3;

	wire vertical_tile_13_15_to_tile_14_15_0;
	wire vertical_tile_13_15_to_tile_14_15_1;
	wire vertical_tile_13_15_to_tile_14_15_2;
	wire vertical_tile_13_15_to_tile_14_15_3;
	wire vertical_tile_14_15_to_tile_13_15_0;
	wire vertical_tile_14_15_to_tile_13_15_1;
	wire vertical_tile_14_15_to_tile_13_15_2;
	wire vertical_tile_14_15_to_tile_13_15_3;

	wire vertical_tile_13_16_to_tile_14_16_0;
	wire vertical_tile_13_16_to_tile_14_16_1;
	wire vertical_tile_13_16_to_tile_14_16_2;
	wire vertical_tile_13_16_to_tile_14_16_3;
	wire vertical_tile_14_16_to_tile_13_16_0;
	wire vertical_tile_14_16_to_tile_13_16_1;
	wire vertical_tile_14_16_to_tile_13_16_2;
	wire vertical_tile_14_16_to_tile_13_16_3;

	wire vertical_tile_13_17_to_tile_14_17_0;
	wire vertical_tile_13_17_to_tile_14_17_1;
	wire vertical_tile_13_17_to_tile_14_17_2;
	wire vertical_tile_13_17_to_tile_14_17_3;
	wire vertical_tile_14_17_to_tile_13_17_0;
	wire vertical_tile_14_17_to_tile_13_17_1;
	wire vertical_tile_14_17_to_tile_13_17_2;
	wire vertical_tile_14_17_to_tile_13_17_3;

	wire vertical_tile_13_18_to_tile_14_18_0;
	wire vertical_tile_13_18_to_tile_14_18_1;
	wire vertical_tile_13_18_to_tile_14_18_2;
	wire vertical_tile_13_18_to_tile_14_18_3;
	wire vertical_tile_14_18_to_tile_13_18_0;
	wire vertical_tile_14_18_to_tile_13_18_1;
	wire vertical_tile_14_18_to_tile_13_18_2;
	wire vertical_tile_14_18_to_tile_13_18_3;

	wire vertical_tile_13_19_to_tile_14_19_0;
	wire vertical_tile_13_19_to_tile_14_19_1;
	wire vertical_tile_13_19_to_tile_14_19_2;
	wire vertical_tile_13_19_to_tile_14_19_3;
	wire vertical_tile_14_19_to_tile_13_19_0;
	wire vertical_tile_14_19_to_tile_13_19_1;
	wire vertical_tile_14_19_to_tile_13_19_2;
	wire vertical_tile_14_19_to_tile_13_19_3;

	wire vertical_tile_13_20_to_tile_14_20_0;
	wire vertical_tile_13_20_to_tile_14_20_1;
	wire vertical_tile_13_20_to_tile_14_20_2;
	wire vertical_tile_13_20_to_tile_14_20_3;
	wire vertical_tile_14_20_to_tile_13_20_0;
	wire vertical_tile_14_20_to_tile_13_20_1;
	wire vertical_tile_14_20_to_tile_13_20_2;
	wire vertical_tile_14_20_to_tile_13_20_3;

	wire vertical_tile_13_21_to_tile_14_21_0;
	wire vertical_tile_13_21_to_tile_14_21_1;
	wire vertical_tile_13_21_to_tile_14_21_2;
	wire vertical_tile_13_21_to_tile_14_21_3;
	wire vertical_tile_14_21_to_tile_13_21_0;
	wire vertical_tile_14_21_to_tile_13_21_1;
	wire vertical_tile_14_21_to_tile_13_21_2;
	wire vertical_tile_14_21_to_tile_13_21_3;

	wire vertical_tile_13_22_to_tile_14_22_0;
	wire vertical_tile_13_22_to_tile_14_22_1;
	wire vertical_tile_13_22_to_tile_14_22_2;
	wire vertical_tile_13_22_to_tile_14_22_3;
	wire vertical_tile_14_22_to_tile_13_22_0;
	wire vertical_tile_14_22_to_tile_13_22_1;
	wire vertical_tile_14_22_to_tile_13_22_2;
	wire vertical_tile_14_22_to_tile_13_22_3;

	wire vertical_tile_13_23_to_tile_14_23_0;
	wire vertical_tile_13_23_to_tile_14_23_1;
	wire vertical_tile_13_23_to_tile_14_23_2;
	wire vertical_tile_13_23_to_tile_14_23_3;
	wire vertical_tile_14_23_to_tile_13_23_0;
	wire vertical_tile_14_23_to_tile_13_23_1;
	wire vertical_tile_14_23_to_tile_13_23_2;
	wire vertical_tile_14_23_to_tile_13_23_3;

	wire vertical_tile_13_24_to_tile_14_24_0;
	wire vertical_tile_13_24_to_tile_14_24_1;
	wire vertical_tile_13_24_to_tile_14_24_2;
	wire vertical_tile_13_24_to_tile_14_24_3;
	wire vertical_tile_14_24_to_tile_13_24_0;
	wire vertical_tile_14_24_to_tile_13_24_1;
	wire vertical_tile_14_24_to_tile_13_24_2;
	wire vertical_tile_14_24_to_tile_13_24_3;

	wire vertical_tile_13_25_to_tile_14_25_0;
	wire vertical_tile_13_25_to_tile_14_25_1;
	wire vertical_tile_13_25_to_tile_14_25_2;
	wire vertical_tile_13_25_to_tile_14_25_3;
	wire vertical_tile_14_25_to_tile_13_25_0;
	wire vertical_tile_14_25_to_tile_13_25_1;
	wire vertical_tile_14_25_to_tile_13_25_2;
	wire vertical_tile_14_25_to_tile_13_25_3;

	wire vertical_tile_13_26_to_tile_14_26_0;
	wire vertical_tile_13_26_to_tile_14_26_1;
	wire vertical_tile_13_26_to_tile_14_26_2;
	wire vertical_tile_13_26_to_tile_14_26_3;
	wire vertical_tile_14_26_to_tile_13_26_0;
	wire vertical_tile_14_26_to_tile_13_26_1;
	wire vertical_tile_14_26_to_tile_13_26_2;
	wire vertical_tile_14_26_to_tile_13_26_3;

	wire vertical_tile_13_27_to_tile_14_27_0;
	wire vertical_tile_13_27_to_tile_14_27_1;
	wire vertical_tile_13_27_to_tile_14_27_2;
	wire vertical_tile_13_27_to_tile_14_27_3;
	wire vertical_tile_14_27_to_tile_13_27_0;
	wire vertical_tile_14_27_to_tile_13_27_1;
	wire vertical_tile_14_27_to_tile_13_27_2;
	wire vertical_tile_14_27_to_tile_13_27_3;

	wire vertical_tile_13_28_to_tile_14_28_0;
	wire vertical_tile_13_28_to_tile_14_28_1;
	wire vertical_tile_13_28_to_tile_14_28_2;
	wire vertical_tile_13_28_to_tile_14_28_3;
	wire vertical_tile_14_28_to_tile_13_28_0;
	wire vertical_tile_14_28_to_tile_13_28_1;
	wire vertical_tile_14_28_to_tile_13_28_2;
	wire vertical_tile_14_28_to_tile_13_28_3;

	wire vertical_tile_13_29_to_tile_14_29_0;
	wire vertical_tile_13_29_to_tile_14_29_1;
	wire vertical_tile_13_29_to_tile_14_29_2;
	wire vertical_tile_13_29_to_tile_14_29_3;
	wire vertical_tile_14_29_to_tile_13_29_0;
	wire vertical_tile_14_29_to_tile_13_29_1;
	wire vertical_tile_14_29_to_tile_13_29_2;
	wire vertical_tile_14_29_to_tile_13_29_3;

	wire vertical_tile_13_30_to_tile_14_30_0;
	wire vertical_tile_13_30_to_tile_14_30_1;
	wire vertical_tile_13_30_to_tile_14_30_2;
	wire vertical_tile_13_30_to_tile_14_30_3;
	wire vertical_tile_14_30_to_tile_13_30_0;
	wire vertical_tile_14_30_to_tile_13_30_1;
	wire vertical_tile_14_30_to_tile_13_30_2;
	wire vertical_tile_14_30_to_tile_13_30_3;

	wire vertical_tile_13_31_to_tile_14_31_0;
	wire vertical_tile_13_31_to_tile_14_31_1;
	wire vertical_tile_13_31_to_tile_14_31_2;
	wire vertical_tile_13_31_to_tile_14_31_3;
	wire vertical_tile_14_31_to_tile_13_31_0;
	wire vertical_tile_14_31_to_tile_13_31_1;
	wire vertical_tile_14_31_to_tile_13_31_2;
	wire vertical_tile_14_31_to_tile_13_31_3;

	wire vertical_tile_14_0_to_tile_15_0_0;
	wire vertical_tile_14_0_to_tile_15_0_1;
	wire vertical_tile_14_0_to_tile_15_0_2;
	wire vertical_tile_14_0_to_tile_15_0_3;
	wire vertical_tile_15_0_to_tile_14_0_0;
	wire vertical_tile_15_0_to_tile_14_0_1;
	wire vertical_tile_15_0_to_tile_14_0_2;
	wire vertical_tile_15_0_to_tile_14_0_3;

	wire vertical_tile_14_1_to_tile_15_1_0;
	wire vertical_tile_14_1_to_tile_15_1_1;
	wire vertical_tile_14_1_to_tile_15_1_2;
	wire vertical_tile_14_1_to_tile_15_1_3;
	wire vertical_tile_15_1_to_tile_14_1_0;
	wire vertical_tile_15_1_to_tile_14_1_1;
	wire vertical_tile_15_1_to_tile_14_1_2;
	wire vertical_tile_15_1_to_tile_14_1_3;

	wire vertical_tile_14_2_to_tile_15_2_0;
	wire vertical_tile_14_2_to_tile_15_2_1;
	wire vertical_tile_14_2_to_tile_15_2_2;
	wire vertical_tile_14_2_to_tile_15_2_3;
	wire vertical_tile_15_2_to_tile_14_2_0;
	wire vertical_tile_15_2_to_tile_14_2_1;
	wire vertical_tile_15_2_to_tile_14_2_2;
	wire vertical_tile_15_2_to_tile_14_2_3;

	wire vertical_tile_14_3_to_tile_15_3_0;
	wire vertical_tile_14_3_to_tile_15_3_1;
	wire vertical_tile_14_3_to_tile_15_3_2;
	wire vertical_tile_14_3_to_tile_15_3_3;
	wire vertical_tile_15_3_to_tile_14_3_0;
	wire vertical_tile_15_3_to_tile_14_3_1;
	wire vertical_tile_15_3_to_tile_14_3_2;
	wire vertical_tile_15_3_to_tile_14_3_3;

	wire vertical_tile_14_4_to_tile_15_4_0;
	wire vertical_tile_14_4_to_tile_15_4_1;
	wire vertical_tile_14_4_to_tile_15_4_2;
	wire vertical_tile_14_4_to_tile_15_4_3;
	wire vertical_tile_15_4_to_tile_14_4_0;
	wire vertical_tile_15_4_to_tile_14_4_1;
	wire vertical_tile_15_4_to_tile_14_4_2;
	wire vertical_tile_15_4_to_tile_14_4_3;

	wire vertical_tile_14_5_to_tile_15_5_0;
	wire vertical_tile_14_5_to_tile_15_5_1;
	wire vertical_tile_14_5_to_tile_15_5_2;
	wire vertical_tile_14_5_to_tile_15_5_3;
	wire vertical_tile_15_5_to_tile_14_5_0;
	wire vertical_tile_15_5_to_tile_14_5_1;
	wire vertical_tile_15_5_to_tile_14_5_2;
	wire vertical_tile_15_5_to_tile_14_5_3;

	wire vertical_tile_14_6_to_tile_15_6_0;
	wire vertical_tile_14_6_to_tile_15_6_1;
	wire vertical_tile_14_6_to_tile_15_6_2;
	wire vertical_tile_14_6_to_tile_15_6_3;
	wire vertical_tile_15_6_to_tile_14_6_0;
	wire vertical_tile_15_6_to_tile_14_6_1;
	wire vertical_tile_15_6_to_tile_14_6_2;
	wire vertical_tile_15_6_to_tile_14_6_3;

	wire vertical_tile_14_7_to_tile_15_7_0;
	wire vertical_tile_14_7_to_tile_15_7_1;
	wire vertical_tile_14_7_to_tile_15_7_2;
	wire vertical_tile_14_7_to_tile_15_7_3;
	wire vertical_tile_15_7_to_tile_14_7_0;
	wire vertical_tile_15_7_to_tile_14_7_1;
	wire vertical_tile_15_7_to_tile_14_7_2;
	wire vertical_tile_15_7_to_tile_14_7_3;

	wire vertical_tile_14_8_to_tile_15_8_0;
	wire vertical_tile_14_8_to_tile_15_8_1;
	wire vertical_tile_14_8_to_tile_15_8_2;
	wire vertical_tile_14_8_to_tile_15_8_3;
	wire vertical_tile_15_8_to_tile_14_8_0;
	wire vertical_tile_15_8_to_tile_14_8_1;
	wire vertical_tile_15_8_to_tile_14_8_2;
	wire vertical_tile_15_8_to_tile_14_8_3;

	wire vertical_tile_14_9_to_tile_15_9_0;
	wire vertical_tile_14_9_to_tile_15_9_1;
	wire vertical_tile_14_9_to_tile_15_9_2;
	wire vertical_tile_14_9_to_tile_15_9_3;
	wire vertical_tile_15_9_to_tile_14_9_0;
	wire vertical_tile_15_9_to_tile_14_9_1;
	wire vertical_tile_15_9_to_tile_14_9_2;
	wire vertical_tile_15_9_to_tile_14_9_3;

	wire vertical_tile_14_10_to_tile_15_10_0;
	wire vertical_tile_14_10_to_tile_15_10_1;
	wire vertical_tile_14_10_to_tile_15_10_2;
	wire vertical_tile_14_10_to_tile_15_10_3;
	wire vertical_tile_15_10_to_tile_14_10_0;
	wire vertical_tile_15_10_to_tile_14_10_1;
	wire vertical_tile_15_10_to_tile_14_10_2;
	wire vertical_tile_15_10_to_tile_14_10_3;

	wire vertical_tile_14_11_to_tile_15_11_0;
	wire vertical_tile_14_11_to_tile_15_11_1;
	wire vertical_tile_14_11_to_tile_15_11_2;
	wire vertical_tile_14_11_to_tile_15_11_3;
	wire vertical_tile_15_11_to_tile_14_11_0;
	wire vertical_tile_15_11_to_tile_14_11_1;
	wire vertical_tile_15_11_to_tile_14_11_2;
	wire vertical_tile_15_11_to_tile_14_11_3;

	wire vertical_tile_14_12_to_tile_15_12_0;
	wire vertical_tile_14_12_to_tile_15_12_1;
	wire vertical_tile_14_12_to_tile_15_12_2;
	wire vertical_tile_14_12_to_tile_15_12_3;
	wire vertical_tile_15_12_to_tile_14_12_0;
	wire vertical_tile_15_12_to_tile_14_12_1;
	wire vertical_tile_15_12_to_tile_14_12_2;
	wire vertical_tile_15_12_to_tile_14_12_3;

	wire vertical_tile_14_13_to_tile_15_13_0;
	wire vertical_tile_14_13_to_tile_15_13_1;
	wire vertical_tile_14_13_to_tile_15_13_2;
	wire vertical_tile_14_13_to_tile_15_13_3;
	wire vertical_tile_15_13_to_tile_14_13_0;
	wire vertical_tile_15_13_to_tile_14_13_1;
	wire vertical_tile_15_13_to_tile_14_13_2;
	wire vertical_tile_15_13_to_tile_14_13_3;

	wire vertical_tile_14_14_to_tile_15_14_0;
	wire vertical_tile_14_14_to_tile_15_14_1;
	wire vertical_tile_14_14_to_tile_15_14_2;
	wire vertical_tile_14_14_to_tile_15_14_3;
	wire vertical_tile_15_14_to_tile_14_14_0;
	wire vertical_tile_15_14_to_tile_14_14_1;
	wire vertical_tile_15_14_to_tile_14_14_2;
	wire vertical_tile_15_14_to_tile_14_14_3;

	wire vertical_tile_14_15_to_tile_15_15_0;
	wire vertical_tile_14_15_to_tile_15_15_1;
	wire vertical_tile_14_15_to_tile_15_15_2;
	wire vertical_tile_14_15_to_tile_15_15_3;
	wire vertical_tile_15_15_to_tile_14_15_0;
	wire vertical_tile_15_15_to_tile_14_15_1;
	wire vertical_tile_15_15_to_tile_14_15_2;
	wire vertical_tile_15_15_to_tile_14_15_3;

	wire vertical_tile_14_16_to_tile_15_16_0;
	wire vertical_tile_14_16_to_tile_15_16_1;
	wire vertical_tile_14_16_to_tile_15_16_2;
	wire vertical_tile_14_16_to_tile_15_16_3;
	wire vertical_tile_15_16_to_tile_14_16_0;
	wire vertical_tile_15_16_to_tile_14_16_1;
	wire vertical_tile_15_16_to_tile_14_16_2;
	wire vertical_tile_15_16_to_tile_14_16_3;

	wire vertical_tile_14_17_to_tile_15_17_0;
	wire vertical_tile_14_17_to_tile_15_17_1;
	wire vertical_tile_14_17_to_tile_15_17_2;
	wire vertical_tile_14_17_to_tile_15_17_3;
	wire vertical_tile_15_17_to_tile_14_17_0;
	wire vertical_tile_15_17_to_tile_14_17_1;
	wire vertical_tile_15_17_to_tile_14_17_2;
	wire vertical_tile_15_17_to_tile_14_17_3;

	wire vertical_tile_14_18_to_tile_15_18_0;
	wire vertical_tile_14_18_to_tile_15_18_1;
	wire vertical_tile_14_18_to_tile_15_18_2;
	wire vertical_tile_14_18_to_tile_15_18_3;
	wire vertical_tile_15_18_to_tile_14_18_0;
	wire vertical_tile_15_18_to_tile_14_18_1;
	wire vertical_tile_15_18_to_tile_14_18_2;
	wire vertical_tile_15_18_to_tile_14_18_3;

	wire vertical_tile_14_19_to_tile_15_19_0;
	wire vertical_tile_14_19_to_tile_15_19_1;
	wire vertical_tile_14_19_to_tile_15_19_2;
	wire vertical_tile_14_19_to_tile_15_19_3;
	wire vertical_tile_15_19_to_tile_14_19_0;
	wire vertical_tile_15_19_to_tile_14_19_1;
	wire vertical_tile_15_19_to_tile_14_19_2;
	wire vertical_tile_15_19_to_tile_14_19_3;

	wire vertical_tile_14_20_to_tile_15_20_0;
	wire vertical_tile_14_20_to_tile_15_20_1;
	wire vertical_tile_14_20_to_tile_15_20_2;
	wire vertical_tile_14_20_to_tile_15_20_3;
	wire vertical_tile_15_20_to_tile_14_20_0;
	wire vertical_tile_15_20_to_tile_14_20_1;
	wire vertical_tile_15_20_to_tile_14_20_2;
	wire vertical_tile_15_20_to_tile_14_20_3;

	wire vertical_tile_14_21_to_tile_15_21_0;
	wire vertical_tile_14_21_to_tile_15_21_1;
	wire vertical_tile_14_21_to_tile_15_21_2;
	wire vertical_tile_14_21_to_tile_15_21_3;
	wire vertical_tile_15_21_to_tile_14_21_0;
	wire vertical_tile_15_21_to_tile_14_21_1;
	wire vertical_tile_15_21_to_tile_14_21_2;
	wire vertical_tile_15_21_to_tile_14_21_3;

	wire vertical_tile_14_22_to_tile_15_22_0;
	wire vertical_tile_14_22_to_tile_15_22_1;
	wire vertical_tile_14_22_to_tile_15_22_2;
	wire vertical_tile_14_22_to_tile_15_22_3;
	wire vertical_tile_15_22_to_tile_14_22_0;
	wire vertical_tile_15_22_to_tile_14_22_1;
	wire vertical_tile_15_22_to_tile_14_22_2;
	wire vertical_tile_15_22_to_tile_14_22_3;

	wire vertical_tile_14_23_to_tile_15_23_0;
	wire vertical_tile_14_23_to_tile_15_23_1;
	wire vertical_tile_14_23_to_tile_15_23_2;
	wire vertical_tile_14_23_to_tile_15_23_3;
	wire vertical_tile_15_23_to_tile_14_23_0;
	wire vertical_tile_15_23_to_tile_14_23_1;
	wire vertical_tile_15_23_to_tile_14_23_2;
	wire vertical_tile_15_23_to_tile_14_23_3;

	wire vertical_tile_14_24_to_tile_15_24_0;
	wire vertical_tile_14_24_to_tile_15_24_1;
	wire vertical_tile_14_24_to_tile_15_24_2;
	wire vertical_tile_14_24_to_tile_15_24_3;
	wire vertical_tile_15_24_to_tile_14_24_0;
	wire vertical_tile_15_24_to_tile_14_24_1;
	wire vertical_tile_15_24_to_tile_14_24_2;
	wire vertical_tile_15_24_to_tile_14_24_3;

	wire vertical_tile_14_25_to_tile_15_25_0;
	wire vertical_tile_14_25_to_tile_15_25_1;
	wire vertical_tile_14_25_to_tile_15_25_2;
	wire vertical_tile_14_25_to_tile_15_25_3;
	wire vertical_tile_15_25_to_tile_14_25_0;
	wire vertical_tile_15_25_to_tile_14_25_1;
	wire vertical_tile_15_25_to_tile_14_25_2;
	wire vertical_tile_15_25_to_tile_14_25_3;

	wire vertical_tile_14_26_to_tile_15_26_0;
	wire vertical_tile_14_26_to_tile_15_26_1;
	wire vertical_tile_14_26_to_tile_15_26_2;
	wire vertical_tile_14_26_to_tile_15_26_3;
	wire vertical_tile_15_26_to_tile_14_26_0;
	wire vertical_tile_15_26_to_tile_14_26_1;
	wire vertical_tile_15_26_to_tile_14_26_2;
	wire vertical_tile_15_26_to_tile_14_26_3;

	wire vertical_tile_14_27_to_tile_15_27_0;
	wire vertical_tile_14_27_to_tile_15_27_1;
	wire vertical_tile_14_27_to_tile_15_27_2;
	wire vertical_tile_14_27_to_tile_15_27_3;
	wire vertical_tile_15_27_to_tile_14_27_0;
	wire vertical_tile_15_27_to_tile_14_27_1;
	wire vertical_tile_15_27_to_tile_14_27_2;
	wire vertical_tile_15_27_to_tile_14_27_3;

	wire vertical_tile_14_28_to_tile_15_28_0;
	wire vertical_tile_14_28_to_tile_15_28_1;
	wire vertical_tile_14_28_to_tile_15_28_2;
	wire vertical_tile_14_28_to_tile_15_28_3;
	wire vertical_tile_15_28_to_tile_14_28_0;
	wire vertical_tile_15_28_to_tile_14_28_1;
	wire vertical_tile_15_28_to_tile_14_28_2;
	wire vertical_tile_15_28_to_tile_14_28_3;

	wire vertical_tile_14_29_to_tile_15_29_0;
	wire vertical_tile_14_29_to_tile_15_29_1;
	wire vertical_tile_14_29_to_tile_15_29_2;
	wire vertical_tile_14_29_to_tile_15_29_3;
	wire vertical_tile_15_29_to_tile_14_29_0;
	wire vertical_tile_15_29_to_tile_14_29_1;
	wire vertical_tile_15_29_to_tile_14_29_2;
	wire vertical_tile_15_29_to_tile_14_29_3;

	wire vertical_tile_14_30_to_tile_15_30_0;
	wire vertical_tile_14_30_to_tile_15_30_1;
	wire vertical_tile_14_30_to_tile_15_30_2;
	wire vertical_tile_14_30_to_tile_15_30_3;
	wire vertical_tile_15_30_to_tile_14_30_0;
	wire vertical_tile_15_30_to_tile_14_30_1;
	wire vertical_tile_15_30_to_tile_14_30_2;
	wire vertical_tile_15_30_to_tile_14_30_3;

	wire vertical_tile_14_31_to_tile_15_31_0;
	wire vertical_tile_14_31_to_tile_15_31_1;
	wire vertical_tile_14_31_to_tile_15_31_2;
	wire vertical_tile_14_31_to_tile_15_31_3;
	wire vertical_tile_15_31_to_tile_14_31_0;
	wire vertical_tile_15_31_to_tile_14_31_1;
	wire vertical_tile_15_31_to_tile_14_31_2;
	wire vertical_tile_15_31_to_tile_14_31_3;

	wire vertical_tile_15_0_to_tile_16_0_0;
	wire vertical_tile_15_0_to_tile_16_0_1;
	wire vertical_tile_15_0_to_tile_16_0_2;
	wire vertical_tile_15_0_to_tile_16_0_3;
	wire vertical_tile_16_0_to_tile_15_0_0;
	wire vertical_tile_16_0_to_tile_15_0_1;
	wire vertical_tile_16_0_to_tile_15_0_2;
	wire vertical_tile_16_0_to_tile_15_0_3;

	wire vertical_tile_15_1_to_tile_16_1_0;
	wire vertical_tile_15_1_to_tile_16_1_1;
	wire vertical_tile_15_1_to_tile_16_1_2;
	wire vertical_tile_15_1_to_tile_16_1_3;
	wire vertical_tile_16_1_to_tile_15_1_0;
	wire vertical_tile_16_1_to_tile_15_1_1;
	wire vertical_tile_16_1_to_tile_15_1_2;
	wire vertical_tile_16_1_to_tile_15_1_3;

	wire vertical_tile_15_2_to_tile_16_2_0;
	wire vertical_tile_15_2_to_tile_16_2_1;
	wire vertical_tile_15_2_to_tile_16_2_2;
	wire vertical_tile_15_2_to_tile_16_2_3;
	wire vertical_tile_16_2_to_tile_15_2_0;
	wire vertical_tile_16_2_to_tile_15_2_1;
	wire vertical_tile_16_2_to_tile_15_2_2;
	wire vertical_tile_16_2_to_tile_15_2_3;

	wire vertical_tile_15_3_to_tile_16_3_0;
	wire vertical_tile_15_3_to_tile_16_3_1;
	wire vertical_tile_15_3_to_tile_16_3_2;
	wire vertical_tile_15_3_to_tile_16_3_3;
	wire vertical_tile_16_3_to_tile_15_3_0;
	wire vertical_tile_16_3_to_tile_15_3_1;
	wire vertical_tile_16_3_to_tile_15_3_2;
	wire vertical_tile_16_3_to_tile_15_3_3;

	wire vertical_tile_15_4_to_tile_16_4_0;
	wire vertical_tile_15_4_to_tile_16_4_1;
	wire vertical_tile_15_4_to_tile_16_4_2;
	wire vertical_tile_15_4_to_tile_16_4_3;
	wire vertical_tile_16_4_to_tile_15_4_0;
	wire vertical_tile_16_4_to_tile_15_4_1;
	wire vertical_tile_16_4_to_tile_15_4_2;
	wire vertical_tile_16_4_to_tile_15_4_3;

	wire vertical_tile_15_5_to_tile_16_5_0;
	wire vertical_tile_15_5_to_tile_16_5_1;
	wire vertical_tile_15_5_to_tile_16_5_2;
	wire vertical_tile_15_5_to_tile_16_5_3;
	wire vertical_tile_16_5_to_tile_15_5_0;
	wire vertical_tile_16_5_to_tile_15_5_1;
	wire vertical_tile_16_5_to_tile_15_5_2;
	wire vertical_tile_16_5_to_tile_15_5_3;

	wire vertical_tile_15_6_to_tile_16_6_0;
	wire vertical_tile_15_6_to_tile_16_6_1;
	wire vertical_tile_15_6_to_tile_16_6_2;
	wire vertical_tile_15_6_to_tile_16_6_3;
	wire vertical_tile_16_6_to_tile_15_6_0;
	wire vertical_tile_16_6_to_tile_15_6_1;
	wire vertical_tile_16_6_to_tile_15_6_2;
	wire vertical_tile_16_6_to_tile_15_6_3;

	wire vertical_tile_15_7_to_tile_16_7_0;
	wire vertical_tile_15_7_to_tile_16_7_1;
	wire vertical_tile_15_7_to_tile_16_7_2;
	wire vertical_tile_15_7_to_tile_16_7_3;
	wire vertical_tile_16_7_to_tile_15_7_0;
	wire vertical_tile_16_7_to_tile_15_7_1;
	wire vertical_tile_16_7_to_tile_15_7_2;
	wire vertical_tile_16_7_to_tile_15_7_3;

	wire vertical_tile_15_8_to_tile_16_8_0;
	wire vertical_tile_15_8_to_tile_16_8_1;
	wire vertical_tile_15_8_to_tile_16_8_2;
	wire vertical_tile_15_8_to_tile_16_8_3;
	wire vertical_tile_16_8_to_tile_15_8_0;
	wire vertical_tile_16_8_to_tile_15_8_1;
	wire vertical_tile_16_8_to_tile_15_8_2;
	wire vertical_tile_16_8_to_tile_15_8_3;

	wire vertical_tile_15_9_to_tile_16_9_0;
	wire vertical_tile_15_9_to_tile_16_9_1;
	wire vertical_tile_15_9_to_tile_16_9_2;
	wire vertical_tile_15_9_to_tile_16_9_3;
	wire vertical_tile_16_9_to_tile_15_9_0;
	wire vertical_tile_16_9_to_tile_15_9_1;
	wire vertical_tile_16_9_to_tile_15_9_2;
	wire vertical_tile_16_9_to_tile_15_9_3;

	wire vertical_tile_15_10_to_tile_16_10_0;
	wire vertical_tile_15_10_to_tile_16_10_1;
	wire vertical_tile_15_10_to_tile_16_10_2;
	wire vertical_tile_15_10_to_tile_16_10_3;
	wire vertical_tile_16_10_to_tile_15_10_0;
	wire vertical_tile_16_10_to_tile_15_10_1;
	wire vertical_tile_16_10_to_tile_15_10_2;
	wire vertical_tile_16_10_to_tile_15_10_3;

	wire vertical_tile_15_11_to_tile_16_11_0;
	wire vertical_tile_15_11_to_tile_16_11_1;
	wire vertical_tile_15_11_to_tile_16_11_2;
	wire vertical_tile_15_11_to_tile_16_11_3;
	wire vertical_tile_16_11_to_tile_15_11_0;
	wire vertical_tile_16_11_to_tile_15_11_1;
	wire vertical_tile_16_11_to_tile_15_11_2;
	wire vertical_tile_16_11_to_tile_15_11_3;

	wire vertical_tile_15_12_to_tile_16_12_0;
	wire vertical_tile_15_12_to_tile_16_12_1;
	wire vertical_tile_15_12_to_tile_16_12_2;
	wire vertical_tile_15_12_to_tile_16_12_3;
	wire vertical_tile_16_12_to_tile_15_12_0;
	wire vertical_tile_16_12_to_tile_15_12_1;
	wire vertical_tile_16_12_to_tile_15_12_2;
	wire vertical_tile_16_12_to_tile_15_12_3;

	wire vertical_tile_15_13_to_tile_16_13_0;
	wire vertical_tile_15_13_to_tile_16_13_1;
	wire vertical_tile_15_13_to_tile_16_13_2;
	wire vertical_tile_15_13_to_tile_16_13_3;
	wire vertical_tile_16_13_to_tile_15_13_0;
	wire vertical_tile_16_13_to_tile_15_13_1;
	wire vertical_tile_16_13_to_tile_15_13_2;
	wire vertical_tile_16_13_to_tile_15_13_3;

	wire vertical_tile_15_14_to_tile_16_14_0;
	wire vertical_tile_15_14_to_tile_16_14_1;
	wire vertical_tile_15_14_to_tile_16_14_2;
	wire vertical_tile_15_14_to_tile_16_14_3;
	wire vertical_tile_16_14_to_tile_15_14_0;
	wire vertical_tile_16_14_to_tile_15_14_1;
	wire vertical_tile_16_14_to_tile_15_14_2;
	wire vertical_tile_16_14_to_tile_15_14_3;

	wire vertical_tile_15_15_to_tile_16_15_0;
	wire vertical_tile_15_15_to_tile_16_15_1;
	wire vertical_tile_15_15_to_tile_16_15_2;
	wire vertical_tile_15_15_to_tile_16_15_3;
	wire vertical_tile_16_15_to_tile_15_15_0;
	wire vertical_tile_16_15_to_tile_15_15_1;
	wire vertical_tile_16_15_to_tile_15_15_2;
	wire vertical_tile_16_15_to_tile_15_15_3;

	wire vertical_tile_15_16_to_tile_16_16_0;
	wire vertical_tile_15_16_to_tile_16_16_1;
	wire vertical_tile_15_16_to_tile_16_16_2;
	wire vertical_tile_15_16_to_tile_16_16_3;
	wire vertical_tile_16_16_to_tile_15_16_0;
	wire vertical_tile_16_16_to_tile_15_16_1;
	wire vertical_tile_16_16_to_tile_15_16_2;
	wire vertical_tile_16_16_to_tile_15_16_3;

	wire vertical_tile_15_17_to_tile_16_17_0;
	wire vertical_tile_15_17_to_tile_16_17_1;
	wire vertical_tile_15_17_to_tile_16_17_2;
	wire vertical_tile_15_17_to_tile_16_17_3;
	wire vertical_tile_16_17_to_tile_15_17_0;
	wire vertical_tile_16_17_to_tile_15_17_1;
	wire vertical_tile_16_17_to_tile_15_17_2;
	wire vertical_tile_16_17_to_tile_15_17_3;

	wire vertical_tile_15_18_to_tile_16_18_0;
	wire vertical_tile_15_18_to_tile_16_18_1;
	wire vertical_tile_15_18_to_tile_16_18_2;
	wire vertical_tile_15_18_to_tile_16_18_3;
	wire vertical_tile_16_18_to_tile_15_18_0;
	wire vertical_tile_16_18_to_tile_15_18_1;
	wire vertical_tile_16_18_to_tile_15_18_2;
	wire vertical_tile_16_18_to_tile_15_18_3;

	wire vertical_tile_15_19_to_tile_16_19_0;
	wire vertical_tile_15_19_to_tile_16_19_1;
	wire vertical_tile_15_19_to_tile_16_19_2;
	wire vertical_tile_15_19_to_tile_16_19_3;
	wire vertical_tile_16_19_to_tile_15_19_0;
	wire vertical_tile_16_19_to_tile_15_19_1;
	wire vertical_tile_16_19_to_tile_15_19_2;
	wire vertical_tile_16_19_to_tile_15_19_3;

	wire vertical_tile_15_20_to_tile_16_20_0;
	wire vertical_tile_15_20_to_tile_16_20_1;
	wire vertical_tile_15_20_to_tile_16_20_2;
	wire vertical_tile_15_20_to_tile_16_20_3;
	wire vertical_tile_16_20_to_tile_15_20_0;
	wire vertical_tile_16_20_to_tile_15_20_1;
	wire vertical_tile_16_20_to_tile_15_20_2;
	wire vertical_tile_16_20_to_tile_15_20_3;

	wire vertical_tile_15_21_to_tile_16_21_0;
	wire vertical_tile_15_21_to_tile_16_21_1;
	wire vertical_tile_15_21_to_tile_16_21_2;
	wire vertical_tile_15_21_to_tile_16_21_3;
	wire vertical_tile_16_21_to_tile_15_21_0;
	wire vertical_tile_16_21_to_tile_15_21_1;
	wire vertical_tile_16_21_to_tile_15_21_2;
	wire vertical_tile_16_21_to_tile_15_21_3;

	wire vertical_tile_15_22_to_tile_16_22_0;
	wire vertical_tile_15_22_to_tile_16_22_1;
	wire vertical_tile_15_22_to_tile_16_22_2;
	wire vertical_tile_15_22_to_tile_16_22_3;
	wire vertical_tile_16_22_to_tile_15_22_0;
	wire vertical_tile_16_22_to_tile_15_22_1;
	wire vertical_tile_16_22_to_tile_15_22_2;
	wire vertical_tile_16_22_to_tile_15_22_3;

	wire vertical_tile_15_23_to_tile_16_23_0;
	wire vertical_tile_15_23_to_tile_16_23_1;
	wire vertical_tile_15_23_to_tile_16_23_2;
	wire vertical_tile_15_23_to_tile_16_23_3;
	wire vertical_tile_16_23_to_tile_15_23_0;
	wire vertical_tile_16_23_to_tile_15_23_1;
	wire vertical_tile_16_23_to_tile_15_23_2;
	wire vertical_tile_16_23_to_tile_15_23_3;

	wire vertical_tile_15_24_to_tile_16_24_0;
	wire vertical_tile_15_24_to_tile_16_24_1;
	wire vertical_tile_15_24_to_tile_16_24_2;
	wire vertical_tile_15_24_to_tile_16_24_3;
	wire vertical_tile_16_24_to_tile_15_24_0;
	wire vertical_tile_16_24_to_tile_15_24_1;
	wire vertical_tile_16_24_to_tile_15_24_2;
	wire vertical_tile_16_24_to_tile_15_24_3;

	wire vertical_tile_15_25_to_tile_16_25_0;
	wire vertical_tile_15_25_to_tile_16_25_1;
	wire vertical_tile_15_25_to_tile_16_25_2;
	wire vertical_tile_15_25_to_tile_16_25_3;
	wire vertical_tile_16_25_to_tile_15_25_0;
	wire vertical_tile_16_25_to_tile_15_25_1;
	wire vertical_tile_16_25_to_tile_15_25_2;
	wire vertical_tile_16_25_to_tile_15_25_3;

	wire vertical_tile_15_26_to_tile_16_26_0;
	wire vertical_tile_15_26_to_tile_16_26_1;
	wire vertical_tile_15_26_to_tile_16_26_2;
	wire vertical_tile_15_26_to_tile_16_26_3;
	wire vertical_tile_16_26_to_tile_15_26_0;
	wire vertical_tile_16_26_to_tile_15_26_1;
	wire vertical_tile_16_26_to_tile_15_26_2;
	wire vertical_tile_16_26_to_tile_15_26_3;

	wire vertical_tile_15_27_to_tile_16_27_0;
	wire vertical_tile_15_27_to_tile_16_27_1;
	wire vertical_tile_15_27_to_tile_16_27_2;
	wire vertical_tile_15_27_to_tile_16_27_3;
	wire vertical_tile_16_27_to_tile_15_27_0;
	wire vertical_tile_16_27_to_tile_15_27_1;
	wire vertical_tile_16_27_to_tile_15_27_2;
	wire vertical_tile_16_27_to_tile_15_27_3;

	wire vertical_tile_15_28_to_tile_16_28_0;
	wire vertical_tile_15_28_to_tile_16_28_1;
	wire vertical_tile_15_28_to_tile_16_28_2;
	wire vertical_tile_15_28_to_tile_16_28_3;
	wire vertical_tile_16_28_to_tile_15_28_0;
	wire vertical_tile_16_28_to_tile_15_28_1;
	wire vertical_tile_16_28_to_tile_15_28_2;
	wire vertical_tile_16_28_to_tile_15_28_3;

	wire vertical_tile_15_29_to_tile_16_29_0;
	wire vertical_tile_15_29_to_tile_16_29_1;
	wire vertical_tile_15_29_to_tile_16_29_2;
	wire vertical_tile_15_29_to_tile_16_29_3;
	wire vertical_tile_16_29_to_tile_15_29_0;
	wire vertical_tile_16_29_to_tile_15_29_1;
	wire vertical_tile_16_29_to_tile_15_29_2;
	wire vertical_tile_16_29_to_tile_15_29_3;

	wire vertical_tile_15_30_to_tile_16_30_0;
	wire vertical_tile_15_30_to_tile_16_30_1;
	wire vertical_tile_15_30_to_tile_16_30_2;
	wire vertical_tile_15_30_to_tile_16_30_3;
	wire vertical_tile_16_30_to_tile_15_30_0;
	wire vertical_tile_16_30_to_tile_15_30_1;
	wire vertical_tile_16_30_to_tile_15_30_2;
	wire vertical_tile_16_30_to_tile_15_30_3;

	wire vertical_tile_15_31_to_tile_16_31_0;
	wire vertical_tile_15_31_to_tile_16_31_1;
	wire vertical_tile_15_31_to_tile_16_31_2;
	wire vertical_tile_15_31_to_tile_16_31_3;
	wire vertical_tile_16_31_to_tile_15_31_0;
	wire vertical_tile_16_31_to_tile_15_31_1;
	wire vertical_tile_16_31_to_tile_15_31_2;
	wire vertical_tile_16_31_to_tile_15_31_3;

	wire vertical_tile_16_0_to_tile_17_0_0;
	wire vertical_tile_16_0_to_tile_17_0_1;
	wire vertical_tile_16_0_to_tile_17_0_2;
	wire vertical_tile_16_0_to_tile_17_0_3;
	wire vertical_tile_17_0_to_tile_16_0_0;
	wire vertical_tile_17_0_to_tile_16_0_1;
	wire vertical_tile_17_0_to_tile_16_0_2;
	wire vertical_tile_17_0_to_tile_16_0_3;

	wire vertical_tile_16_1_to_tile_17_1_0;
	wire vertical_tile_16_1_to_tile_17_1_1;
	wire vertical_tile_16_1_to_tile_17_1_2;
	wire vertical_tile_16_1_to_tile_17_1_3;
	wire vertical_tile_17_1_to_tile_16_1_0;
	wire vertical_tile_17_1_to_tile_16_1_1;
	wire vertical_tile_17_1_to_tile_16_1_2;
	wire vertical_tile_17_1_to_tile_16_1_3;

	wire vertical_tile_16_2_to_tile_17_2_0;
	wire vertical_tile_16_2_to_tile_17_2_1;
	wire vertical_tile_16_2_to_tile_17_2_2;
	wire vertical_tile_16_2_to_tile_17_2_3;
	wire vertical_tile_17_2_to_tile_16_2_0;
	wire vertical_tile_17_2_to_tile_16_2_1;
	wire vertical_tile_17_2_to_tile_16_2_2;
	wire vertical_tile_17_2_to_tile_16_2_3;

	wire vertical_tile_16_3_to_tile_17_3_0;
	wire vertical_tile_16_3_to_tile_17_3_1;
	wire vertical_tile_16_3_to_tile_17_3_2;
	wire vertical_tile_16_3_to_tile_17_3_3;
	wire vertical_tile_17_3_to_tile_16_3_0;
	wire vertical_tile_17_3_to_tile_16_3_1;
	wire vertical_tile_17_3_to_tile_16_3_2;
	wire vertical_tile_17_3_to_tile_16_3_3;

	wire vertical_tile_16_4_to_tile_17_4_0;
	wire vertical_tile_16_4_to_tile_17_4_1;
	wire vertical_tile_16_4_to_tile_17_4_2;
	wire vertical_tile_16_4_to_tile_17_4_3;
	wire vertical_tile_17_4_to_tile_16_4_0;
	wire vertical_tile_17_4_to_tile_16_4_1;
	wire vertical_tile_17_4_to_tile_16_4_2;
	wire vertical_tile_17_4_to_tile_16_4_3;

	wire vertical_tile_16_5_to_tile_17_5_0;
	wire vertical_tile_16_5_to_tile_17_5_1;
	wire vertical_tile_16_5_to_tile_17_5_2;
	wire vertical_tile_16_5_to_tile_17_5_3;
	wire vertical_tile_17_5_to_tile_16_5_0;
	wire vertical_tile_17_5_to_tile_16_5_1;
	wire vertical_tile_17_5_to_tile_16_5_2;
	wire vertical_tile_17_5_to_tile_16_5_3;

	wire vertical_tile_16_6_to_tile_17_6_0;
	wire vertical_tile_16_6_to_tile_17_6_1;
	wire vertical_tile_16_6_to_tile_17_6_2;
	wire vertical_tile_16_6_to_tile_17_6_3;
	wire vertical_tile_17_6_to_tile_16_6_0;
	wire vertical_tile_17_6_to_tile_16_6_1;
	wire vertical_tile_17_6_to_tile_16_6_2;
	wire vertical_tile_17_6_to_tile_16_6_3;

	wire vertical_tile_16_7_to_tile_17_7_0;
	wire vertical_tile_16_7_to_tile_17_7_1;
	wire vertical_tile_16_7_to_tile_17_7_2;
	wire vertical_tile_16_7_to_tile_17_7_3;
	wire vertical_tile_17_7_to_tile_16_7_0;
	wire vertical_tile_17_7_to_tile_16_7_1;
	wire vertical_tile_17_7_to_tile_16_7_2;
	wire vertical_tile_17_7_to_tile_16_7_3;

	wire vertical_tile_16_8_to_tile_17_8_0;
	wire vertical_tile_16_8_to_tile_17_8_1;
	wire vertical_tile_16_8_to_tile_17_8_2;
	wire vertical_tile_16_8_to_tile_17_8_3;
	wire vertical_tile_17_8_to_tile_16_8_0;
	wire vertical_tile_17_8_to_tile_16_8_1;
	wire vertical_tile_17_8_to_tile_16_8_2;
	wire vertical_tile_17_8_to_tile_16_8_3;

	wire vertical_tile_16_9_to_tile_17_9_0;
	wire vertical_tile_16_9_to_tile_17_9_1;
	wire vertical_tile_16_9_to_tile_17_9_2;
	wire vertical_tile_16_9_to_tile_17_9_3;
	wire vertical_tile_17_9_to_tile_16_9_0;
	wire vertical_tile_17_9_to_tile_16_9_1;
	wire vertical_tile_17_9_to_tile_16_9_2;
	wire vertical_tile_17_9_to_tile_16_9_3;

	wire vertical_tile_16_10_to_tile_17_10_0;
	wire vertical_tile_16_10_to_tile_17_10_1;
	wire vertical_tile_16_10_to_tile_17_10_2;
	wire vertical_tile_16_10_to_tile_17_10_3;
	wire vertical_tile_17_10_to_tile_16_10_0;
	wire vertical_tile_17_10_to_tile_16_10_1;
	wire vertical_tile_17_10_to_tile_16_10_2;
	wire vertical_tile_17_10_to_tile_16_10_3;

	wire vertical_tile_16_11_to_tile_17_11_0;
	wire vertical_tile_16_11_to_tile_17_11_1;
	wire vertical_tile_16_11_to_tile_17_11_2;
	wire vertical_tile_16_11_to_tile_17_11_3;
	wire vertical_tile_17_11_to_tile_16_11_0;
	wire vertical_tile_17_11_to_tile_16_11_1;
	wire vertical_tile_17_11_to_tile_16_11_2;
	wire vertical_tile_17_11_to_tile_16_11_3;

	wire vertical_tile_16_12_to_tile_17_12_0;
	wire vertical_tile_16_12_to_tile_17_12_1;
	wire vertical_tile_16_12_to_tile_17_12_2;
	wire vertical_tile_16_12_to_tile_17_12_3;
	wire vertical_tile_17_12_to_tile_16_12_0;
	wire vertical_tile_17_12_to_tile_16_12_1;
	wire vertical_tile_17_12_to_tile_16_12_2;
	wire vertical_tile_17_12_to_tile_16_12_3;

	wire vertical_tile_16_13_to_tile_17_13_0;
	wire vertical_tile_16_13_to_tile_17_13_1;
	wire vertical_tile_16_13_to_tile_17_13_2;
	wire vertical_tile_16_13_to_tile_17_13_3;
	wire vertical_tile_17_13_to_tile_16_13_0;
	wire vertical_tile_17_13_to_tile_16_13_1;
	wire vertical_tile_17_13_to_tile_16_13_2;
	wire vertical_tile_17_13_to_tile_16_13_3;

	wire vertical_tile_16_14_to_tile_17_14_0;
	wire vertical_tile_16_14_to_tile_17_14_1;
	wire vertical_tile_16_14_to_tile_17_14_2;
	wire vertical_tile_16_14_to_tile_17_14_3;
	wire vertical_tile_17_14_to_tile_16_14_0;
	wire vertical_tile_17_14_to_tile_16_14_1;
	wire vertical_tile_17_14_to_tile_16_14_2;
	wire vertical_tile_17_14_to_tile_16_14_3;

	wire vertical_tile_16_15_to_tile_17_15_0;
	wire vertical_tile_16_15_to_tile_17_15_1;
	wire vertical_tile_16_15_to_tile_17_15_2;
	wire vertical_tile_16_15_to_tile_17_15_3;
	wire vertical_tile_17_15_to_tile_16_15_0;
	wire vertical_tile_17_15_to_tile_16_15_1;
	wire vertical_tile_17_15_to_tile_16_15_2;
	wire vertical_tile_17_15_to_tile_16_15_3;

	wire vertical_tile_16_16_to_tile_17_16_0;
	wire vertical_tile_16_16_to_tile_17_16_1;
	wire vertical_tile_16_16_to_tile_17_16_2;
	wire vertical_tile_16_16_to_tile_17_16_3;
	wire vertical_tile_17_16_to_tile_16_16_0;
	wire vertical_tile_17_16_to_tile_16_16_1;
	wire vertical_tile_17_16_to_tile_16_16_2;
	wire vertical_tile_17_16_to_tile_16_16_3;

	wire vertical_tile_16_17_to_tile_17_17_0;
	wire vertical_tile_16_17_to_tile_17_17_1;
	wire vertical_tile_16_17_to_tile_17_17_2;
	wire vertical_tile_16_17_to_tile_17_17_3;
	wire vertical_tile_17_17_to_tile_16_17_0;
	wire vertical_tile_17_17_to_tile_16_17_1;
	wire vertical_tile_17_17_to_tile_16_17_2;
	wire vertical_tile_17_17_to_tile_16_17_3;

	wire vertical_tile_16_18_to_tile_17_18_0;
	wire vertical_tile_16_18_to_tile_17_18_1;
	wire vertical_tile_16_18_to_tile_17_18_2;
	wire vertical_tile_16_18_to_tile_17_18_3;
	wire vertical_tile_17_18_to_tile_16_18_0;
	wire vertical_tile_17_18_to_tile_16_18_1;
	wire vertical_tile_17_18_to_tile_16_18_2;
	wire vertical_tile_17_18_to_tile_16_18_3;

	wire vertical_tile_16_19_to_tile_17_19_0;
	wire vertical_tile_16_19_to_tile_17_19_1;
	wire vertical_tile_16_19_to_tile_17_19_2;
	wire vertical_tile_16_19_to_tile_17_19_3;
	wire vertical_tile_17_19_to_tile_16_19_0;
	wire vertical_tile_17_19_to_tile_16_19_1;
	wire vertical_tile_17_19_to_tile_16_19_2;
	wire vertical_tile_17_19_to_tile_16_19_3;

	wire vertical_tile_16_20_to_tile_17_20_0;
	wire vertical_tile_16_20_to_tile_17_20_1;
	wire vertical_tile_16_20_to_tile_17_20_2;
	wire vertical_tile_16_20_to_tile_17_20_3;
	wire vertical_tile_17_20_to_tile_16_20_0;
	wire vertical_tile_17_20_to_tile_16_20_1;
	wire vertical_tile_17_20_to_tile_16_20_2;
	wire vertical_tile_17_20_to_tile_16_20_3;

	wire vertical_tile_16_21_to_tile_17_21_0;
	wire vertical_tile_16_21_to_tile_17_21_1;
	wire vertical_tile_16_21_to_tile_17_21_2;
	wire vertical_tile_16_21_to_tile_17_21_3;
	wire vertical_tile_17_21_to_tile_16_21_0;
	wire vertical_tile_17_21_to_tile_16_21_1;
	wire vertical_tile_17_21_to_tile_16_21_2;
	wire vertical_tile_17_21_to_tile_16_21_3;

	wire vertical_tile_16_22_to_tile_17_22_0;
	wire vertical_tile_16_22_to_tile_17_22_1;
	wire vertical_tile_16_22_to_tile_17_22_2;
	wire vertical_tile_16_22_to_tile_17_22_3;
	wire vertical_tile_17_22_to_tile_16_22_0;
	wire vertical_tile_17_22_to_tile_16_22_1;
	wire vertical_tile_17_22_to_tile_16_22_2;
	wire vertical_tile_17_22_to_tile_16_22_3;

	wire vertical_tile_16_23_to_tile_17_23_0;
	wire vertical_tile_16_23_to_tile_17_23_1;
	wire vertical_tile_16_23_to_tile_17_23_2;
	wire vertical_tile_16_23_to_tile_17_23_3;
	wire vertical_tile_17_23_to_tile_16_23_0;
	wire vertical_tile_17_23_to_tile_16_23_1;
	wire vertical_tile_17_23_to_tile_16_23_2;
	wire vertical_tile_17_23_to_tile_16_23_3;

	wire vertical_tile_16_24_to_tile_17_24_0;
	wire vertical_tile_16_24_to_tile_17_24_1;
	wire vertical_tile_16_24_to_tile_17_24_2;
	wire vertical_tile_16_24_to_tile_17_24_3;
	wire vertical_tile_17_24_to_tile_16_24_0;
	wire vertical_tile_17_24_to_tile_16_24_1;
	wire vertical_tile_17_24_to_tile_16_24_2;
	wire vertical_tile_17_24_to_tile_16_24_3;

	wire vertical_tile_16_25_to_tile_17_25_0;
	wire vertical_tile_16_25_to_tile_17_25_1;
	wire vertical_tile_16_25_to_tile_17_25_2;
	wire vertical_tile_16_25_to_tile_17_25_3;
	wire vertical_tile_17_25_to_tile_16_25_0;
	wire vertical_tile_17_25_to_tile_16_25_1;
	wire vertical_tile_17_25_to_tile_16_25_2;
	wire vertical_tile_17_25_to_tile_16_25_3;

	wire vertical_tile_16_26_to_tile_17_26_0;
	wire vertical_tile_16_26_to_tile_17_26_1;
	wire vertical_tile_16_26_to_tile_17_26_2;
	wire vertical_tile_16_26_to_tile_17_26_3;
	wire vertical_tile_17_26_to_tile_16_26_0;
	wire vertical_tile_17_26_to_tile_16_26_1;
	wire vertical_tile_17_26_to_tile_16_26_2;
	wire vertical_tile_17_26_to_tile_16_26_3;

	wire vertical_tile_16_27_to_tile_17_27_0;
	wire vertical_tile_16_27_to_tile_17_27_1;
	wire vertical_tile_16_27_to_tile_17_27_2;
	wire vertical_tile_16_27_to_tile_17_27_3;
	wire vertical_tile_17_27_to_tile_16_27_0;
	wire vertical_tile_17_27_to_tile_16_27_1;
	wire vertical_tile_17_27_to_tile_16_27_2;
	wire vertical_tile_17_27_to_tile_16_27_3;

	wire vertical_tile_16_28_to_tile_17_28_0;
	wire vertical_tile_16_28_to_tile_17_28_1;
	wire vertical_tile_16_28_to_tile_17_28_2;
	wire vertical_tile_16_28_to_tile_17_28_3;
	wire vertical_tile_17_28_to_tile_16_28_0;
	wire vertical_tile_17_28_to_tile_16_28_1;
	wire vertical_tile_17_28_to_tile_16_28_2;
	wire vertical_tile_17_28_to_tile_16_28_3;

	wire vertical_tile_16_29_to_tile_17_29_0;
	wire vertical_tile_16_29_to_tile_17_29_1;
	wire vertical_tile_16_29_to_tile_17_29_2;
	wire vertical_tile_16_29_to_tile_17_29_3;
	wire vertical_tile_17_29_to_tile_16_29_0;
	wire vertical_tile_17_29_to_tile_16_29_1;
	wire vertical_tile_17_29_to_tile_16_29_2;
	wire vertical_tile_17_29_to_tile_16_29_3;

	wire vertical_tile_16_30_to_tile_17_30_0;
	wire vertical_tile_16_30_to_tile_17_30_1;
	wire vertical_tile_16_30_to_tile_17_30_2;
	wire vertical_tile_16_30_to_tile_17_30_3;
	wire vertical_tile_17_30_to_tile_16_30_0;
	wire vertical_tile_17_30_to_tile_16_30_1;
	wire vertical_tile_17_30_to_tile_16_30_2;
	wire vertical_tile_17_30_to_tile_16_30_3;

	wire vertical_tile_16_31_to_tile_17_31_0;
	wire vertical_tile_16_31_to_tile_17_31_1;
	wire vertical_tile_16_31_to_tile_17_31_2;
	wire vertical_tile_16_31_to_tile_17_31_3;
	wire vertical_tile_17_31_to_tile_16_31_0;
	wire vertical_tile_17_31_to_tile_16_31_1;
	wire vertical_tile_17_31_to_tile_16_31_2;
	wire vertical_tile_17_31_to_tile_16_31_3;

	wire vertical_tile_17_0_to_tile_18_0_0;
	wire vertical_tile_17_0_to_tile_18_0_1;
	wire vertical_tile_17_0_to_tile_18_0_2;
	wire vertical_tile_17_0_to_tile_18_0_3;
	wire vertical_tile_18_0_to_tile_17_0_0;
	wire vertical_tile_18_0_to_tile_17_0_1;
	wire vertical_tile_18_0_to_tile_17_0_2;
	wire vertical_tile_18_0_to_tile_17_0_3;

	wire vertical_tile_17_1_to_tile_18_1_0;
	wire vertical_tile_17_1_to_tile_18_1_1;
	wire vertical_tile_17_1_to_tile_18_1_2;
	wire vertical_tile_17_1_to_tile_18_1_3;
	wire vertical_tile_18_1_to_tile_17_1_0;
	wire vertical_tile_18_1_to_tile_17_1_1;
	wire vertical_tile_18_1_to_tile_17_1_2;
	wire vertical_tile_18_1_to_tile_17_1_3;

	wire vertical_tile_17_2_to_tile_18_2_0;
	wire vertical_tile_17_2_to_tile_18_2_1;
	wire vertical_tile_17_2_to_tile_18_2_2;
	wire vertical_tile_17_2_to_tile_18_2_3;
	wire vertical_tile_18_2_to_tile_17_2_0;
	wire vertical_tile_18_2_to_tile_17_2_1;
	wire vertical_tile_18_2_to_tile_17_2_2;
	wire vertical_tile_18_2_to_tile_17_2_3;

	wire vertical_tile_17_3_to_tile_18_3_0;
	wire vertical_tile_17_3_to_tile_18_3_1;
	wire vertical_tile_17_3_to_tile_18_3_2;
	wire vertical_tile_17_3_to_tile_18_3_3;
	wire vertical_tile_18_3_to_tile_17_3_0;
	wire vertical_tile_18_3_to_tile_17_3_1;
	wire vertical_tile_18_3_to_tile_17_3_2;
	wire vertical_tile_18_3_to_tile_17_3_3;

	wire vertical_tile_17_4_to_tile_18_4_0;
	wire vertical_tile_17_4_to_tile_18_4_1;
	wire vertical_tile_17_4_to_tile_18_4_2;
	wire vertical_tile_17_4_to_tile_18_4_3;
	wire vertical_tile_18_4_to_tile_17_4_0;
	wire vertical_tile_18_4_to_tile_17_4_1;
	wire vertical_tile_18_4_to_tile_17_4_2;
	wire vertical_tile_18_4_to_tile_17_4_3;

	wire vertical_tile_17_5_to_tile_18_5_0;
	wire vertical_tile_17_5_to_tile_18_5_1;
	wire vertical_tile_17_5_to_tile_18_5_2;
	wire vertical_tile_17_5_to_tile_18_5_3;
	wire vertical_tile_18_5_to_tile_17_5_0;
	wire vertical_tile_18_5_to_tile_17_5_1;
	wire vertical_tile_18_5_to_tile_17_5_2;
	wire vertical_tile_18_5_to_tile_17_5_3;

	wire vertical_tile_17_6_to_tile_18_6_0;
	wire vertical_tile_17_6_to_tile_18_6_1;
	wire vertical_tile_17_6_to_tile_18_6_2;
	wire vertical_tile_17_6_to_tile_18_6_3;
	wire vertical_tile_18_6_to_tile_17_6_0;
	wire vertical_tile_18_6_to_tile_17_6_1;
	wire vertical_tile_18_6_to_tile_17_6_2;
	wire vertical_tile_18_6_to_tile_17_6_3;

	wire vertical_tile_17_7_to_tile_18_7_0;
	wire vertical_tile_17_7_to_tile_18_7_1;
	wire vertical_tile_17_7_to_tile_18_7_2;
	wire vertical_tile_17_7_to_tile_18_7_3;
	wire vertical_tile_18_7_to_tile_17_7_0;
	wire vertical_tile_18_7_to_tile_17_7_1;
	wire vertical_tile_18_7_to_tile_17_7_2;
	wire vertical_tile_18_7_to_tile_17_7_3;

	wire vertical_tile_17_8_to_tile_18_8_0;
	wire vertical_tile_17_8_to_tile_18_8_1;
	wire vertical_tile_17_8_to_tile_18_8_2;
	wire vertical_tile_17_8_to_tile_18_8_3;
	wire vertical_tile_18_8_to_tile_17_8_0;
	wire vertical_tile_18_8_to_tile_17_8_1;
	wire vertical_tile_18_8_to_tile_17_8_2;
	wire vertical_tile_18_8_to_tile_17_8_3;

	wire vertical_tile_17_9_to_tile_18_9_0;
	wire vertical_tile_17_9_to_tile_18_9_1;
	wire vertical_tile_17_9_to_tile_18_9_2;
	wire vertical_tile_17_9_to_tile_18_9_3;
	wire vertical_tile_18_9_to_tile_17_9_0;
	wire vertical_tile_18_9_to_tile_17_9_1;
	wire vertical_tile_18_9_to_tile_17_9_2;
	wire vertical_tile_18_9_to_tile_17_9_3;

	wire vertical_tile_17_10_to_tile_18_10_0;
	wire vertical_tile_17_10_to_tile_18_10_1;
	wire vertical_tile_17_10_to_tile_18_10_2;
	wire vertical_tile_17_10_to_tile_18_10_3;
	wire vertical_tile_18_10_to_tile_17_10_0;
	wire vertical_tile_18_10_to_tile_17_10_1;
	wire vertical_tile_18_10_to_tile_17_10_2;
	wire vertical_tile_18_10_to_tile_17_10_3;

	wire vertical_tile_17_11_to_tile_18_11_0;
	wire vertical_tile_17_11_to_tile_18_11_1;
	wire vertical_tile_17_11_to_tile_18_11_2;
	wire vertical_tile_17_11_to_tile_18_11_3;
	wire vertical_tile_18_11_to_tile_17_11_0;
	wire vertical_tile_18_11_to_tile_17_11_1;
	wire vertical_tile_18_11_to_tile_17_11_2;
	wire vertical_tile_18_11_to_tile_17_11_3;

	wire vertical_tile_17_12_to_tile_18_12_0;
	wire vertical_tile_17_12_to_tile_18_12_1;
	wire vertical_tile_17_12_to_tile_18_12_2;
	wire vertical_tile_17_12_to_tile_18_12_3;
	wire vertical_tile_18_12_to_tile_17_12_0;
	wire vertical_tile_18_12_to_tile_17_12_1;
	wire vertical_tile_18_12_to_tile_17_12_2;
	wire vertical_tile_18_12_to_tile_17_12_3;

	wire vertical_tile_17_13_to_tile_18_13_0;
	wire vertical_tile_17_13_to_tile_18_13_1;
	wire vertical_tile_17_13_to_tile_18_13_2;
	wire vertical_tile_17_13_to_tile_18_13_3;
	wire vertical_tile_18_13_to_tile_17_13_0;
	wire vertical_tile_18_13_to_tile_17_13_1;
	wire vertical_tile_18_13_to_tile_17_13_2;
	wire vertical_tile_18_13_to_tile_17_13_3;

	wire vertical_tile_17_14_to_tile_18_14_0;
	wire vertical_tile_17_14_to_tile_18_14_1;
	wire vertical_tile_17_14_to_tile_18_14_2;
	wire vertical_tile_17_14_to_tile_18_14_3;
	wire vertical_tile_18_14_to_tile_17_14_0;
	wire vertical_tile_18_14_to_tile_17_14_1;
	wire vertical_tile_18_14_to_tile_17_14_2;
	wire vertical_tile_18_14_to_tile_17_14_3;

	wire vertical_tile_17_15_to_tile_18_15_0;
	wire vertical_tile_17_15_to_tile_18_15_1;
	wire vertical_tile_17_15_to_tile_18_15_2;
	wire vertical_tile_17_15_to_tile_18_15_3;
	wire vertical_tile_18_15_to_tile_17_15_0;
	wire vertical_tile_18_15_to_tile_17_15_1;
	wire vertical_tile_18_15_to_tile_17_15_2;
	wire vertical_tile_18_15_to_tile_17_15_3;

	wire vertical_tile_17_16_to_tile_18_16_0;
	wire vertical_tile_17_16_to_tile_18_16_1;
	wire vertical_tile_17_16_to_tile_18_16_2;
	wire vertical_tile_17_16_to_tile_18_16_3;
	wire vertical_tile_18_16_to_tile_17_16_0;
	wire vertical_tile_18_16_to_tile_17_16_1;
	wire vertical_tile_18_16_to_tile_17_16_2;
	wire vertical_tile_18_16_to_tile_17_16_3;

	wire vertical_tile_17_17_to_tile_18_17_0;
	wire vertical_tile_17_17_to_tile_18_17_1;
	wire vertical_tile_17_17_to_tile_18_17_2;
	wire vertical_tile_17_17_to_tile_18_17_3;
	wire vertical_tile_18_17_to_tile_17_17_0;
	wire vertical_tile_18_17_to_tile_17_17_1;
	wire vertical_tile_18_17_to_tile_17_17_2;
	wire vertical_tile_18_17_to_tile_17_17_3;

	wire vertical_tile_17_18_to_tile_18_18_0;
	wire vertical_tile_17_18_to_tile_18_18_1;
	wire vertical_tile_17_18_to_tile_18_18_2;
	wire vertical_tile_17_18_to_tile_18_18_3;
	wire vertical_tile_18_18_to_tile_17_18_0;
	wire vertical_tile_18_18_to_tile_17_18_1;
	wire vertical_tile_18_18_to_tile_17_18_2;
	wire vertical_tile_18_18_to_tile_17_18_3;

	wire vertical_tile_17_19_to_tile_18_19_0;
	wire vertical_tile_17_19_to_tile_18_19_1;
	wire vertical_tile_17_19_to_tile_18_19_2;
	wire vertical_tile_17_19_to_tile_18_19_3;
	wire vertical_tile_18_19_to_tile_17_19_0;
	wire vertical_tile_18_19_to_tile_17_19_1;
	wire vertical_tile_18_19_to_tile_17_19_2;
	wire vertical_tile_18_19_to_tile_17_19_3;

	wire vertical_tile_17_20_to_tile_18_20_0;
	wire vertical_tile_17_20_to_tile_18_20_1;
	wire vertical_tile_17_20_to_tile_18_20_2;
	wire vertical_tile_17_20_to_tile_18_20_3;
	wire vertical_tile_18_20_to_tile_17_20_0;
	wire vertical_tile_18_20_to_tile_17_20_1;
	wire vertical_tile_18_20_to_tile_17_20_2;
	wire vertical_tile_18_20_to_tile_17_20_3;

	wire vertical_tile_17_21_to_tile_18_21_0;
	wire vertical_tile_17_21_to_tile_18_21_1;
	wire vertical_tile_17_21_to_tile_18_21_2;
	wire vertical_tile_17_21_to_tile_18_21_3;
	wire vertical_tile_18_21_to_tile_17_21_0;
	wire vertical_tile_18_21_to_tile_17_21_1;
	wire vertical_tile_18_21_to_tile_17_21_2;
	wire vertical_tile_18_21_to_tile_17_21_3;

	wire vertical_tile_17_22_to_tile_18_22_0;
	wire vertical_tile_17_22_to_tile_18_22_1;
	wire vertical_tile_17_22_to_tile_18_22_2;
	wire vertical_tile_17_22_to_tile_18_22_3;
	wire vertical_tile_18_22_to_tile_17_22_0;
	wire vertical_tile_18_22_to_tile_17_22_1;
	wire vertical_tile_18_22_to_tile_17_22_2;
	wire vertical_tile_18_22_to_tile_17_22_3;

	wire vertical_tile_17_23_to_tile_18_23_0;
	wire vertical_tile_17_23_to_tile_18_23_1;
	wire vertical_tile_17_23_to_tile_18_23_2;
	wire vertical_tile_17_23_to_tile_18_23_3;
	wire vertical_tile_18_23_to_tile_17_23_0;
	wire vertical_tile_18_23_to_tile_17_23_1;
	wire vertical_tile_18_23_to_tile_17_23_2;
	wire vertical_tile_18_23_to_tile_17_23_3;

	wire vertical_tile_17_24_to_tile_18_24_0;
	wire vertical_tile_17_24_to_tile_18_24_1;
	wire vertical_tile_17_24_to_tile_18_24_2;
	wire vertical_tile_17_24_to_tile_18_24_3;
	wire vertical_tile_18_24_to_tile_17_24_0;
	wire vertical_tile_18_24_to_tile_17_24_1;
	wire vertical_tile_18_24_to_tile_17_24_2;
	wire vertical_tile_18_24_to_tile_17_24_3;

	wire vertical_tile_17_25_to_tile_18_25_0;
	wire vertical_tile_17_25_to_tile_18_25_1;
	wire vertical_tile_17_25_to_tile_18_25_2;
	wire vertical_tile_17_25_to_tile_18_25_3;
	wire vertical_tile_18_25_to_tile_17_25_0;
	wire vertical_tile_18_25_to_tile_17_25_1;
	wire vertical_tile_18_25_to_tile_17_25_2;
	wire vertical_tile_18_25_to_tile_17_25_3;

	wire vertical_tile_17_26_to_tile_18_26_0;
	wire vertical_tile_17_26_to_tile_18_26_1;
	wire vertical_tile_17_26_to_tile_18_26_2;
	wire vertical_tile_17_26_to_tile_18_26_3;
	wire vertical_tile_18_26_to_tile_17_26_0;
	wire vertical_tile_18_26_to_tile_17_26_1;
	wire vertical_tile_18_26_to_tile_17_26_2;
	wire vertical_tile_18_26_to_tile_17_26_3;

	wire vertical_tile_17_27_to_tile_18_27_0;
	wire vertical_tile_17_27_to_tile_18_27_1;
	wire vertical_tile_17_27_to_tile_18_27_2;
	wire vertical_tile_17_27_to_tile_18_27_3;
	wire vertical_tile_18_27_to_tile_17_27_0;
	wire vertical_tile_18_27_to_tile_17_27_1;
	wire vertical_tile_18_27_to_tile_17_27_2;
	wire vertical_tile_18_27_to_tile_17_27_3;

	wire vertical_tile_17_28_to_tile_18_28_0;
	wire vertical_tile_17_28_to_tile_18_28_1;
	wire vertical_tile_17_28_to_tile_18_28_2;
	wire vertical_tile_17_28_to_tile_18_28_3;
	wire vertical_tile_18_28_to_tile_17_28_0;
	wire vertical_tile_18_28_to_tile_17_28_1;
	wire vertical_tile_18_28_to_tile_17_28_2;
	wire vertical_tile_18_28_to_tile_17_28_3;

	wire vertical_tile_17_29_to_tile_18_29_0;
	wire vertical_tile_17_29_to_tile_18_29_1;
	wire vertical_tile_17_29_to_tile_18_29_2;
	wire vertical_tile_17_29_to_tile_18_29_3;
	wire vertical_tile_18_29_to_tile_17_29_0;
	wire vertical_tile_18_29_to_tile_17_29_1;
	wire vertical_tile_18_29_to_tile_17_29_2;
	wire vertical_tile_18_29_to_tile_17_29_3;

	wire vertical_tile_17_30_to_tile_18_30_0;
	wire vertical_tile_17_30_to_tile_18_30_1;
	wire vertical_tile_17_30_to_tile_18_30_2;
	wire vertical_tile_17_30_to_tile_18_30_3;
	wire vertical_tile_18_30_to_tile_17_30_0;
	wire vertical_tile_18_30_to_tile_17_30_1;
	wire vertical_tile_18_30_to_tile_17_30_2;
	wire vertical_tile_18_30_to_tile_17_30_3;

	wire vertical_tile_17_31_to_tile_18_31_0;
	wire vertical_tile_17_31_to_tile_18_31_1;
	wire vertical_tile_17_31_to_tile_18_31_2;
	wire vertical_tile_17_31_to_tile_18_31_3;
	wire vertical_tile_18_31_to_tile_17_31_0;
	wire vertical_tile_18_31_to_tile_17_31_1;
	wire vertical_tile_18_31_to_tile_17_31_2;
	wire vertical_tile_18_31_to_tile_17_31_3;

	wire vertical_tile_18_0_to_tile_19_0_0;
	wire vertical_tile_18_0_to_tile_19_0_1;
	wire vertical_tile_18_0_to_tile_19_0_2;
	wire vertical_tile_18_0_to_tile_19_0_3;
	wire vertical_tile_19_0_to_tile_18_0_0;
	wire vertical_tile_19_0_to_tile_18_0_1;
	wire vertical_tile_19_0_to_tile_18_0_2;
	wire vertical_tile_19_0_to_tile_18_0_3;

	wire vertical_tile_18_1_to_tile_19_1_0;
	wire vertical_tile_18_1_to_tile_19_1_1;
	wire vertical_tile_18_1_to_tile_19_1_2;
	wire vertical_tile_18_1_to_tile_19_1_3;
	wire vertical_tile_19_1_to_tile_18_1_0;
	wire vertical_tile_19_1_to_tile_18_1_1;
	wire vertical_tile_19_1_to_tile_18_1_2;
	wire vertical_tile_19_1_to_tile_18_1_3;

	wire vertical_tile_18_2_to_tile_19_2_0;
	wire vertical_tile_18_2_to_tile_19_2_1;
	wire vertical_tile_18_2_to_tile_19_2_2;
	wire vertical_tile_18_2_to_tile_19_2_3;
	wire vertical_tile_19_2_to_tile_18_2_0;
	wire vertical_tile_19_2_to_tile_18_2_1;
	wire vertical_tile_19_2_to_tile_18_2_2;
	wire vertical_tile_19_2_to_tile_18_2_3;

	wire vertical_tile_18_3_to_tile_19_3_0;
	wire vertical_tile_18_3_to_tile_19_3_1;
	wire vertical_tile_18_3_to_tile_19_3_2;
	wire vertical_tile_18_3_to_tile_19_3_3;
	wire vertical_tile_19_3_to_tile_18_3_0;
	wire vertical_tile_19_3_to_tile_18_3_1;
	wire vertical_tile_19_3_to_tile_18_3_2;
	wire vertical_tile_19_3_to_tile_18_3_3;

	wire vertical_tile_18_4_to_tile_19_4_0;
	wire vertical_tile_18_4_to_tile_19_4_1;
	wire vertical_tile_18_4_to_tile_19_4_2;
	wire vertical_tile_18_4_to_tile_19_4_3;
	wire vertical_tile_19_4_to_tile_18_4_0;
	wire vertical_tile_19_4_to_tile_18_4_1;
	wire vertical_tile_19_4_to_tile_18_4_2;
	wire vertical_tile_19_4_to_tile_18_4_3;

	wire vertical_tile_18_5_to_tile_19_5_0;
	wire vertical_tile_18_5_to_tile_19_5_1;
	wire vertical_tile_18_5_to_tile_19_5_2;
	wire vertical_tile_18_5_to_tile_19_5_3;
	wire vertical_tile_19_5_to_tile_18_5_0;
	wire vertical_tile_19_5_to_tile_18_5_1;
	wire vertical_tile_19_5_to_tile_18_5_2;
	wire vertical_tile_19_5_to_tile_18_5_3;

	wire vertical_tile_18_6_to_tile_19_6_0;
	wire vertical_tile_18_6_to_tile_19_6_1;
	wire vertical_tile_18_6_to_tile_19_6_2;
	wire vertical_tile_18_6_to_tile_19_6_3;
	wire vertical_tile_19_6_to_tile_18_6_0;
	wire vertical_tile_19_6_to_tile_18_6_1;
	wire vertical_tile_19_6_to_tile_18_6_2;
	wire vertical_tile_19_6_to_tile_18_6_3;

	wire vertical_tile_18_7_to_tile_19_7_0;
	wire vertical_tile_18_7_to_tile_19_7_1;
	wire vertical_tile_18_7_to_tile_19_7_2;
	wire vertical_tile_18_7_to_tile_19_7_3;
	wire vertical_tile_19_7_to_tile_18_7_0;
	wire vertical_tile_19_7_to_tile_18_7_1;
	wire vertical_tile_19_7_to_tile_18_7_2;
	wire vertical_tile_19_7_to_tile_18_7_3;

	wire vertical_tile_18_8_to_tile_19_8_0;
	wire vertical_tile_18_8_to_tile_19_8_1;
	wire vertical_tile_18_8_to_tile_19_8_2;
	wire vertical_tile_18_8_to_tile_19_8_3;
	wire vertical_tile_19_8_to_tile_18_8_0;
	wire vertical_tile_19_8_to_tile_18_8_1;
	wire vertical_tile_19_8_to_tile_18_8_2;
	wire vertical_tile_19_8_to_tile_18_8_3;

	wire vertical_tile_18_9_to_tile_19_9_0;
	wire vertical_tile_18_9_to_tile_19_9_1;
	wire vertical_tile_18_9_to_tile_19_9_2;
	wire vertical_tile_18_9_to_tile_19_9_3;
	wire vertical_tile_19_9_to_tile_18_9_0;
	wire vertical_tile_19_9_to_tile_18_9_1;
	wire vertical_tile_19_9_to_tile_18_9_2;
	wire vertical_tile_19_9_to_tile_18_9_3;

	wire vertical_tile_18_10_to_tile_19_10_0;
	wire vertical_tile_18_10_to_tile_19_10_1;
	wire vertical_tile_18_10_to_tile_19_10_2;
	wire vertical_tile_18_10_to_tile_19_10_3;
	wire vertical_tile_19_10_to_tile_18_10_0;
	wire vertical_tile_19_10_to_tile_18_10_1;
	wire vertical_tile_19_10_to_tile_18_10_2;
	wire vertical_tile_19_10_to_tile_18_10_3;

	wire vertical_tile_18_11_to_tile_19_11_0;
	wire vertical_tile_18_11_to_tile_19_11_1;
	wire vertical_tile_18_11_to_tile_19_11_2;
	wire vertical_tile_18_11_to_tile_19_11_3;
	wire vertical_tile_19_11_to_tile_18_11_0;
	wire vertical_tile_19_11_to_tile_18_11_1;
	wire vertical_tile_19_11_to_tile_18_11_2;
	wire vertical_tile_19_11_to_tile_18_11_3;

	wire vertical_tile_18_12_to_tile_19_12_0;
	wire vertical_tile_18_12_to_tile_19_12_1;
	wire vertical_tile_18_12_to_tile_19_12_2;
	wire vertical_tile_18_12_to_tile_19_12_3;
	wire vertical_tile_19_12_to_tile_18_12_0;
	wire vertical_tile_19_12_to_tile_18_12_1;
	wire vertical_tile_19_12_to_tile_18_12_2;
	wire vertical_tile_19_12_to_tile_18_12_3;

	wire vertical_tile_18_13_to_tile_19_13_0;
	wire vertical_tile_18_13_to_tile_19_13_1;
	wire vertical_tile_18_13_to_tile_19_13_2;
	wire vertical_tile_18_13_to_tile_19_13_3;
	wire vertical_tile_19_13_to_tile_18_13_0;
	wire vertical_tile_19_13_to_tile_18_13_1;
	wire vertical_tile_19_13_to_tile_18_13_2;
	wire vertical_tile_19_13_to_tile_18_13_3;

	wire vertical_tile_18_14_to_tile_19_14_0;
	wire vertical_tile_18_14_to_tile_19_14_1;
	wire vertical_tile_18_14_to_tile_19_14_2;
	wire vertical_tile_18_14_to_tile_19_14_3;
	wire vertical_tile_19_14_to_tile_18_14_0;
	wire vertical_tile_19_14_to_tile_18_14_1;
	wire vertical_tile_19_14_to_tile_18_14_2;
	wire vertical_tile_19_14_to_tile_18_14_3;

	wire vertical_tile_18_15_to_tile_19_15_0;
	wire vertical_tile_18_15_to_tile_19_15_1;
	wire vertical_tile_18_15_to_tile_19_15_2;
	wire vertical_tile_18_15_to_tile_19_15_3;
	wire vertical_tile_19_15_to_tile_18_15_0;
	wire vertical_tile_19_15_to_tile_18_15_1;
	wire vertical_tile_19_15_to_tile_18_15_2;
	wire vertical_tile_19_15_to_tile_18_15_3;

	wire vertical_tile_18_16_to_tile_19_16_0;
	wire vertical_tile_18_16_to_tile_19_16_1;
	wire vertical_tile_18_16_to_tile_19_16_2;
	wire vertical_tile_18_16_to_tile_19_16_3;
	wire vertical_tile_19_16_to_tile_18_16_0;
	wire vertical_tile_19_16_to_tile_18_16_1;
	wire vertical_tile_19_16_to_tile_18_16_2;
	wire vertical_tile_19_16_to_tile_18_16_3;

	wire vertical_tile_18_17_to_tile_19_17_0;
	wire vertical_tile_18_17_to_tile_19_17_1;
	wire vertical_tile_18_17_to_tile_19_17_2;
	wire vertical_tile_18_17_to_tile_19_17_3;
	wire vertical_tile_19_17_to_tile_18_17_0;
	wire vertical_tile_19_17_to_tile_18_17_1;
	wire vertical_tile_19_17_to_tile_18_17_2;
	wire vertical_tile_19_17_to_tile_18_17_3;

	wire vertical_tile_18_18_to_tile_19_18_0;
	wire vertical_tile_18_18_to_tile_19_18_1;
	wire vertical_tile_18_18_to_tile_19_18_2;
	wire vertical_tile_18_18_to_tile_19_18_3;
	wire vertical_tile_19_18_to_tile_18_18_0;
	wire vertical_tile_19_18_to_tile_18_18_1;
	wire vertical_tile_19_18_to_tile_18_18_2;
	wire vertical_tile_19_18_to_tile_18_18_3;

	wire vertical_tile_18_19_to_tile_19_19_0;
	wire vertical_tile_18_19_to_tile_19_19_1;
	wire vertical_tile_18_19_to_tile_19_19_2;
	wire vertical_tile_18_19_to_tile_19_19_3;
	wire vertical_tile_19_19_to_tile_18_19_0;
	wire vertical_tile_19_19_to_tile_18_19_1;
	wire vertical_tile_19_19_to_tile_18_19_2;
	wire vertical_tile_19_19_to_tile_18_19_3;

	wire vertical_tile_18_20_to_tile_19_20_0;
	wire vertical_tile_18_20_to_tile_19_20_1;
	wire vertical_tile_18_20_to_tile_19_20_2;
	wire vertical_tile_18_20_to_tile_19_20_3;
	wire vertical_tile_19_20_to_tile_18_20_0;
	wire vertical_tile_19_20_to_tile_18_20_1;
	wire vertical_tile_19_20_to_tile_18_20_2;
	wire vertical_tile_19_20_to_tile_18_20_3;

	wire vertical_tile_18_21_to_tile_19_21_0;
	wire vertical_tile_18_21_to_tile_19_21_1;
	wire vertical_tile_18_21_to_tile_19_21_2;
	wire vertical_tile_18_21_to_tile_19_21_3;
	wire vertical_tile_19_21_to_tile_18_21_0;
	wire vertical_tile_19_21_to_tile_18_21_1;
	wire vertical_tile_19_21_to_tile_18_21_2;
	wire vertical_tile_19_21_to_tile_18_21_3;

	wire vertical_tile_18_22_to_tile_19_22_0;
	wire vertical_tile_18_22_to_tile_19_22_1;
	wire vertical_tile_18_22_to_tile_19_22_2;
	wire vertical_tile_18_22_to_tile_19_22_3;
	wire vertical_tile_19_22_to_tile_18_22_0;
	wire vertical_tile_19_22_to_tile_18_22_1;
	wire vertical_tile_19_22_to_tile_18_22_2;
	wire vertical_tile_19_22_to_tile_18_22_3;

	wire vertical_tile_18_23_to_tile_19_23_0;
	wire vertical_tile_18_23_to_tile_19_23_1;
	wire vertical_tile_18_23_to_tile_19_23_2;
	wire vertical_tile_18_23_to_tile_19_23_3;
	wire vertical_tile_19_23_to_tile_18_23_0;
	wire vertical_tile_19_23_to_tile_18_23_1;
	wire vertical_tile_19_23_to_tile_18_23_2;
	wire vertical_tile_19_23_to_tile_18_23_3;

	wire vertical_tile_18_24_to_tile_19_24_0;
	wire vertical_tile_18_24_to_tile_19_24_1;
	wire vertical_tile_18_24_to_tile_19_24_2;
	wire vertical_tile_18_24_to_tile_19_24_3;
	wire vertical_tile_19_24_to_tile_18_24_0;
	wire vertical_tile_19_24_to_tile_18_24_1;
	wire vertical_tile_19_24_to_tile_18_24_2;
	wire vertical_tile_19_24_to_tile_18_24_3;

	wire vertical_tile_18_25_to_tile_19_25_0;
	wire vertical_tile_18_25_to_tile_19_25_1;
	wire vertical_tile_18_25_to_tile_19_25_2;
	wire vertical_tile_18_25_to_tile_19_25_3;
	wire vertical_tile_19_25_to_tile_18_25_0;
	wire vertical_tile_19_25_to_tile_18_25_1;
	wire vertical_tile_19_25_to_tile_18_25_2;
	wire vertical_tile_19_25_to_tile_18_25_3;

	wire vertical_tile_18_26_to_tile_19_26_0;
	wire vertical_tile_18_26_to_tile_19_26_1;
	wire vertical_tile_18_26_to_tile_19_26_2;
	wire vertical_tile_18_26_to_tile_19_26_3;
	wire vertical_tile_19_26_to_tile_18_26_0;
	wire vertical_tile_19_26_to_tile_18_26_1;
	wire vertical_tile_19_26_to_tile_18_26_2;
	wire vertical_tile_19_26_to_tile_18_26_3;

	wire vertical_tile_18_27_to_tile_19_27_0;
	wire vertical_tile_18_27_to_tile_19_27_1;
	wire vertical_tile_18_27_to_tile_19_27_2;
	wire vertical_tile_18_27_to_tile_19_27_3;
	wire vertical_tile_19_27_to_tile_18_27_0;
	wire vertical_tile_19_27_to_tile_18_27_1;
	wire vertical_tile_19_27_to_tile_18_27_2;
	wire vertical_tile_19_27_to_tile_18_27_3;

	wire vertical_tile_18_28_to_tile_19_28_0;
	wire vertical_tile_18_28_to_tile_19_28_1;
	wire vertical_tile_18_28_to_tile_19_28_2;
	wire vertical_tile_18_28_to_tile_19_28_3;
	wire vertical_tile_19_28_to_tile_18_28_0;
	wire vertical_tile_19_28_to_tile_18_28_1;
	wire vertical_tile_19_28_to_tile_18_28_2;
	wire vertical_tile_19_28_to_tile_18_28_3;

	wire vertical_tile_18_29_to_tile_19_29_0;
	wire vertical_tile_18_29_to_tile_19_29_1;
	wire vertical_tile_18_29_to_tile_19_29_2;
	wire vertical_tile_18_29_to_tile_19_29_3;
	wire vertical_tile_19_29_to_tile_18_29_0;
	wire vertical_tile_19_29_to_tile_18_29_1;
	wire vertical_tile_19_29_to_tile_18_29_2;
	wire vertical_tile_19_29_to_tile_18_29_3;

	wire vertical_tile_18_30_to_tile_19_30_0;
	wire vertical_tile_18_30_to_tile_19_30_1;
	wire vertical_tile_18_30_to_tile_19_30_2;
	wire vertical_tile_18_30_to_tile_19_30_3;
	wire vertical_tile_19_30_to_tile_18_30_0;
	wire vertical_tile_19_30_to_tile_18_30_1;
	wire vertical_tile_19_30_to_tile_18_30_2;
	wire vertical_tile_19_30_to_tile_18_30_3;

	wire vertical_tile_18_31_to_tile_19_31_0;
	wire vertical_tile_18_31_to_tile_19_31_1;
	wire vertical_tile_18_31_to_tile_19_31_2;
	wire vertical_tile_18_31_to_tile_19_31_3;
	wire vertical_tile_19_31_to_tile_18_31_0;
	wire vertical_tile_19_31_to_tile_18_31_1;
	wire vertical_tile_19_31_to_tile_18_31_2;
	wire vertical_tile_19_31_to_tile_18_31_3;

	wire vertical_tile_19_0_to_tile_20_0_0;
	wire vertical_tile_19_0_to_tile_20_0_1;
	wire vertical_tile_19_0_to_tile_20_0_2;
	wire vertical_tile_19_0_to_tile_20_0_3;
	wire vertical_tile_20_0_to_tile_19_0_0;
	wire vertical_tile_20_0_to_tile_19_0_1;
	wire vertical_tile_20_0_to_tile_19_0_2;
	wire vertical_tile_20_0_to_tile_19_0_3;

	wire vertical_tile_19_1_to_tile_20_1_0;
	wire vertical_tile_19_1_to_tile_20_1_1;
	wire vertical_tile_19_1_to_tile_20_1_2;
	wire vertical_tile_19_1_to_tile_20_1_3;
	wire vertical_tile_20_1_to_tile_19_1_0;
	wire vertical_tile_20_1_to_tile_19_1_1;
	wire vertical_tile_20_1_to_tile_19_1_2;
	wire vertical_tile_20_1_to_tile_19_1_3;

	wire vertical_tile_19_2_to_tile_20_2_0;
	wire vertical_tile_19_2_to_tile_20_2_1;
	wire vertical_tile_19_2_to_tile_20_2_2;
	wire vertical_tile_19_2_to_tile_20_2_3;
	wire vertical_tile_20_2_to_tile_19_2_0;
	wire vertical_tile_20_2_to_tile_19_2_1;
	wire vertical_tile_20_2_to_tile_19_2_2;
	wire vertical_tile_20_2_to_tile_19_2_3;

	wire vertical_tile_19_3_to_tile_20_3_0;
	wire vertical_tile_19_3_to_tile_20_3_1;
	wire vertical_tile_19_3_to_tile_20_3_2;
	wire vertical_tile_19_3_to_tile_20_3_3;
	wire vertical_tile_20_3_to_tile_19_3_0;
	wire vertical_tile_20_3_to_tile_19_3_1;
	wire vertical_tile_20_3_to_tile_19_3_2;
	wire vertical_tile_20_3_to_tile_19_3_3;

	wire vertical_tile_19_4_to_tile_20_4_0;
	wire vertical_tile_19_4_to_tile_20_4_1;
	wire vertical_tile_19_4_to_tile_20_4_2;
	wire vertical_tile_19_4_to_tile_20_4_3;
	wire vertical_tile_20_4_to_tile_19_4_0;
	wire vertical_tile_20_4_to_tile_19_4_1;
	wire vertical_tile_20_4_to_tile_19_4_2;
	wire vertical_tile_20_4_to_tile_19_4_3;

	wire vertical_tile_19_5_to_tile_20_5_0;
	wire vertical_tile_19_5_to_tile_20_5_1;
	wire vertical_tile_19_5_to_tile_20_5_2;
	wire vertical_tile_19_5_to_tile_20_5_3;
	wire vertical_tile_20_5_to_tile_19_5_0;
	wire vertical_tile_20_5_to_tile_19_5_1;
	wire vertical_tile_20_5_to_tile_19_5_2;
	wire vertical_tile_20_5_to_tile_19_5_3;

	wire vertical_tile_19_6_to_tile_20_6_0;
	wire vertical_tile_19_6_to_tile_20_6_1;
	wire vertical_tile_19_6_to_tile_20_6_2;
	wire vertical_tile_19_6_to_tile_20_6_3;
	wire vertical_tile_20_6_to_tile_19_6_0;
	wire vertical_tile_20_6_to_tile_19_6_1;
	wire vertical_tile_20_6_to_tile_19_6_2;
	wire vertical_tile_20_6_to_tile_19_6_3;

	wire vertical_tile_19_7_to_tile_20_7_0;
	wire vertical_tile_19_7_to_tile_20_7_1;
	wire vertical_tile_19_7_to_tile_20_7_2;
	wire vertical_tile_19_7_to_tile_20_7_3;
	wire vertical_tile_20_7_to_tile_19_7_0;
	wire vertical_tile_20_7_to_tile_19_7_1;
	wire vertical_tile_20_7_to_tile_19_7_2;
	wire vertical_tile_20_7_to_tile_19_7_3;

	wire vertical_tile_19_8_to_tile_20_8_0;
	wire vertical_tile_19_8_to_tile_20_8_1;
	wire vertical_tile_19_8_to_tile_20_8_2;
	wire vertical_tile_19_8_to_tile_20_8_3;
	wire vertical_tile_20_8_to_tile_19_8_0;
	wire vertical_tile_20_8_to_tile_19_8_1;
	wire vertical_tile_20_8_to_tile_19_8_2;
	wire vertical_tile_20_8_to_tile_19_8_3;

	wire vertical_tile_19_9_to_tile_20_9_0;
	wire vertical_tile_19_9_to_tile_20_9_1;
	wire vertical_tile_19_9_to_tile_20_9_2;
	wire vertical_tile_19_9_to_tile_20_9_3;
	wire vertical_tile_20_9_to_tile_19_9_0;
	wire vertical_tile_20_9_to_tile_19_9_1;
	wire vertical_tile_20_9_to_tile_19_9_2;
	wire vertical_tile_20_9_to_tile_19_9_3;

	wire vertical_tile_19_10_to_tile_20_10_0;
	wire vertical_tile_19_10_to_tile_20_10_1;
	wire vertical_tile_19_10_to_tile_20_10_2;
	wire vertical_tile_19_10_to_tile_20_10_3;
	wire vertical_tile_20_10_to_tile_19_10_0;
	wire vertical_tile_20_10_to_tile_19_10_1;
	wire vertical_tile_20_10_to_tile_19_10_2;
	wire vertical_tile_20_10_to_tile_19_10_3;

	wire vertical_tile_19_11_to_tile_20_11_0;
	wire vertical_tile_19_11_to_tile_20_11_1;
	wire vertical_tile_19_11_to_tile_20_11_2;
	wire vertical_tile_19_11_to_tile_20_11_3;
	wire vertical_tile_20_11_to_tile_19_11_0;
	wire vertical_tile_20_11_to_tile_19_11_1;
	wire vertical_tile_20_11_to_tile_19_11_2;
	wire vertical_tile_20_11_to_tile_19_11_3;

	wire vertical_tile_19_12_to_tile_20_12_0;
	wire vertical_tile_19_12_to_tile_20_12_1;
	wire vertical_tile_19_12_to_tile_20_12_2;
	wire vertical_tile_19_12_to_tile_20_12_3;
	wire vertical_tile_20_12_to_tile_19_12_0;
	wire vertical_tile_20_12_to_tile_19_12_1;
	wire vertical_tile_20_12_to_tile_19_12_2;
	wire vertical_tile_20_12_to_tile_19_12_3;

	wire vertical_tile_19_13_to_tile_20_13_0;
	wire vertical_tile_19_13_to_tile_20_13_1;
	wire vertical_tile_19_13_to_tile_20_13_2;
	wire vertical_tile_19_13_to_tile_20_13_3;
	wire vertical_tile_20_13_to_tile_19_13_0;
	wire vertical_tile_20_13_to_tile_19_13_1;
	wire vertical_tile_20_13_to_tile_19_13_2;
	wire vertical_tile_20_13_to_tile_19_13_3;

	wire vertical_tile_19_14_to_tile_20_14_0;
	wire vertical_tile_19_14_to_tile_20_14_1;
	wire vertical_tile_19_14_to_tile_20_14_2;
	wire vertical_tile_19_14_to_tile_20_14_3;
	wire vertical_tile_20_14_to_tile_19_14_0;
	wire vertical_tile_20_14_to_tile_19_14_1;
	wire vertical_tile_20_14_to_tile_19_14_2;
	wire vertical_tile_20_14_to_tile_19_14_3;

	wire vertical_tile_19_15_to_tile_20_15_0;
	wire vertical_tile_19_15_to_tile_20_15_1;
	wire vertical_tile_19_15_to_tile_20_15_2;
	wire vertical_tile_19_15_to_tile_20_15_3;
	wire vertical_tile_20_15_to_tile_19_15_0;
	wire vertical_tile_20_15_to_tile_19_15_1;
	wire vertical_tile_20_15_to_tile_19_15_2;
	wire vertical_tile_20_15_to_tile_19_15_3;

	wire vertical_tile_19_16_to_tile_20_16_0;
	wire vertical_tile_19_16_to_tile_20_16_1;
	wire vertical_tile_19_16_to_tile_20_16_2;
	wire vertical_tile_19_16_to_tile_20_16_3;
	wire vertical_tile_20_16_to_tile_19_16_0;
	wire vertical_tile_20_16_to_tile_19_16_1;
	wire vertical_tile_20_16_to_tile_19_16_2;
	wire vertical_tile_20_16_to_tile_19_16_3;

	wire vertical_tile_19_17_to_tile_20_17_0;
	wire vertical_tile_19_17_to_tile_20_17_1;
	wire vertical_tile_19_17_to_tile_20_17_2;
	wire vertical_tile_19_17_to_tile_20_17_3;
	wire vertical_tile_20_17_to_tile_19_17_0;
	wire vertical_tile_20_17_to_tile_19_17_1;
	wire vertical_tile_20_17_to_tile_19_17_2;
	wire vertical_tile_20_17_to_tile_19_17_3;

	wire vertical_tile_19_18_to_tile_20_18_0;
	wire vertical_tile_19_18_to_tile_20_18_1;
	wire vertical_tile_19_18_to_tile_20_18_2;
	wire vertical_tile_19_18_to_tile_20_18_3;
	wire vertical_tile_20_18_to_tile_19_18_0;
	wire vertical_tile_20_18_to_tile_19_18_1;
	wire vertical_tile_20_18_to_tile_19_18_2;
	wire vertical_tile_20_18_to_tile_19_18_3;

	wire vertical_tile_19_19_to_tile_20_19_0;
	wire vertical_tile_19_19_to_tile_20_19_1;
	wire vertical_tile_19_19_to_tile_20_19_2;
	wire vertical_tile_19_19_to_tile_20_19_3;
	wire vertical_tile_20_19_to_tile_19_19_0;
	wire vertical_tile_20_19_to_tile_19_19_1;
	wire vertical_tile_20_19_to_tile_19_19_2;
	wire vertical_tile_20_19_to_tile_19_19_3;

	wire vertical_tile_19_20_to_tile_20_20_0;
	wire vertical_tile_19_20_to_tile_20_20_1;
	wire vertical_tile_19_20_to_tile_20_20_2;
	wire vertical_tile_19_20_to_tile_20_20_3;
	wire vertical_tile_20_20_to_tile_19_20_0;
	wire vertical_tile_20_20_to_tile_19_20_1;
	wire vertical_tile_20_20_to_tile_19_20_2;
	wire vertical_tile_20_20_to_tile_19_20_3;

	wire vertical_tile_19_21_to_tile_20_21_0;
	wire vertical_tile_19_21_to_tile_20_21_1;
	wire vertical_tile_19_21_to_tile_20_21_2;
	wire vertical_tile_19_21_to_tile_20_21_3;
	wire vertical_tile_20_21_to_tile_19_21_0;
	wire vertical_tile_20_21_to_tile_19_21_1;
	wire vertical_tile_20_21_to_tile_19_21_2;
	wire vertical_tile_20_21_to_tile_19_21_3;

	wire vertical_tile_19_22_to_tile_20_22_0;
	wire vertical_tile_19_22_to_tile_20_22_1;
	wire vertical_tile_19_22_to_tile_20_22_2;
	wire vertical_tile_19_22_to_tile_20_22_3;
	wire vertical_tile_20_22_to_tile_19_22_0;
	wire vertical_tile_20_22_to_tile_19_22_1;
	wire vertical_tile_20_22_to_tile_19_22_2;
	wire vertical_tile_20_22_to_tile_19_22_3;

	wire vertical_tile_19_23_to_tile_20_23_0;
	wire vertical_tile_19_23_to_tile_20_23_1;
	wire vertical_tile_19_23_to_tile_20_23_2;
	wire vertical_tile_19_23_to_tile_20_23_3;
	wire vertical_tile_20_23_to_tile_19_23_0;
	wire vertical_tile_20_23_to_tile_19_23_1;
	wire vertical_tile_20_23_to_tile_19_23_2;
	wire vertical_tile_20_23_to_tile_19_23_3;

	wire vertical_tile_19_24_to_tile_20_24_0;
	wire vertical_tile_19_24_to_tile_20_24_1;
	wire vertical_tile_19_24_to_tile_20_24_2;
	wire vertical_tile_19_24_to_tile_20_24_3;
	wire vertical_tile_20_24_to_tile_19_24_0;
	wire vertical_tile_20_24_to_tile_19_24_1;
	wire vertical_tile_20_24_to_tile_19_24_2;
	wire vertical_tile_20_24_to_tile_19_24_3;

	wire vertical_tile_19_25_to_tile_20_25_0;
	wire vertical_tile_19_25_to_tile_20_25_1;
	wire vertical_tile_19_25_to_tile_20_25_2;
	wire vertical_tile_19_25_to_tile_20_25_3;
	wire vertical_tile_20_25_to_tile_19_25_0;
	wire vertical_tile_20_25_to_tile_19_25_1;
	wire vertical_tile_20_25_to_tile_19_25_2;
	wire vertical_tile_20_25_to_tile_19_25_3;

	wire vertical_tile_19_26_to_tile_20_26_0;
	wire vertical_tile_19_26_to_tile_20_26_1;
	wire vertical_tile_19_26_to_tile_20_26_2;
	wire vertical_tile_19_26_to_tile_20_26_3;
	wire vertical_tile_20_26_to_tile_19_26_0;
	wire vertical_tile_20_26_to_tile_19_26_1;
	wire vertical_tile_20_26_to_tile_19_26_2;
	wire vertical_tile_20_26_to_tile_19_26_3;

	wire vertical_tile_19_27_to_tile_20_27_0;
	wire vertical_tile_19_27_to_tile_20_27_1;
	wire vertical_tile_19_27_to_tile_20_27_2;
	wire vertical_tile_19_27_to_tile_20_27_3;
	wire vertical_tile_20_27_to_tile_19_27_0;
	wire vertical_tile_20_27_to_tile_19_27_1;
	wire vertical_tile_20_27_to_tile_19_27_2;
	wire vertical_tile_20_27_to_tile_19_27_3;

	wire vertical_tile_19_28_to_tile_20_28_0;
	wire vertical_tile_19_28_to_tile_20_28_1;
	wire vertical_tile_19_28_to_tile_20_28_2;
	wire vertical_tile_19_28_to_tile_20_28_3;
	wire vertical_tile_20_28_to_tile_19_28_0;
	wire vertical_tile_20_28_to_tile_19_28_1;
	wire vertical_tile_20_28_to_tile_19_28_2;
	wire vertical_tile_20_28_to_tile_19_28_3;

	wire vertical_tile_19_29_to_tile_20_29_0;
	wire vertical_tile_19_29_to_tile_20_29_1;
	wire vertical_tile_19_29_to_tile_20_29_2;
	wire vertical_tile_19_29_to_tile_20_29_3;
	wire vertical_tile_20_29_to_tile_19_29_0;
	wire vertical_tile_20_29_to_tile_19_29_1;
	wire vertical_tile_20_29_to_tile_19_29_2;
	wire vertical_tile_20_29_to_tile_19_29_3;

	wire vertical_tile_19_30_to_tile_20_30_0;
	wire vertical_tile_19_30_to_tile_20_30_1;
	wire vertical_tile_19_30_to_tile_20_30_2;
	wire vertical_tile_19_30_to_tile_20_30_3;
	wire vertical_tile_20_30_to_tile_19_30_0;
	wire vertical_tile_20_30_to_tile_19_30_1;
	wire vertical_tile_20_30_to_tile_19_30_2;
	wire vertical_tile_20_30_to_tile_19_30_3;

	wire vertical_tile_19_31_to_tile_20_31_0;
	wire vertical_tile_19_31_to_tile_20_31_1;
	wire vertical_tile_19_31_to_tile_20_31_2;
	wire vertical_tile_19_31_to_tile_20_31_3;
	wire vertical_tile_20_31_to_tile_19_31_0;
	wire vertical_tile_20_31_to_tile_19_31_1;
	wire vertical_tile_20_31_to_tile_19_31_2;
	wire vertical_tile_20_31_to_tile_19_31_3;

	wire vertical_tile_20_0_to_tile_21_0_0;
	wire vertical_tile_20_0_to_tile_21_0_1;
	wire vertical_tile_20_0_to_tile_21_0_2;
	wire vertical_tile_20_0_to_tile_21_0_3;
	wire vertical_tile_21_0_to_tile_20_0_0;
	wire vertical_tile_21_0_to_tile_20_0_1;
	wire vertical_tile_21_0_to_tile_20_0_2;
	wire vertical_tile_21_0_to_tile_20_0_3;

	wire vertical_tile_20_1_to_tile_21_1_0;
	wire vertical_tile_20_1_to_tile_21_1_1;
	wire vertical_tile_20_1_to_tile_21_1_2;
	wire vertical_tile_20_1_to_tile_21_1_3;
	wire vertical_tile_21_1_to_tile_20_1_0;
	wire vertical_tile_21_1_to_tile_20_1_1;
	wire vertical_tile_21_1_to_tile_20_1_2;
	wire vertical_tile_21_1_to_tile_20_1_3;

	wire vertical_tile_20_2_to_tile_21_2_0;
	wire vertical_tile_20_2_to_tile_21_2_1;
	wire vertical_tile_20_2_to_tile_21_2_2;
	wire vertical_tile_20_2_to_tile_21_2_3;
	wire vertical_tile_21_2_to_tile_20_2_0;
	wire vertical_tile_21_2_to_tile_20_2_1;
	wire vertical_tile_21_2_to_tile_20_2_2;
	wire vertical_tile_21_2_to_tile_20_2_3;

	wire vertical_tile_20_3_to_tile_21_3_0;
	wire vertical_tile_20_3_to_tile_21_3_1;
	wire vertical_tile_20_3_to_tile_21_3_2;
	wire vertical_tile_20_3_to_tile_21_3_3;
	wire vertical_tile_21_3_to_tile_20_3_0;
	wire vertical_tile_21_3_to_tile_20_3_1;
	wire vertical_tile_21_3_to_tile_20_3_2;
	wire vertical_tile_21_3_to_tile_20_3_3;

	wire vertical_tile_20_4_to_tile_21_4_0;
	wire vertical_tile_20_4_to_tile_21_4_1;
	wire vertical_tile_20_4_to_tile_21_4_2;
	wire vertical_tile_20_4_to_tile_21_4_3;
	wire vertical_tile_21_4_to_tile_20_4_0;
	wire vertical_tile_21_4_to_tile_20_4_1;
	wire vertical_tile_21_4_to_tile_20_4_2;
	wire vertical_tile_21_4_to_tile_20_4_3;

	wire vertical_tile_20_5_to_tile_21_5_0;
	wire vertical_tile_20_5_to_tile_21_5_1;
	wire vertical_tile_20_5_to_tile_21_5_2;
	wire vertical_tile_20_5_to_tile_21_5_3;
	wire vertical_tile_21_5_to_tile_20_5_0;
	wire vertical_tile_21_5_to_tile_20_5_1;
	wire vertical_tile_21_5_to_tile_20_5_2;
	wire vertical_tile_21_5_to_tile_20_5_3;

	wire vertical_tile_20_6_to_tile_21_6_0;
	wire vertical_tile_20_6_to_tile_21_6_1;
	wire vertical_tile_20_6_to_tile_21_6_2;
	wire vertical_tile_20_6_to_tile_21_6_3;
	wire vertical_tile_21_6_to_tile_20_6_0;
	wire vertical_tile_21_6_to_tile_20_6_1;
	wire vertical_tile_21_6_to_tile_20_6_2;
	wire vertical_tile_21_6_to_tile_20_6_3;

	wire vertical_tile_20_7_to_tile_21_7_0;
	wire vertical_tile_20_7_to_tile_21_7_1;
	wire vertical_tile_20_7_to_tile_21_7_2;
	wire vertical_tile_20_7_to_tile_21_7_3;
	wire vertical_tile_21_7_to_tile_20_7_0;
	wire vertical_tile_21_7_to_tile_20_7_1;
	wire vertical_tile_21_7_to_tile_20_7_2;
	wire vertical_tile_21_7_to_tile_20_7_3;

	wire vertical_tile_20_8_to_tile_21_8_0;
	wire vertical_tile_20_8_to_tile_21_8_1;
	wire vertical_tile_20_8_to_tile_21_8_2;
	wire vertical_tile_20_8_to_tile_21_8_3;
	wire vertical_tile_21_8_to_tile_20_8_0;
	wire vertical_tile_21_8_to_tile_20_8_1;
	wire vertical_tile_21_8_to_tile_20_8_2;
	wire vertical_tile_21_8_to_tile_20_8_3;

	wire vertical_tile_20_9_to_tile_21_9_0;
	wire vertical_tile_20_9_to_tile_21_9_1;
	wire vertical_tile_20_9_to_tile_21_9_2;
	wire vertical_tile_20_9_to_tile_21_9_3;
	wire vertical_tile_21_9_to_tile_20_9_0;
	wire vertical_tile_21_9_to_tile_20_9_1;
	wire vertical_tile_21_9_to_tile_20_9_2;
	wire vertical_tile_21_9_to_tile_20_9_3;

	wire vertical_tile_20_10_to_tile_21_10_0;
	wire vertical_tile_20_10_to_tile_21_10_1;
	wire vertical_tile_20_10_to_tile_21_10_2;
	wire vertical_tile_20_10_to_tile_21_10_3;
	wire vertical_tile_21_10_to_tile_20_10_0;
	wire vertical_tile_21_10_to_tile_20_10_1;
	wire vertical_tile_21_10_to_tile_20_10_2;
	wire vertical_tile_21_10_to_tile_20_10_3;

	wire vertical_tile_20_11_to_tile_21_11_0;
	wire vertical_tile_20_11_to_tile_21_11_1;
	wire vertical_tile_20_11_to_tile_21_11_2;
	wire vertical_tile_20_11_to_tile_21_11_3;
	wire vertical_tile_21_11_to_tile_20_11_0;
	wire vertical_tile_21_11_to_tile_20_11_1;
	wire vertical_tile_21_11_to_tile_20_11_2;
	wire vertical_tile_21_11_to_tile_20_11_3;

	wire vertical_tile_20_12_to_tile_21_12_0;
	wire vertical_tile_20_12_to_tile_21_12_1;
	wire vertical_tile_20_12_to_tile_21_12_2;
	wire vertical_tile_20_12_to_tile_21_12_3;
	wire vertical_tile_21_12_to_tile_20_12_0;
	wire vertical_tile_21_12_to_tile_20_12_1;
	wire vertical_tile_21_12_to_tile_20_12_2;
	wire vertical_tile_21_12_to_tile_20_12_3;

	wire vertical_tile_20_13_to_tile_21_13_0;
	wire vertical_tile_20_13_to_tile_21_13_1;
	wire vertical_tile_20_13_to_tile_21_13_2;
	wire vertical_tile_20_13_to_tile_21_13_3;
	wire vertical_tile_21_13_to_tile_20_13_0;
	wire vertical_tile_21_13_to_tile_20_13_1;
	wire vertical_tile_21_13_to_tile_20_13_2;
	wire vertical_tile_21_13_to_tile_20_13_3;

	wire vertical_tile_20_14_to_tile_21_14_0;
	wire vertical_tile_20_14_to_tile_21_14_1;
	wire vertical_tile_20_14_to_tile_21_14_2;
	wire vertical_tile_20_14_to_tile_21_14_3;
	wire vertical_tile_21_14_to_tile_20_14_0;
	wire vertical_tile_21_14_to_tile_20_14_1;
	wire vertical_tile_21_14_to_tile_20_14_2;
	wire vertical_tile_21_14_to_tile_20_14_3;

	wire vertical_tile_20_15_to_tile_21_15_0;
	wire vertical_tile_20_15_to_tile_21_15_1;
	wire vertical_tile_20_15_to_tile_21_15_2;
	wire vertical_tile_20_15_to_tile_21_15_3;
	wire vertical_tile_21_15_to_tile_20_15_0;
	wire vertical_tile_21_15_to_tile_20_15_1;
	wire vertical_tile_21_15_to_tile_20_15_2;
	wire vertical_tile_21_15_to_tile_20_15_3;

	wire vertical_tile_20_16_to_tile_21_16_0;
	wire vertical_tile_20_16_to_tile_21_16_1;
	wire vertical_tile_20_16_to_tile_21_16_2;
	wire vertical_tile_20_16_to_tile_21_16_3;
	wire vertical_tile_21_16_to_tile_20_16_0;
	wire vertical_tile_21_16_to_tile_20_16_1;
	wire vertical_tile_21_16_to_tile_20_16_2;
	wire vertical_tile_21_16_to_tile_20_16_3;

	wire vertical_tile_20_17_to_tile_21_17_0;
	wire vertical_tile_20_17_to_tile_21_17_1;
	wire vertical_tile_20_17_to_tile_21_17_2;
	wire vertical_tile_20_17_to_tile_21_17_3;
	wire vertical_tile_21_17_to_tile_20_17_0;
	wire vertical_tile_21_17_to_tile_20_17_1;
	wire vertical_tile_21_17_to_tile_20_17_2;
	wire vertical_tile_21_17_to_tile_20_17_3;

	wire vertical_tile_20_18_to_tile_21_18_0;
	wire vertical_tile_20_18_to_tile_21_18_1;
	wire vertical_tile_20_18_to_tile_21_18_2;
	wire vertical_tile_20_18_to_tile_21_18_3;
	wire vertical_tile_21_18_to_tile_20_18_0;
	wire vertical_tile_21_18_to_tile_20_18_1;
	wire vertical_tile_21_18_to_tile_20_18_2;
	wire vertical_tile_21_18_to_tile_20_18_3;

	wire vertical_tile_20_19_to_tile_21_19_0;
	wire vertical_tile_20_19_to_tile_21_19_1;
	wire vertical_tile_20_19_to_tile_21_19_2;
	wire vertical_tile_20_19_to_tile_21_19_3;
	wire vertical_tile_21_19_to_tile_20_19_0;
	wire vertical_tile_21_19_to_tile_20_19_1;
	wire vertical_tile_21_19_to_tile_20_19_2;
	wire vertical_tile_21_19_to_tile_20_19_3;

	wire vertical_tile_20_20_to_tile_21_20_0;
	wire vertical_tile_20_20_to_tile_21_20_1;
	wire vertical_tile_20_20_to_tile_21_20_2;
	wire vertical_tile_20_20_to_tile_21_20_3;
	wire vertical_tile_21_20_to_tile_20_20_0;
	wire vertical_tile_21_20_to_tile_20_20_1;
	wire vertical_tile_21_20_to_tile_20_20_2;
	wire vertical_tile_21_20_to_tile_20_20_3;

	wire vertical_tile_20_21_to_tile_21_21_0;
	wire vertical_tile_20_21_to_tile_21_21_1;
	wire vertical_tile_20_21_to_tile_21_21_2;
	wire vertical_tile_20_21_to_tile_21_21_3;
	wire vertical_tile_21_21_to_tile_20_21_0;
	wire vertical_tile_21_21_to_tile_20_21_1;
	wire vertical_tile_21_21_to_tile_20_21_2;
	wire vertical_tile_21_21_to_tile_20_21_3;

	wire vertical_tile_20_22_to_tile_21_22_0;
	wire vertical_tile_20_22_to_tile_21_22_1;
	wire vertical_tile_20_22_to_tile_21_22_2;
	wire vertical_tile_20_22_to_tile_21_22_3;
	wire vertical_tile_21_22_to_tile_20_22_0;
	wire vertical_tile_21_22_to_tile_20_22_1;
	wire vertical_tile_21_22_to_tile_20_22_2;
	wire vertical_tile_21_22_to_tile_20_22_3;

	wire vertical_tile_20_23_to_tile_21_23_0;
	wire vertical_tile_20_23_to_tile_21_23_1;
	wire vertical_tile_20_23_to_tile_21_23_2;
	wire vertical_tile_20_23_to_tile_21_23_3;
	wire vertical_tile_21_23_to_tile_20_23_0;
	wire vertical_tile_21_23_to_tile_20_23_1;
	wire vertical_tile_21_23_to_tile_20_23_2;
	wire vertical_tile_21_23_to_tile_20_23_3;

	wire vertical_tile_20_24_to_tile_21_24_0;
	wire vertical_tile_20_24_to_tile_21_24_1;
	wire vertical_tile_20_24_to_tile_21_24_2;
	wire vertical_tile_20_24_to_tile_21_24_3;
	wire vertical_tile_21_24_to_tile_20_24_0;
	wire vertical_tile_21_24_to_tile_20_24_1;
	wire vertical_tile_21_24_to_tile_20_24_2;
	wire vertical_tile_21_24_to_tile_20_24_3;

	wire vertical_tile_20_25_to_tile_21_25_0;
	wire vertical_tile_20_25_to_tile_21_25_1;
	wire vertical_tile_20_25_to_tile_21_25_2;
	wire vertical_tile_20_25_to_tile_21_25_3;
	wire vertical_tile_21_25_to_tile_20_25_0;
	wire vertical_tile_21_25_to_tile_20_25_1;
	wire vertical_tile_21_25_to_tile_20_25_2;
	wire vertical_tile_21_25_to_tile_20_25_3;

	wire vertical_tile_20_26_to_tile_21_26_0;
	wire vertical_tile_20_26_to_tile_21_26_1;
	wire vertical_tile_20_26_to_tile_21_26_2;
	wire vertical_tile_20_26_to_tile_21_26_3;
	wire vertical_tile_21_26_to_tile_20_26_0;
	wire vertical_tile_21_26_to_tile_20_26_1;
	wire vertical_tile_21_26_to_tile_20_26_2;
	wire vertical_tile_21_26_to_tile_20_26_3;

	wire vertical_tile_20_27_to_tile_21_27_0;
	wire vertical_tile_20_27_to_tile_21_27_1;
	wire vertical_tile_20_27_to_tile_21_27_2;
	wire vertical_tile_20_27_to_tile_21_27_3;
	wire vertical_tile_21_27_to_tile_20_27_0;
	wire vertical_tile_21_27_to_tile_20_27_1;
	wire vertical_tile_21_27_to_tile_20_27_2;
	wire vertical_tile_21_27_to_tile_20_27_3;

	wire vertical_tile_20_28_to_tile_21_28_0;
	wire vertical_tile_20_28_to_tile_21_28_1;
	wire vertical_tile_20_28_to_tile_21_28_2;
	wire vertical_tile_20_28_to_tile_21_28_3;
	wire vertical_tile_21_28_to_tile_20_28_0;
	wire vertical_tile_21_28_to_tile_20_28_1;
	wire vertical_tile_21_28_to_tile_20_28_2;
	wire vertical_tile_21_28_to_tile_20_28_3;

	wire vertical_tile_20_29_to_tile_21_29_0;
	wire vertical_tile_20_29_to_tile_21_29_1;
	wire vertical_tile_20_29_to_tile_21_29_2;
	wire vertical_tile_20_29_to_tile_21_29_3;
	wire vertical_tile_21_29_to_tile_20_29_0;
	wire vertical_tile_21_29_to_tile_20_29_1;
	wire vertical_tile_21_29_to_tile_20_29_2;
	wire vertical_tile_21_29_to_tile_20_29_3;

	wire vertical_tile_20_30_to_tile_21_30_0;
	wire vertical_tile_20_30_to_tile_21_30_1;
	wire vertical_tile_20_30_to_tile_21_30_2;
	wire vertical_tile_20_30_to_tile_21_30_3;
	wire vertical_tile_21_30_to_tile_20_30_0;
	wire vertical_tile_21_30_to_tile_20_30_1;
	wire vertical_tile_21_30_to_tile_20_30_2;
	wire vertical_tile_21_30_to_tile_20_30_3;

	wire vertical_tile_20_31_to_tile_21_31_0;
	wire vertical_tile_20_31_to_tile_21_31_1;
	wire vertical_tile_20_31_to_tile_21_31_2;
	wire vertical_tile_20_31_to_tile_21_31_3;
	wire vertical_tile_21_31_to_tile_20_31_0;
	wire vertical_tile_21_31_to_tile_20_31_1;
	wire vertical_tile_21_31_to_tile_20_31_2;
	wire vertical_tile_21_31_to_tile_20_31_3;

	wire vertical_tile_21_0_to_tile_22_0_0;
	wire vertical_tile_21_0_to_tile_22_0_1;
	wire vertical_tile_21_0_to_tile_22_0_2;
	wire vertical_tile_21_0_to_tile_22_0_3;
	wire vertical_tile_22_0_to_tile_21_0_0;
	wire vertical_tile_22_0_to_tile_21_0_1;
	wire vertical_tile_22_0_to_tile_21_0_2;
	wire vertical_tile_22_0_to_tile_21_0_3;

	wire vertical_tile_21_1_to_tile_22_1_0;
	wire vertical_tile_21_1_to_tile_22_1_1;
	wire vertical_tile_21_1_to_tile_22_1_2;
	wire vertical_tile_21_1_to_tile_22_1_3;
	wire vertical_tile_22_1_to_tile_21_1_0;
	wire vertical_tile_22_1_to_tile_21_1_1;
	wire vertical_tile_22_1_to_tile_21_1_2;
	wire vertical_tile_22_1_to_tile_21_1_3;

	wire vertical_tile_21_2_to_tile_22_2_0;
	wire vertical_tile_21_2_to_tile_22_2_1;
	wire vertical_tile_21_2_to_tile_22_2_2;
	wire vertical_tile_21_2_to_tile_22_2_3;
	wire vertical_tile_22_2_to_tile_21_2_0;
	wire vertical_tile_22_2_to_tile_21_2_1;
	wire vertical_tile_22_2_to_tile_21_2_2;
	wire vertical_tile_22_2_to_tile_21_2_3;

	wire vertical_tile_21_3_to_tile_22_3_0;
	wire vertical_tile_21_3_to_tile_22_3_1;
	wire vertical_tile_21_3_to_tile_22_3_2;
	wire vertical_tile_21_3_to_tile_22_3_3;
	wire vertical_tile_22_3_to_tile_21_3_0;
	wire vertical_tile_22_3_to_tile_21_3_1;
	wire vertical_tile_22_3_to_tile_21_3_2;
	wire vertical_tile_22_3_to_tile_21_3_3;

	wire vertical_tile_21_4_to_tile_22_4_0;
	wire vertical_tile_21_4_to_tile_22_4_1;
	wire vertical_tile_21_4_to_tile_22_4_2;
	wire vertical_tile_21_4_to_tile_22_4_3;
	wire vertical_tile_22_4_to_tile_21_4_0;
	wire vertical_tile_22_4_to_tile_21_4_1;
	wire vertical_tile_22_4_to_tile_21_4_2;
	wire vertical_tile_22_4_to_tile_21_4_3;

	wire vertical_tile_21_5_to_tile_22_5_0;
	wire vertical_tile_21_5_to_tile_22_5_1;
	wire vertical_tile_21_5_to_tile_22_5_2;
	wire vertical_tile_21_5_to_tile_22_5_3;
	wire vertical_tile_22_5_to_tile_21_5_0;
	wire vertical_tile_22_5_to_tile_21_5_1;
	wire vertical_tile_22_5_to_tile_21_5_2;
	wire vertical_tile_22_5_to_tile_21_5_3;

	wire vertical_tile_21_6_to_tile_22_6_0;
	wire vertical_tile_21_6_to_tile_22_6_1;
	wire vertical_tile_21_6_to_tile_22_6_2;
	wire vertical_tile_21_6_to_tile_22_6_3;
	wire vertical_tile_22_6_to_tile_21_6_0;
	wire vertical_tile_22_6_to_tile_21_6_1;
	wire vertical_tile_22_6_to_tile_21_6_2;
	wire vertical_tile_22_6_to_tile_21_6_3;

	wire vertical_tile_21_7_to_tile_22_7_0;
	wire vertical_tile_21_7_to_tile_22_7_1;
	wire vertical_tile_21_7_to_tile_22_7_2;
	wire vertical_tile_21_7_to_tile_22_7_3;
	wire vertical_tile_22_7_to_tile_21_7_0;
	wire vertical_tile_22_7_to_tile_21_7_1;
	wire vertical_tile_22_7_to_tile_21_7_2;
	wire vertical_tile_22_7_to_tile_21_7_3;

	wire vertical_tile_21_8_to_tile_22_8_0;
	wire vertical_tile_21_8_to_tile_22_8_1;
	wire vertical_tile_21_8_to_tile_22_8_2;
	wire vertical_tile_21_8_to_tile_22_8_3;
	wire vertical_tile_22_8_to_tile_21_8_0;
	wire vertical_tile_22_8_to_tile_21_8_1;
	wire vertical_tile_22_8_to_tile_21_8_2;
	wire vertical_tile_22_8_to_tile_21_8_3;

	wire vertical_tile_21_9_to_tile_22_9_0;
	wire vertical_tile_21_9_to_tile_22_9_1;
	wire vertical_tile_21_9_to_tile_22_9_2;
	wire vertical_tile_21_9_to_tile_22_9_3;
	wire vertical_tile_22_9_to_tile_21_9_0;
	wire vertical_tile_22_9_to_tile_21_9_1;
	wire vertical_tile_22_9_to_tile_21_9_2;
	wire vertical_tile_22_9_to_tile_21_9_3;

	wire vertical_tile_21_10_to_tile_22_10_0;
	wire vertical_tile_21_10_to_tile_22_10_1;
	wire vertical_tile_21_10_to_tile_22_10_2;
	wire vertical_tile_21_10_to_tile_22_10_3;
	wire vertical_tile_22_10_to_tile_21_10_0;
	wire vertical_tile_22_10_to_tile_21_10_1;
	wire vertical_tile_22_10_to_tile_21_10_2;
	wire vertical_tile_22_10_to_tile_21_10_3;

	wire vertical_tile_21_11_to_tile_22_11_0;
	wire vertical_tile_21_11_to_tile_22_11_1;
	wire vertical_tile_21_11_to_tile_22_11_2;
	wire vertical_tile_21_11_to_tile_22_11_3;
	wire vertical_tile_22_11_to_tile_21_11_0;
	wire vertical_tile_22_11_to_tile_21_11_1;
	wire vertical_tile_22_11_to_tile_21_11_2;
	wire vertical_tile_22_11_to_tile_21_11_3;

	wire vertical_tile_21_12_to_tile_22_12_0;
	wire vertical_tile_21_12_to_tile_22_12_1;
	wire vertical_tile_21_12_to_tile_22_12_2;
	wire vertical_tile_21_12_to_tile_22_12_3;
	wire vertical_tile_22_12_to_tile_21_12_0;
	wire vertical_tile_22_12_to_tile_21_12_1;
	wire vertical_tile_22_12_to_tile_21_12_2;
	wire vertical_tile_22_12_to_tile_21_12_3;

	wire vertical_tile_21_13_to_tile_22_13_0;
	wire vertical_tile_21_13_to_tile_22_13_1;
	wire vertical_tile_21_13_to_tile_22_13_2;
	wire vertical_tile_21_13_to_tile_22_13_3;
	wire vertical_tile_22_13_to_tile_21_13_0;
	wire vertical_tile_22_13_to_tile_21_13_1;
	wire vertical_tile_22_13_to_tile_21_13_2;
	wire vertical_tile_22_13_to_tile_21_13_3;

	wire vertical_tile_21_14_to_tile_22_14_0;
	wire vertical_tile_21_14_to_tile_22_14_1;
	wire vertical_tile_21_14_to_tile_22_14_2;
	wire vertical_tile_21_14_to_tile_22_14_3;
	wire vertical_tile_22_14_to_tile_21_14_0;
	wire vertical_tile_22_14_to_tile_21_14_1;
	wire vertical_tile_22_14_to_tile_21_14_2;
	wire vertical_tile_22_14_to_tile_21_14_3;

	wire vertical_tile_21_15_to_tile_22_15_0;
	wire vertical_tile_21_15_to_tile_22_15_1;
	wire vertical_tile_21_15_to_tile_22_15_2;
	wire vertical_tile_21_15_to_tile_22_15_3;
	wire vertical_tile_22_15_to_tile_21_15_0;
	wire vertical_tile_22_15_to_tile_21_15_1;
	wire vertical_tile_22_15_to_tile_21_15_2;
	wire vertical_tile_22_15_to_tile_21_15_3;

	wire vertical_tile_21_16_to_tile_22_16_0;
	wire vertical_tile_21_16_to_tile_22_16_1;
	wire vertical_tile_21_16_to_tile_22_16_2;
	wire vertical_tile_21_16_to_tile_22_16_3;
	wire vertical_tile_22_16_to_tile_21_16_0;
	wire vertical_tile_22_16_to_tile_21_16_1;
	wire vertical_tile_22_16_to_tile_21_16_2;
	wire vertical_tile_22_16_to_tile_21_16_3;

	wire vertical_tile_21_17_to_tile_22_17_0;
	wire vertical_tile_21_17_to_tile_22_17_1;
	wire vertical_tile_21_17_to_tile_22_17_2;
	wire vertical_tile_21_17_to_tile_22_17_3;
	wire vertical_tile_22_17_to_tile_21_17_0;
	wire vertical_tile_22_17_to_tile_21_17_1;
	wire vertical_tile_22_17_to_tile_21_17_2;
	wire vertical_tile_22_17_to_tile_21_17_3;

	wire vertical_tile_21_18_to_tile_22_18_0;
	wire vertical_tile_21_18_to_tile_22_18_1;
	wire vertical_tile_21_18_to_tile_22_18_2;
	wire vertical_tile_21_18_to_tile_22_18_3;
	wire vertical_tile_22_18_to_tile_21_18_0;
	wire vertical_tile_22_18_to_tile_21_18_1;
	wire vertical_tile_22_18_to_tile_21_18_2;
	wire vertical_tile_22_18_to_tile_21_18_3;

	wire vertical_tile_21_19_to_tile_22_19_0;
	wire vertical_tile_21_19_to_tile_22_19_1;
	wire vertical_tile_21_19_to_tile_22_19_2;
	wire vertical_tile_21_19_to_tile_22_19_3;
	wire vertical_tile_22_19_to_tile_21_19_0;
	wire vertical_tile_22_19_to_tile_21_19_1;
	wire vertical_tile_22_19_to_tile_21_19_2;
	wire vertical_tile_22_19_to_tile_21_19_3;

	wire vertical_tile_21_20_to_tile_22_20_0;
	wire vertical_tile_21_20_to_tile_22_20_1;
	wire vertical_tile_21_20_to_tile_22_20_2;
	wire vertical_tile_21_20_to_tile_22_20_3;
	wire vertical_tile_22_20_to_tile_21_20_0;
	wire vertical_tile_22_20_to_tile_21_20_1;
	wire vertical_tile_22_20_to_tile_21_20_2;
	wire vertical_tile_22_20_to_tile_21_20_3;

	wire vertical_tile_21_21_to_tile_22_21_0;
	wire vertical_tile_21_21_to_tile_22_21_1;
	wire vertical_tile_21_21_to_tile_22_21_2;
	wire vertical_tile_21_21_to_tile_22_21_3;
	wire vertical_tile_22_21_to_tile_21_21_0;
	wire vertical_tile_22_21_to_tile_21_21_1;
	wire vertical_tile_22_21_to_tile_21_21_2;
	wire vertical_tile_22_21_to_tile_21_21_3;

	wire vertical_tile_21_22_to_tile_22_22_0;
	wire vertical_tile_21_22_to_tile_22_22_1;
	wire vertical_tile_21_22_to_tile_22_22_2;
	wire vertical_tile_21_22_to_tile_22_22_3;
	wire vertical_tile_22_22_to_tile_21_22_0;
	wire vertical_tile_22_22_to_tile_21_22_1;
	wire vertical_tile_22_22_to_tile_21_22_2;
	wire vertical_tile_22_22_to_tile_21_22_3;

	wire vertical_tile_21_23_to_tile_22_23_0;
	wire vertical_tile_21_23_to_tile_22_23_1;
	wire vertical_tile_21_23_to_tile_22_23_2;
	wire vertical_tile_21_23_to_tile_22_23_3;
	wire vertical_tile_22_23_to_tile_21_23_0;
	wire vertical_tile_22_23_to_tile_21_23_1;
	wire vertical_tile_22_23_to_tile_21_23_2;
	wire vertical_tile_22_23_to_tile_21_23_3;

	wire vertical_tile_21_24_to_tile_22_24_0;
	wire vertical_tile_21_24_to_tile_22_24_1;
	wire vertical_tile_21_24_to_tile_22_24_2;
	wire vertical_tile_21_24_to_tile_22_24_3;
	wire vertical_tile_22_24_to_tile_21_24_0;
	wire vertical_tile_22_24_to_tile_21_24_1;
	wire vertical_tile_22_24_to_tile_21_24_2;
	wire vertical_tile_22_24_to_tile_21_24_3;

	wire vertical_tile_21_25_to_tile_22_25_0;
	wire vertical_tile_21_25_to_tile_22_25_1;
	wire vertical_tile_21_25_to_tile_22_25_2;
	wire vertical_tile_21_25_to_tile_22_25_3;
	wire vertical_tile_22_25_to_tile_21_25_0;
	wire vertical_tile_22_25_to_tile_21_25_1;
	wire vertical_tile_22_25_to_tile_21_25_2;
	wire vertical_tile_22_25_to_tile_21_25_3;

	wire vertical_tile_21_26_to_tile_22_26_0;
	wire vertical_tile_21_26_to_tile_22_26_1;
	wire vertical_tile_21_26_to_tile_22_26_2;
	wire vertical_tile_21_26_to_tile_22_26_3;
	wire vertical_tile_22_26_to_tile_21_26_0;
	wire vertical_tile_22_26_to_tile_21_26_1;
	wire vertical_tile_22_26_to_tile_21_26_2;
	wire vertical_tile_22_26_to_tile_21_26_3;

	wire vertical_tile_21_27_to_tile_22_27_0;
	wire vertical_tile_21_27_to_tile_22_27_1;
	wire vertical_tile_21_27_to_tile_22_27_2;
	wire vertical_tile_21_27_to_tile_22_27_3;
	wire vertical_tile_22_27_to_tile_21_27_0;
	wire vertical_tile_22_27_to_tile_21_27_1;
	wire vertical_tile_22_27_to_tile_21_27_2;
	wire vertical_tile_22_27_to_tile_21_27_3;

	wire vertical_tile_21_28_to_tile_22_28_0;
	wire vertical_tile_21_28_to_tile_22_28_1;
	wire vertical_tile_21_28_to_tile_22_28_2;
	wire vertical_tile_21_28_to_tile_22_28_3;
	wire vertical_tile_22_28_to_tile_21_28_0;
	wire vertical_tile_22_28_to_tile_21_28_1;
	wire vertical_tile_22_28_to_tile_21_28_2;
	wire vertical_tile_22_28_to_tile_21_28_3;

	wire vertical_tile_21_29_to_tile_22_29_0;
	wire vertical_tile_21_29_to_tile_22_29_1;
	wire vertical_tile_21_29_to_tile_22_29_2;
	wire vertical_tile_21_29_to_tile_22_29_3;
	wire vertical_tile_22_29_to_tile_21_29_0;
	wire vertical_tile_22_29_to_tile_21_29_1;
	wire vertical_tile_22_29_to_tile_21_29_2;
	wire vertical_tile_22_29_to_tile_21_29_3;

	wire vertical_tile_21_30_to_tile_22_30_0;
	wire vertical_tile_21_30_to_tile_22_30_1;
	wire vertical_tile_21_30_to_tile_22_30_2;
	wire vertical_tile_21_30_to_tile_22_30_3;
	wire vertical_tile_22_30_to_tile_21_30_0;
	wire vertical_tile_22_30_to_tile_21_30_1;
	wire vertical_tile_22_30_to_tile_21_30_2;
	wire vertical_tile_22_30_to_tile_21_30_3;

	wire vertical_tile_21_31_to_tile_22_31_0;
	wire vertical_tile_21_31_to_tile_22_31_1;
	wire vertical_tile_21_31_to_tile_22_31_2;
	wire vertical_tile_21_31_to_tile_22_31_3;
	wire vertical_tile_22_31_to_tile_21_31_0;
	wire vertical_tile_22_31_to_tile_21_31_1;
	wire vertical_tile_22_31_to_tile_21_31_2;
	wire vertical_tile_22_31_to_tile_21_31_3;

	wire vertical_tile_22_0_to_tile_23_0_0;
	wire vertical_tile_22_0_to_tile_23_0_1;
	wire vertical_tile_22_0_to_tile_23_0_2;
	wire vertical_tile_22_0_to_tile_23_0_3;
	wire vertical_tile_23_0_to_tile_22_0_0;
	wire vertical_tile_23_0_to_tile_22_0_1;
	wire vertical_tile_23_0_to_tile_22_0_2;
	wire vertical_tile_23_0_to_tile_22_0_3;

	wire vertical_tile_22_1_to_tile_23_1_0;
	wire vertical_tile_22_1_to_tile_23_1_1;
	wire vertical_tile_22_1_to_tile_23_1_2;
	wire vertical_tile_22_1_to_tile_23_1_3;
	wire vertical_tile_23_1_to_tile_22_1_0;
	wire vertical_tile_23_1_to_tile_22_1_1;
	wire vertical_tile_23_1_to_tile_22_1_2;
	wire vertical_tile_23_1_to_tile_22_1_3;

	wire vertical_tile_22_2_to_tile_23_2_0;
	wire vertical_tile_22_2_to_tile_23_2_1;
	wire vertical_tile_22_2_to_tile_23_2_2;
	wire vertical_tile_22_2_to_tile_23_2_3;
	wire vertical_tile_23_2_to_tile_22_2_0;
	wire vertical_tile_23_2_to_tile_22_2_1;
	wire vertical_tile_23_2_to_tile_22_2_2;
	wire vertical_tile_23_2_to_tile_22_2_3;

	wire vertical_tile_22_3_to_tile_23_3_0;
	wire vertical_tile_22_3_to_tile_23_3_1;
	wire vertical_tile_22_3_to_tile_23_3_2;
	wire vertical_tile_22_3_to_tile_23_3_3;
	wire vertical_tile_23_3_to_tile_22_3_0;
	wire vertical_tile_23_3_to_tile_22_3_1;
	wire vertical_tile_23_3_to_tile_22_3_2;
	wire vertical_tile_23_3_to_tile_22_3_3;

	wire vertical_tile_22_4_to_tile_23_4_0;
	wire vertical_tile_22_4_to_tile_23_4_1;
	wire vertical_tile_22_4_to_tile_23_4_2;
	wire vertical_tile_22_4_to_tile_23_4_3;
	wire vertical_tile_23_4_to_tile_22_4_0;
	wire vertical_tile_23_4_to_tile_22_4_1;
	wire vertical_tile_23_4_to_tile_22_4_2;
	wire vertical_tile_23_4_to_tile_22_4_3;

	wire vertical_tile_22_5_to_tile_23_5_0;
	wire vertical_tile_22_5_to_tile_23_5_1;
	wire vertical_tile_22_5_to_tile_23_5_2;
	wire vertical_tile_22_5_to_tile_23_5_3;
	wire vertical_tile_23_5_to_tile_22_5_0;
	wire vertical_tile_23_5_to_tile_22_5_1;
	wire vertical_tile_23_5_to_tile_22_5_2;
	wire vertical_tile_23_5_to_tile_22_5_3;

	wire vertical_tile_22_6_to_tile_23_6_0;
	wire vertical_tile_22_6_to_tile_23_6_1;
	wire vertical_tile_22_6_to_tile_23_6_2;
	wire vertical_tile_22_6_to_tile_23_6_3;
	wire vertical_tile_23_6_to_tile_22_6_0;
	wire vertical_tile_23_6_to_tile_22_6_1;
	wire vertical_tile_23_6_to_tile_22_6_2;
	wire vertical_tile_23_6_to_tile_22_6_3;

	wire vertical_tile_22_7_to_tile_23_7_0;
	wire vertical_tile_22_7_to_tile_23_7_1;
	wire vertical_tile_22_7_to_tile_23_7_2;
	wire vertical_tile_22_7_to_tile_23_7_3;
	wire vertical_tile_23_7_to_tile_22_7_0;
	wire vertical_tile_23_7_to_tile_22_7_1;
	wire vertical_tile_23_7_to_tile_22_7_2;
	wire vertical_tile_23_7_to_tile_22_7_3;

	wire vertical_tile_22_8_to_tile_23_8_0;
	wire vertical_tile_22_8_to_tile_23_8_1;
	wire vertical_tile_22_8_to_tile_23_8_2;
	wire vertical_tile_22_8_to_tile_23_8_3;
	wire vertical_tile_23_8_to_tile_22_8_0;
	wire vertical_tile_23_8_to_tile_22_8_1;
	wire vertical_tile_23_8_to_tile_22_8_2;
	wire vertical_tile_23_8_to_tile_22_8_3;

	wire vertical_tile_22_9_to_tile_23_9_0;
	wire vertical_tile_22_9_to_tile_23_9_1;
	wire vertical_tile_22_9_to_tile_23_9_2;
	wire vertical_tile_22_9_to_tile_23_9_3;
	wire vertical_tile_23_9_to_tile_22_9_0;
	wire vertical_tile_23_9_to_tile_22_9_1;
	wire vertical_tile_23_9_to_tile_22_9_2;
	wire vertical_tile_23_9_to_tile_22_9_3;

	wire vertical_tile_22_10_to_tile_23_10_0;
	wire vertical_tile_22_10_to_tile_23_10_1;
	wire vertical_tile_22_10_to_tile_23_10_2;
	wire vertical_tile_22_10_to_tile_23_10_3;
	wire vertical_tile_23_10_to_tile_22_10_0;
	wire vertical_tile_23_10_to_tile_22_10_1;
	wire vertical_tile_23_10_to_tile_22_10_2;
	wire vertical_tile_23_10_to_tile_22_10_3;

	wire vertical_tile_22_11_to_tile_23_11_0;
	wire vertical_tile_22_11_to_tile_23_11_1;
	wire vertical_tile_22_11_to_tile_23_11_2;
	wire vertical_tile_22_11_to_tile_23_11_3;
	wire vertical_tile_23_11_to_tile_22_11_0;
	wire vertical_tile_23_11_to_tile_22_11_1;
	wire vertical_tile_23_11_to_tile_22_11_2;
	wire vertical_tile_23_11_to_tile_22_11_3;

	wire vertical_tile_22_12_to_tile_23_12_0;
	wire vertical_tile_22_12_to_tile_23_12_1;
	wire vertical_tile_22_12_to_tile_23_12_2;
	wire vertical_tile_22_12_to_tile_23_12_3;
	wire vertical_tile_23_12_to_tile_22_12_0;
	wire vertical_tile_23_12_to_tile_22_12_1;
	wire vertical_tile_23_12_to_tile_22_12_2;
	wire vertical_tile_23_12_to_tile_22_12_3;

	wire vertical_tile_22_13_to_tile_23_13_0;
	wire vertical_tile_22_13_to_tile_23_13_1;
	wire vertical_tile_22_13_to_tile_23_13_2;
	wire vertical_tile_22_13_to_tile_23_13_3;
	wire vertical_tile_23_13_to_tile_22_13_0;
	wire vertical_tile_23_13_to_tile_22_13_1;
	wire vertical_tile_23_13_to_tile_22_13_2;
	wire vertical_tile_23_13_to_tile_22_13_3;

	wire vertical_tile_22_14_to_tile_23_14_0;
	wire vertical_tile_22_14_to_tile_23_14_1;
	wire vertical_tile_22_14_to_tile_23_14_2;
	wire vertical_tile_22_14_to_tile_23_14_3;
	wire vertical_tile_23_14_to_tile_22_14_0;
	wire vertical_tile_23_14_to_tile_22_14_1;
	wire vertical_tile_23_14_to_tile_22_14_2;
	wire vertical_tile_23_14_to_tile_22_14_3;

	wire vertical_tile_22_15_to_tile_23_15_0;
	wire vertical_tile_22_15_to_tile_23_15_1;
	wire vertical_tile_22_15_to_tile_23_15_2;
	wire vertical_tile_22_15_to_tile_23_15_3;
	wire vertical_tile_23_15_to_tile_22_15_0;
	wire vertical_tile_23_15_to_tile_22_15_1;
	wire vertical_tile_23_15_to_tile_22_15_2;
	wire vertical_tile_23_15_to_tile_22_15_3;

	wire vertical_tile_22_16_to_tile_23_16_0;
	wire vertical_tile_22_16_to_tile_23_16_1;
	wire vertical_tile_22_16_to_tile_23_16_2;
	wire vertical_tile_22_16_to_tile_23_16_3;
	wire vertical_tile_23_16_to_tile_22_16_0;
	wire vertical_tile_23_16_to_tile_22_16_1;
	wire vertical_tile_23_16_to_tile_22_16_2;
	wire vertical_tile_23_16_to_tile_22_16_3;

	wire vertical_tile_22_17_to_tile_23_17_0;
	wire vertical_tile_22_17_to_tile_23_17_1;
	wire vertical_tile_22_17_to_tile_23_17_2;
	wire vertical_tile_22_17_to_tile_23_17_3;
	wire vertical_tile_23_17_to_tile_22_17_0;
	wire vertical_tile_23_17_to_tile_22_17_1;
	wire vertical_tile_23_17_to_tile_22_17_2;
	wire vertical_tile_23_17_to_tile_22_17_3;

	wire vertical_tile_22_18_to_tile_23_18_0;
	wire vertical_tile_22_18_to_tile_23_18_1;
	wire vertical_tile_22_18_to_tile_23_18_2;
	wire vertical_tile_22_18_to_tile_23_18_3;
	wire vertical_tile_23_18_to_tile_22_18_0;
	wire vertical_tile_23_18_to_tile_22_18_1;
	wire vertical_tile_23_18_to_tile_22_18_2;
	wire vertical_tile_23_18_to_tile_22_18_3;

	wire vertical_tile_22_19_to_tile_23_19_0;
	wire vertical_tile_22_19_to_tile_23_19_1;
	wire vertical_tile_22_19_to_tile_23_19_2;
	wire vertical_tile_22_19_to_tile_23_19_3;
	wire vertical_tile_23_19_to_tile_22_19_0;
	wire vertical_tile_23_19_to_tile_22_19_1;
	wire vertical_tile_23_19_to_tile_22_19_2;
	wire vertical_tile_23_19_to_tile_22_19_3;

	wire vertical_tile_22_20_to_tile_23_20_0;
	wire vertical_tile_22_20_to_tile_23_20_1;
	wire vertical_tile_22_20_to_tile_23_20_2;
	wire vertical_tile_22_20_to_tile_23_20_3;
	wire vertical_tile_23_20_to_tile_22_20_0;
	wire vertical_tile_23_20_to_tile_22_20_1;
	wire vertical_tile_23_20_to_tile_22_20_2;
	wire vertical_tile_23_20_to_tile_22_20_3;

	wire vertical_tile_22_21_to_tile_23_21_0;
	wire vertical_tile_22_21_to_tile_23_21_1;
	wire vertical_tile_22_21_to_tile_23_21_2;
	wire vertical_tile_22_21_to_tile_23_21_3;
	wire vertical_tile_23_21_to_tile_22_21_0;
	wire vertical_tile_23_21_to_tile_22_21_1;
	wire vertical_tile_23_21_to_tile_22_21_2;
	wire vertical_tile_23_21_to_tile_22_21_3;

	wire vertical_tile_22_22_to_tile_23_22_0;
	wire vertical_tile_22_22_to_tile_23_22_1;
	wire vertical_tile_22_22_to_tile_23_22_2;
	wire vertical_tile_22_22_to_tile_23_22_3;
	wire vertical_tile_23_22_to_tile_22_22_0;
	wire vertical_tile_23_22_to_tile_22_22_1;
	wire vertical_tile_23_22_to_tile_22_22_2;
	wire vertical_tile_23_22_to_tile_22_22_3;

	wire vertical_tile_22_23_to_tile_23_23_0;
	wire vertical_tile_22_23_to_tile_23_23_1;
	wire vertical_tile_22_23_to_tile_23_23_2;
	wire vertical_tile_22_23_to_tile_23_23_3;
	wire vertical_tile_23_23_to_tile_22_23_0;
	wire vertical_tile_23_23_to_tile_22_23_1;
	wire vertical_tile_23_23_to_tile_22_23_2;
	wire vertical_tile_23_23_to_tile_22_23_3;

	wire vertical_tile_22_24_to_tile_23_24_0;
	wire vertical_tile_22_24_to_tile_23_24_1;
	wire vertical_tile_22_24_to_tile_23_24_2;
	wire vertical_tile_22_24_to_tile_23_24_3;
	wire vertical_tile_23_24_to_tile_22_24_0;
	wire vertical_tile_23_24_to_tile_22_24_1;
	wire vertical_tile_23_24_to_tile_22_24_2;
	wire vertical_tile_23_24_to_tile_22_24_3;

	wire vertical_tile_22_25_to_tile_23_25_0;
	wire vertical_tile_22_25_to_tile_23_25_1;
	wire vertical_tile_22_25_to_tile_23_25_2;
	wire vertical_tile_22_25_to_tile_23_25_3;
	wire vertical_tile_23_25_to_tile_22_25_0;
	wire vertical_tile_23_25_to_tile_22_25_1;
	wire vertical_tile_23_25_to_tile_22_25_2;
	wire vertical_tile_23_25_to_tile_22_25_3;

	wire vertical_tile_22_26_to_tile_23_26_0;
	wire vertical_tile_22_26_to_tile_23_26_1;
	wire vertical_tile_22_26_to_tile_23_26_2;
	wire vertical_tile_22_26_to_tile_23_26_3;
	wire vertical_tile_23_26_to_tile_22_26_0;
	wire vertical_tile_23_26_to_tile_22_26_1;
	wire vertical_tile_23_26_to_tile_22_26_2;
	wire vertical_tile_23_26_to_tile_22_26_3;

	wire vertical_tile_22_27_to_tile_23_27_0;
	wire vertical_tile_22_27_to_tile_23_27_1;
	wire vertical_tile_22_27_to_tile_23_27_2;
	wire vertical_tile_22_27_to_tile_23_27_3;
	wire vertical_tile_23_27_to_tile_22_27_0;
	wire vertical_tile_23_27_to_tile_22_27_1;
	wire vertical_tile_23_27_to_tile_22_27_2;
	wire vertical_tile_23_27_to_tile_22_27_3;

	wire vertical_tile_22_28_to_tile_23_28_0;
	wire vertical_tile_22_28_to_tile_23_28_1;
	wire vertical_tile_22_28_to_tile_23_28_2;
	wire vertical_tile_22_28_to_tile_23_28_3;
	wire vertical_tile_23_28_to_tile_22_28_0;
	wire vertical_tile_23_28_to_tile_22_28_1;
	wire vertical_tile_23_28_to_tile_22_28_2;
	wire vertical_tile_23_28_to_tile_22_28_3;

	wire vertical_tile_22_29_to_tile_23_29_0;
	wire vertical_tile_22_29_to_tile_23_29_1;
	wire vertical_tile_22_29_to_tile_23_29_2;
	wire vertical_tile_22_29_to_tile_23_29_3;
	wire vertical_tile_23_29_to_tile_22_29_0;
	wire vertical_tile_23_29_to_tile_22_29_1;
	wire vertical_tile_23_29_to_tile_22_29_2;
	wire vertical_tile_23_29_to_tile_22_29_3;

	wire vertical_tile_22_30_to_tile_23_30_0;
	wire vertical_tile_22_30_to_tile_23_30_1;
	wire vertical_tile_22_30_to_tile_23_30_2;
	wire vertical_tile_22_30_to_tile_23_30_3;
	wire vertical_tile_23_30_to_tile_22_30_0;
	wire vertical_tile_23_30_to_tile_22_30_1;
	wire vertical_tile_23_30_to_tile_22_30_2;
	wire vertical_tile_23_30_to_tile_22_30_3;

	wire vertical_tile_22_31_to_tile_23_31_0;
	wire vertical_tile_22_31_to_tile_23_31_1;
	wire vertical_tile_22_31_to_tile_23_31_2;
	wire vertical_tile_22_31_to_tile_23_31_3;
	wire vertical_tile_23_31_to_tile_22_31_0;
	wire vertical_tile_23_31_to_tile_22_31_1;
	wire vertical_tile_23_31_to_tile_22_31_2;
	wire vertical_tile_23_31_to_tile_22_31_3;

	wire vertical_tile_23_0_to_tile_24_0_0;
	wire vertical_tile_23_0_to_tile_24_0_1;
	wire vertical_tile_23_0_to_tile_24_0_2;
	wire vertical_tile_23_0_to_tile_24_0_3;
	wire vertical_tile_24_0_to_tile_23_0_0;
	wire vertical_tile_24_0_to_tile_23_0_1;
	wire vertical_tile_24_0_to_tile_23_0_2;
	wire vertical_tile_24_0_to_tile_23_0_3;

	wire vertical_tile_23_1_to_tile_24_1_0;
	wire vertical_tile_23_1_to_tile_24_1_1;
	wire vertical_tile_23_1_to_tile_24_1_2;
	wire vertical_tile_23_1_to_tile_24_1_3;
	wire vertical_tile_24_1_to_tile_23_1_0;
	wire vertical_tile_24_1_to_tile_23_1_1;
	wire vertical_tile_24_1_to_tile_23_1_2;
	wire vertical_tile_24_1_to_tile_23_1_3;

	wire vertical_tile_23_2_to_tile_24_2_0;
	wire vertical_tile_23_2_to_tile_24_2_1;
	wire vertical_tile_23_2_to_tile_24_2_2;
	wire vertical_tile_23_2_to_tile_24_2_3;
	wire vertical_tile_24_2_to_tile_23_2_0;
	wire vertical_tile_24_2_to_tile_23_2_1;
	wire vertical_tile_24_2_to_tile_23_2_2;
	wire vertical_tile_24_2_to_tile_23_2_3;

	wire vertical_tile_23_3_to_tile_24_3_0;
	wire vertical_tile_23_3_to_tile_24_3_1;
	wire vertical_tile_23_3_to_tile_24_3_2;
	wire vertical_tile_23_3_to_tile_24_3_3;
	wire vertical_tile_24_3_to_tile_23_3_0;
	wire vertical_tile_24_3_to_tile_23_3_1;
	wire vertical_tile_24_3_to_tile_23_3_2;
	wire vertical_tile_24_3_to_tile_23_3_3;

	wire vertical_tile_23_4_to_tile_24_4_0;
	wire vertical_tile_23_4_to_tile_24_4_1;
	wire vertical_tile_23_4_to_tile_24_4_2;
	wire vertical_tile_23_4_to_tile_24_4_3;
	wire vertical_tile_24_4_to_tile_23_4_0;
	wire vertical_tile_24_4_to_tile_23_4_1;
	wire vertical_tile_24_4_to_tile_23_4_2;
	wire vertical_tile_24_4_to_tile_23_4_3;

	wire vertical_tile_23_5_to_tile_24_5_0;
	wire vertical_tile_23_5_to_tile_24_5_1;
	wire vertical_tile_23_5_to_tile_24_5_2;
	wire vertical_tile_23_5_to_tile_24_5_3;
	wire vertical_tile_24_5_to_tile_23_5_0;
	wire vertical_tile_24_5_to_tile_23_5_1;
	wire vertical_tile_24_5_to_tile_23_5_2;
	wire vertical_tile_24_5_to_tile_23_5_3;

	wire vertical_tile_23_6_to_tile_24_6_0;
	wire vertical_tile_23_6_to_tile_24_6_1;
	wire vertical_tile_23_6_to_tile_24_6_2;
	wire vertical_tile_23_6_to_tile_24_6_3;
	wire vertical_tile_24_6_to_tile_23_6_0;
	wire vertical_tile_24_6_to_tile_23_6_1;
	wire vertical_tile_24_6_to_tile_23_6_2;
	wire vertical_tile_24_6_to_tile_23_6_3;

	wire vertical_tile_23_7_to_tile_24_7_0;
	wire vertical_tile_23_7_to_tile_24_7_1;
	wire vertical_tile_23_7_to_tile_24_7_2;
	wire vertical_tile_23_7_to_tile_24_7_3;
	wire vertical_tile_24_7_to_tile_23_7_0;
	wire vertical_tile_24_7_to_tile_23_7_1;
	wire vertical_tile_24_7_to_tile_23_7_2;
	wire vertical_tile_24_7_to_tile_23_7_3;

	wire vertical_tile_23_8_to_tile_24_8_0;
	wire vertical_tile_23_8_to_tile_24_8_1;
	wire vertical_tile_23_8_to_tile_24_8_2;
	wire vertical_tile_23_8_to_tile_24_8_3;
	wire vertical_tile_24_8_to_tile_23_8_0;
	wire vertical_tile_24_8_to_tile_23_8_1;
	wire vertical_tile_24_8_to_tile_23_8_2;
	wire vertical_tile_24_8_to_tile_23_8_3;

	wire vertical_tile_23_9_to_tile_24_9_0;
	wire vertical_tile_23_9_to_tile_24_9_1;
	wire vertical_tile_23_9_to_tile_24_9_2;
	wire vertical_tile_23_9_to_tile_24_9_3;
	wire vertical_tile_24_9_to_tile_23_9_0;
	wire vertical_tile_24_9_to_tile_23_9_1;
	wire vertical_tile_24_9_to_tile_23_9_2;
	wire vertical_tile_24_9_to_tile_23_9_3;

	wire vertical_tile_23_10_to_tile_24_10_0;
	wire vertical_tile_23_10_to_tile_24_10_1;
	wire vertical_tile_23_10_to_tile_24_10_2;
	wire vertical_tile_23_10_to_tile_24_10_3;
	wire vertical_tile_24_10_to_tile_23_10_0;
	wire vertical_tile_24_10_to_tile_23_10_1;
	wire vertical_tile_24_10_to_tile_23_10_2;
	wire vertical_tile_24_10_to_tile_23_10_3;

	wire vertical_tile_23_11_to_tile_24_11_0;
	wire vertical_tile_23_11_to_tile_24_11_1;
	wire vertical_tile_23_11_to_tile_24_11_2;
	wire vertical_tile_23_11_to_tile_24_11_3;
	wire vertical_tile_24_11_to_tile_23_11_0;
	wire vertical_tile_24_11_to_tile_23_11_1;
	wire vertical_tile_24_11_to_tile_23_11_2;
	wire vertical_tile_24_11_to_tile_23_11_3;

	wire vertical_tile_23_12_to_tile_24_12_0;
	wire vertical_tile_23_12_to_tile_24_12_1;
	wire vertical_tile_23_12_to_tile_24_12_2;
	wire vertical_tile_23_12_to_tile_24_12_3;
	wire vertical_tile_24_12_to_tile_23_12_0;
	wire vertical_tile_24_12_to_tile_23_12_1;
	wire vertical_tile_24_12_to_tile_23_12_2;
	wire vertical_tile_24_12_to_tile_23_12_3;

	wire vertical_tile_23_13_to_tile_24_13_0;
	wire vertical_tile_23_13_to_tile_24_13_1;
	wire vertical_tile_23_13_to_tile_24_13_2;
	wire vertical_tile_23_13_to_tile_24_13_3;
	wire vertical_tile_24_13_to_tile_23_13_0;
	wire vertical_tile_24_13_to_tile_23_13_1;
	wire vertical_tile_24_13_to_tile_23_13_2;
	wire vertical_tile_24_13_to_tile_23_13_3;

	wire vertical_tile_23_14_to_tile_24_14_0;
	wire vertical_tile_23_14_to_tile_24_14_1;
	wire vertical_tile_23_14_to_tile_24_14_2;
	wire vertical_tile_23_14_to_tile_24_14_3;
	wire vertical_tile_24_14_to_tile_23_14_0;
	wire vertical_tile_24_14_to_tile_23_14_1;
	wire vertical_tile_24_14_to_tile_23_14_2;
	wire vertical_tile_24_14_to_tile_23_14_3;

	wire vertical_tile_23_15_to_tile_24_15_0;
	wire vertical_tile_23_15_to_tile_24_15_1;
	wire vertical_tile_23_15_to_tile_24_15_2;
	wire vertical_tile_23_15_to_tile_24_15_3;
	wire vertical_tile_24_15_to_tile_23_15_0;
	wire vertical_tile_24_15_to_tile_23_15_1;
	wire vertical_tile_24_15_to_tile_23_15_2;
	wire vertical_tile_24_15_to_tile_23_15_3;

	wire vertical_tile_23_16_to_tile_24_16_0;
	wire vertical_tile_23_16_to_tile_24_16_1;
	wire vertical_tile_23_16_to_tile_24_16_2;
	wire vertical_tile_23_16_to_tile_24_16_3;
	wire vertical_tile_24_16_to_tile_23_16_0;
	wire vertical_tile_24_16_to_tile_23_16_1;
	wire vertical_tile_24_16_to_tile_23_16_2;
	wire vertical_tile_24_16_to_tile_23_16_3;

	wire vertical_tile_23_17_to_tile_24_17_0;
	wire vertical_tile_23_17_to_tile_24_17_1;
	wire vertical_tile_23_17_to_tile_24_17_2;
	wire vertical_tile_23_17_to_tile_24_17_3;
	wire vertical_tile_24_17_to_tile_23_17_0;
	wire vertical_tile_24_17_to_tile_23_17_1;
	wire vertical_tile_24_17_to_tile_23_17_2;
	wire vertical_tile_24_17_to_tile_23_17_3;

	wire vertical_tile_23_18_to_tile_24_18_0;
	wire vertical_tile_23_18_to_tile_24_18_1;
	wire vertical_tile_23_18_to_tile_24_18_2;
	wire vertical_tile_23_18_to_tile_24_18_3;
	wire vertical_tile_24_18_to_tile_23_18_0;
	wire vertical_tile_24_18_to_tile_23_18_1;
	wire vertical_tile_24_18_to_tile_23_18_2;
	wire vertical_tile_24_18_to_tile_23_18_3;

	wire vertical_tile_23_19_to_tile_24_19_0;
	wire vertical_tile_23_19_to_tile_24_19_1;
	wire vertical_tile_23_19_to_tile_24_19_2;
	wire vertical_tile_23_19_to_tile_24_19_3;
	wire vertical_tile_24_19_to_tile_23_19_0;
	wire vertical_tile_24_19_to_tile_23_19_1;
	wire vertical_tile_24_19_to_tile_23_19_2;
	wire vertical_tile_24_19_to_tile_23_19_3;

	wire vertical_tile_23_20_to_tile_24_20_0;
	wire vertical_tile_23_20_to_tile_24_20_1;
	wire vertical_tile_23_20_to_tile_24_20_2;
	wire vertical_tile_23_20_to_tile_24_20_3;
	wire vertical_tile_24_20_to_tile_23_20_0;
	wire vertical_tile_24_20_to_tile_23_20_1;
	wire vertical_tile_24_20_to_tile_23_20_2;
	wire vertical_tile_24_20_to_tile_23_20_3;

	wire vertical_tile_23_21_to_tile_24_21_0;
	wire vertical_tile_23_21_to_tile_24_21_1;
	wire vertical_tile_23_21_to_tile_24_21_2;
	wire vertical_tile_23_21_to_tile_24_21_3;
	wire vertical_tile_24_21_to_tile_23_21_0;
	wire vertical_tile_24_21_to_tile_23_21_1;
	wire vertical_tile_24_21_to_tile_23_21_2;
	wire vertical_tile_24_21_to_tile_23_21_3;

	wire vertical_tile_23_22_to_tile_24_22_0;
	wire vertical_tile_23_22_to_tile_24_22_1;
	wire vertical_tile_23_22_to_tile_24_22_2;
	wire vertical_tile_23_22_to_tile_24_22_3;
	wire vertical_tile_24_22_to_tile_23_22_0;
	wire vertical_tile_24_22_to_tile_23_22_1;
	wire vertical_tile_24_22_to_tile_23_22_2;
	wire vertical_tile_24_22_to_tile_23_22_3;

	wire vertical_tile_23_23_to_tile_24_23_0;
	wire vertical_tile_23_23_to_tile_24_23_1;
	wire vertical_tile_23_23_to_tile_24_23_2;
	wire vertical_tile_23_23_to_tile_24_23_3;
	wire vertical_tile_24_23_to_tile_23_23_0;
	wire vertical_tile_24_23_to_tile_23_23_1;
	wire vertical_tile_24_23_to_tile_23_23_2;
	wire vertical_tile_24_23_to_tile_23_23_3;

	wire vertical_tile_23_24_to_tile_24_24_0;
	wire vertical_tile_23_24_to_tile_24_24_1;
	wire vertical_tile_23_24_to_tile_24_24_2;
	wire vertical_tile_23_24_to_tile_24_24_3;
	wire vertical_tile_24_24_to_tile_23_24_0;
	wire vertical_tile_24_24_to_tile_23_24_1;
	wire vertical_tile_24_24_to_tile_23_24_2;
	wire vertical_tile_24_24_to_tile_23_24_3;

	wire vertical_tile_23_25_to_tile_24_25_0;
	wire vertical_tile_23_25_to_tile_24_25_1;
	wire vertical_tile_23_25_to_tile_24_25_2;
	wire vertical_tile_23_25_to_tile_24_25_3;
	wire vertical_tile_24_25_to_tile_23_25_0;
	wire vertical_tile_24_25_to_tile_23_25_1;
	wire vertical_tile_24_25_to_tile_23_25_2;
	wire vertical_tile_24_25_to_tile_23_25_3;

	wire vertical_tile_23_26_to_tile_24_26_0;
	wire vertical_tile_23_26_to_tile_24_26_1;
	wire vertical_tile_23_26_to_tile_24_26_2;
	wire vertical_tile_23_26_to_tile_24_26_3;
	wire vertical_tile_24_26_to_tile_23_26_0;
	wire vertical_tile_24_26_to_tile_23_26_1;
	wire vertical_tile_24_26_to_tile_23_26_2;
	wire vertical_tile_24_26_to_tile_23_26_3;

	wire vertical_tile_23_27_to_tile_24_27_0;
	wire vertical_tile_23_27_to_tile_24_27_1;
	wire vertical_tile_23_27_to_tile_24_27_2;
	wire vertical_tile_23_27_to_tile_24_27_3;
	wire vertical_tile_24_27_to_tile_23_27_0;
	wire vertical_tile_24_27_to_tile_23_27_1;
	wire vertical_tile_24_27_to_tile_23_27_2;
	wire vertical_tile_24_27_to_tile_23_27_3;

	wire vertical_tile_23_28_to_tile_24_28_0;
	wire vertical_tile_23_28_to_tile_24_28_1;
	wire vertical_tile_23_28_to_tile_24_28_2;
	wire vertical_tile_23_28_to_tile_24_28_3;
	wire vertical_tile_24_28_to_tile_23_28_0;
	wire vertical_tile_24_28_to_tile_23_28_1;
	wire vertical_tile_24_28_to_tile_23_28_2;
	wire vertical_tile_24_28_to_tile_23_28_3;

	wire vertical_tile_23_29_to_tile_24_29_0;
	wire vertical_tile_23_29_to_tile_24_29_1;
	wire vertical_tile_23_29_to_tile_24_29_2;
	wire vertical_tile_23_29_to_tile_24_29_3;
	wire vertical_tile_24_29_to_tile_23_29_0;
	wire vertical_tile_24_29_to_tile_23_29_1;
	wire vertical_tile_24_29_to_tile_23_29_2;
	wire vertical_tile_24_29_to_tile_23_29_3;

	wire vertical_tile_23_30_to_tile_24_30_0;
	wire vertical_tile_23_30_to_tile_24_30_1;
	wire vertical_tile_23_30_to_tile_24_30_2;
	wire vertical_tile_23_30_to_tile_24_30_3;
	wire vertical_tile_24_30_to_tile_23_30_0;
	wire vertical_tile_24_30_to_tile_23_30_1;
	wire vertical_tile_24_30_to_tile_23_30_2;
	wire vertical_tile_24_30_to_tile_23_30_3;

	wire vertical_tile_23_31_to_tile_24_31_0;
	wire vertical_tile_23_31_to_tile_24_31_1;
	wire vertical_tile_23_31_to_tile_24_31_2;
	wire vertical_tile_23_31_to_tile_24_31_3;
	wire vertical_tile_24_31_to_tile_23_31_0;
	wire vertical_tile_24_31_to_tile_23_31_1;
	wire vertical_tile_24_31_to_tile_23_31_2;
	wire vertical_tile_24_31_to_tile_23_31_3;

	wire vertical_tile_24_0_to_tile_25_0_0;
	wire vertical_tile_24_0_to_tile_25_0_1;
	wire vertical_tile_24_0_to_tile_25_0_2;
	wire vertical_tile_24_0_to_tile_25_0_3;
	wire vertical_tile_25_0_to_tile_24_0_0;
	wire vertical_tile_25_0_to_tile_24_0_1;
	wire vertical_tile_25_0_to_tile_24_0_2;
	wire vertical_tile_25_0_to_tile_24_0_3;

	wire vertical_tile_24_1_to_tile_25_1_0;
	wire vertical_tile_24_1_to_tile_25_1_1;
	wire vertical_tile_24_1_to_tile_25_1_2;
	wire vertical_tile_24_1_to_tile_25_1_3;
	wire vertical_tile_25_1_to_tile_24_1_0;
	wire vertical_tile_25_1_to_tile_24_1_1;
	wire vertical_tile_25_1_to_tile_24_1_2;
	wire vertical_tile_25_1_to_tile_24_1_3;

	wire vertical_tile_24_2_to_tile_25_2_0;
	wire vertical_tile_24_2_to_tile_25_2_1;
	wire vertical_tile_24_2_to_tile_25_2_2;
	wire vertical_tile_24_2_to_tile_25_2_3;
	wire vertical_tile_25_2_to_tile_24_2_0;
	wire vertical_tile_25_2_to_tile_24_2_1;
	wire vertical_tile_25_2_to_tile_24_2_2;
	wire vertical_tile_25_2_to_tile_24_2_3;

	wire vertical_tile_24_3_to_tile_25_3_0;
	wire vertical_tile_24_3_to_tile_25_3_1;
	wire vertical_tile_24_3_to_tile_25_3_2;
	wire vertical_tile_24_3_to_tile_25_3_3;
	wire vertical_tile_25_3_to_tile_24_3_0;
	wire vertical_tile_25_3_to_tile_24_3_1;
	wire vertical_tile_25_3_to_tile_24_3_2;
	wire vertical_tile_25_3_to_tile_24_3_3;

	wire vertical_tile_24_4_to_tile_25_4_0;
	wire vertical_tile_24_4_to_tile_25_4_1;
	wire vertical_tile_24_4_to_tile_25_4_2;
	wire vertical_tile_24_4_to_tile_25_4_3;
	wire vertical_tile_25_4_to_tile_24_4_0;
	wire vertical_tile_25_4_to_tile_24_4_1;
	wire vertical_tile_25_4_to_tile_24_4_2;
	wire vertical_tile_25_4_to_tile_24_4_3;

	wire vertical_tile_24_5_to_tile_25_5_0;
	wire vertical_tile_24_5_to_tile_25_5_1;
	wire vertical_tile_24_5_to_tile_25_5_2;
	wire vertical_tile_24_5_to_tile_25_5_3;
	wire vertical_tile_25_5_to_tile_24_5_0;
	wire vertical_tile_25_5_to_tile_24_5_1;
	wire vertical_tile_25_5_to_tile_24_5_2;
	wire vertical_tile_25_5_to_tile_24_5_3;

	wire vertical_tile_24_6_to_tile_25_6_0;
	wire vertical_tile_24_6_to_tile_25_6_1;
	wire vertical_tile_24_6_to_tile_25_6_2;
	wire vertical_tile_24_6_to_tile_25_6_3;
	wire vertical_tile_25_6_to_tile_24_6_0;
	wire vertical_tile_25_6_to_tile_24_6_1;
	wire vertical_tile_25_6_to_tile_24_6_2;
	wire vertical_tile_25_6_to_tile_24_6_3;

	wire vertical_tile_24_7_to_tile_25_7_0;
	wire vertical_tile_24_7_to_tile_25_7_1;
	wire vertical_tile_24_7_to_tile_25_7_2;
	wire vertical_tile_24_7_to_tile_25_7_3;
	wire vertical_tile_25_7_to_tile_24_7_0;
	wire vertical_tile_25_7_to_tile_24_7_1;
	wire vertical_tile_25_7_to_tile_24_7_2;
	wire vertical_tile_25_7_to_tile_24_7_3;

	wire vertical_tile_24_8_to_tile_25_8_0;
	wire vertical_tile_24_8_to_tile_25_8_1;
	wire vertical_tile_24_8_to_tile_25_8_2;
	wire vertical_tile_24_8_to_tile_25_8_3;
	wire vertical_tile_25_8_to_tile_24_8_0;
	wire vertical_tile_25_8_to_tile_24_8_1;
	wire vertical_tile_25_8_to_tile_24_8_2;
	wire vertical_tile_25_8_to_tile_24_8_3;

	wire vertical_tile_24_9_to_tile_25_9_0;
	wire vertical_tile_24_9_to_tile_25_9_1;
	wire vertical_tile_24_9_to_tile_25_9_2;
	wire vertical_tile_24_9_to_tile_25_9_3;
	wire vertical_tile_25_9_to_tile_24_9_0;
	wire vertical_tile_25_9_to_tile_24_9_1;
	wire vertical_tile_25_9_to_tile_24_9_2;
	wire vertical_tile_25_9_to_tile_24_9_3;

	wire vertical_tile_24_10_to_tile_25_10_0;
	wire vertical_tile_24_10_to_tile_25_10_1;
	wire vertical_tile_24_10_to_tile_25_10_2;
	wire vertical_tile_24_10_to_tile_25_10_3;
	wire vertical_tile_25_10_to_tile_24_10_0;
	wire vertical_tile_25_10_to_tile_24_10_1;
	wire vertical_tile_25_10_to_tile_24_10_2;
	wire vertical_tile_25_10_to_tile_24_10_3;

	wire vertical_tile_24_11_to_tile_25_11_0;
	wire vertical_tile_24_11_to_tile_25_11_1;
	wire vertical_tile_24_11_to_tile_25_11_2;
	wire vertical_tile_24_11_to_tile_25_11_3;
	wire vertical_tile_25_11_to_tile_24_11_0;
	wire vertical_tile_25_11_to_tile_24_11_1;
	wire vertical_tile_25_11_to_tile_24_11_2;
	wire vertical_tile_25_11_to_tile_24_11_3;

	wire vertical_tile_24_12_to_tile_25_12_0;
	wire vertical_tile_24_12_to_tile_25_12_1;
	wire vertical_tile_24_12_to_tile_25_12_2;
	wire vertical_tile_24_12_to_tile_25_12_3;
	wire vertical_tile_25_12_to_tile_24_12_0;
	wire vertical_tile_25_12_to_tile_24_12_1;
	wire vertical_tile_25_12_to_tile_24_12_2;
	wire vertical_tile_25_12_to_tile_24_12_3;

	wire vertical_tile_24_13_to_tile_25_13_0;
	wire vertical_tile_24_13_to_tile_25_13_1;
	wire vertical_tile_24_13_to_tile_25_13_2;
	wire vertical_tile_24_13_to_tile_25_13_3;
	wire vertical_tile_25_13_to_tile_24_13_0;
	wire vertical_tile_25_13_to_tile_24_13_1;
	wire vertical_tile_25_13_to_tile_24_13_2;
	wire vertical_tile_25_13_to_tile_24_13_3;

	wire vertical_tile_24_14_to_tile_25_14_0;
	wire vertical_tile_24_14_to_tile_25_14_1;
	wire vertical_tile_24_14_to_tile_25_14_2;
	wire vertical_tile_24_14_to_tile_25_14_3;
	wire vertical_tile_25_14_to_tile_24_14_0;
	wire vertical_tile_25_14_to_tile_24_14_1;
	wire vertical_tile_25_14_to_tile_24_14_2;
	wire vertical_tile_25_14_to_tile_24_14_3;

	wire vertical_tile_24_15_to_tile_25_15_0;
	wire vertical_tile_24_15_to_tile_25_15_1;
	wire vertical_tile_24_15_to_tile_25_15_2;
	wire vertical_tile_24_15_to_tile_25_15_3;
	wire vertical_tile_25_15_to_tile_24_15_0;
	wire vertical_tile_25_15_to_tile_24_15_1;
	wire vertical_tile_25_15_to_tile_24_15_2;
	wire vertical_tile_25_15_to_tile_24_15_3;

	wire vertical_tile_24_16_to_tile_25_16_0;
	wire vertical_tile_24_16_to_tile_25_16_1;
	wire vertical_tile_24_16_to_tile_25_16_2;
	wire vertical_tile_24_16_to_tile_25_16_3;
	wire vertical_tile_25_16_to_tile_24_16_0;
	wire vertical_tile_25_16_to_tile_24_16_1;
	wire vertical_tile_25_16_to_tile_24_16_2;
	wire vertical_tile_25_16_to_tile_24_16_3;

	wire vertical_tile_24_17_to_tile_25_17_0;
	wire vertical_tile_24_17_to_tile_25_17_1;
	wire vertical_tile_24_17_to_tile_25_17_2;
	wire vertical_tile_24_17_to_tile_25_17_3;
	wire vertical_tile_25_17_to_tile_24_17_0;
	wire vertical_tile_25_17_to_tile_24_17_1;
	wire vertical_tile_25_17_to_tile_24_17_2;
	wire vertical_tile_25_17_to_tile_24_17_3;

	wire vertical_tile_24_18_to_tile_25_18_0;
	wire vertical_tile_24_18_to_tile_25_18_1;
	wire vertical_tile_24_18_to_tile_25_18_2;
	wire vertical_tile_24_18_to_tile_25_18_3;
	wire vertical_tile_25_18_to_tile_24_18_0;
	wire vertical_tile_25_18_to_tile_24_18_1;
	wire vertical_tile_25_18_to_tile_24_18_2;
	wire vertical_tile_25_18_to_tile_24_18_3;

	wire vertical_tile_24_19_to_tile_25_19_0;
	wire vertical_tile_24_19_to_tile_25_19_1;
	wire vertical_tile_24_19_to_tile_25_19_2;
	wire vertical_tile_24_19_to_tile_25_19_3;
	wire vertical_tile_25_19_to_tile_24_19_0;
	wire vertical_tile_25_19_to_tile_24_19_1;
	wire vertical_tile_25_19_to_tile_24_19_2;
	wire vertical_tile_25_19_to_tile_24_19_3;

	wire vertical_tile_24_20_to_tile_25_20_0;
	wire vertical_tile_24_20_to_tile_25_20_1;
	wire vertical_tile_24_20_to_tile_25_20_2;
	wire vertical_tile_24_20_to_tile_25_20_3;
	wire vertical_tile_25_20_to_tile_24_20_0;
	wire vertical_tile_25_20_to_tile_24_20_1;
	wire vertical_tile_25_20_to_tile_24_20_2;
	wire vertical_tile_25_20_to_tile_24_20_3;

	wire vertical_tile_24_21_to_tile_25_21_0;
	wire vertical_tile_24_21_to_tile_25_21_1;
	wire vertical_tile_24_21_to_tile_25_21_2;
	wire vertical_tile_24_21_to_tile_25_21_3;
	wire vertical_tile_25_21_to_tile_24_21_0;
	wire vertical_tile_25_21_to_tile_24_21_1;
	wire vertical_tile_25_21_to_tile_24_21_2;
	wire vertical_tile_25_21_to_tile_24_21_3;

	wire vertical_tile_24_22_to_tile_25_22_0;
	wire vertical_tile_24_22_to_tile_25_22_1;
	wire vertical_tile_24_22_to_tile_25_22_2;
	wire vertical_tile_24_22_to_tile_25_22_3;
	wire vertical_tile_25_22_to_tile_24_22_0;
	wire vertical_tile_25_22_to_tile_24_22_1;
	wire vertical_tile_25_22_to_tile_24_22_2;
	wire vertical_tile_25_22_to_tile_24_22_3;

	wire vertical_tile_24_23_to_tile_25_23_0;
	wire vertical_tile_24_23_to_tile_25_23_1;
	wire vertical_tile_24_23_to_tile_25_23_2;
	wire vertical_tile_24_23_to_tile_25_23_3;
	wire vertical_tile_25_23_to_tile_24_23_0;
	wire vertical_tile_25_23_to_tile_24_23_1;
	wire vertical_tile_25_23_to_tile_24_23_2;
	wire vertical_tile_25_23_to_tile_24_23_3;

	wire vertical_tile_24_24_to_tile_25_24_0;
	wire vertical_tile_24_24_to_tile_25_24_1;
	wire vertical_tile_24_24_to_tile_25_24_2;
	wire vertical_tile_24_24_to_tile_25_24_3;
	wire vertical_tile_25_24_to_tile_24_24_0;
	wire vertical_tile_25_24_to_tile_24_24_1;
	wire vertical_tile_25_24_to_tile_24_24_2;
	wire vertical_tile_25_24_to_tile_24_24_3;

	wire vertical_tile_24_25_to_tile_25_25_0;
	wire vertical_tile_24_25_to_tile_25_25_1;
	wire vertical_tile_24_25_to_tile_25_25_2;
	wire vertical_tile_24_25_to_tile_25_25_3;
	wire vertical_tile_25_25_to_tile_24_25_0;
	wire vertical_tile_25_25_to_tile_24_25_1;
	wire vertical_tile_25_25_to_tile_24_25_2;
	wire vertical_tile_25_25_to_tile_24_25_3;

	wire vertical_tile_24_26_to_tile_25_26_0;
	wire vertical_tile_24_26_to_tile_25_26_1;
	wire vertical_tile_24_26_to_tile_25_26_2;
	wire vertical_tile_24_26_to_tile_25_26_3;
	wire vertical_tile_25_26_to_tile_24_26_0;
	wire vertical_tile_25_26_to_tile_24_26_1;
	wire vertical_tile_25_26_to_tile_24_26_2;
	wire vertical_tile_25_26_to_tile_24_26_3;

	wire vertical_tile_24_27_to_tile_25_27_0;
	wire vertical_tile_24_27_to_tile_25_27_1;
	wire vertical_tile_24_27_to_tile_25_27_2;
	wire vertical_tile_24_27_to_tile_25_27_3;
	wire vertical_tile_25_27_to_tile_24_27_0;
	wire vertical_tile_25_27_to_tile_24_27_1;
	wire vertical_tile_25_27_to_tile_24_27_2;
	wire vertical_tile_25_27_to_tile_24_27_3;

	wire vertical_tile_24_28_to_tile_25_28_0;
	wire vertical_tile_24_28_to_tile_25_28_1;
	wire vertical_tile_24_28_to_tile_25_28_2;
	wire vertical_tile_24_28_to_tile_25_28_3;
	wire vertical_tile_25_28_to_tile_24_28_0;
	wire vertical_tile_25_28_to_tile_24_28_1;
	wire vertical_tile_25_28_to_tile_24_28_2;
	wire vertical_tile_25_28_to_tile_24_28_3;

	wire vertical_tile_24_29_to_tile_25_29_0;
	wire vertical_tile_24_29_to_tile_25_29_1;
	wire vertical_tile_24_29_to_tile_25_29_2;
	wire vertical_tile_24_29_to_tile_25_29_3;
	wire vertical_tile_25_29_to_tile_24_29_0;
	wire vertical_tile_25_29_to_tile_24_29_1;
	wire vertical_tile_25_29_to_tile_24_29_2;
	wire vertical_tile_25_29_to_tile_24_29_3;

	wire vertical_tile_24_30_to_tile_25_30_0;
	wire vertical_tile_24_30_to_tile_25_30_1;
	wire vertical_tile_24_30_to_tile_25_30_2;
	wire vertical_tile_24_30_to_tile_25_30_3;
	wire vertical_tile_25_30_to_tile_24_30_0;
	wire vertical_tile_25_30_to_tile_24_30_1;
	wire vertical_tile_25_30_to_tile_24_30_2;
	wire vertical_tile_25_30_to_tile_24_30_3;

	wire vertical_tile_24_31_to_tile_25_31_0;
	wire vertical_tile_24_31_to_tile_25_31_1;
	wire vertical_tile_24_31_to_tile_25_31_2;
	wire vertical_tile_24_31_to_tile_25_31_3;
	wire vertical_tile_25_31_to_tile_24_31_0;
	wire vertical_tile_25_31_to_tile_24_31_1;
	wire vertical_tile_25_31_to_tile_24_31_2;
	wire vertical_tile_25_31_to_tile_24_31_3;

	wire vertical_tile_25_0_to_tile_26_0_0;
	wire vertical_tile_25_0_to_tile_26_0_1;
	wire vertical_tile_25_0_to_tile_26_0_2;
	wire vertical_tile_25_0_to_tile_26_0_3;
	wire vertical_tile_26_0_to_tile_25_0_0;
	wire vertical_tile_26_0_to_tile_25_0_1;
	wire vertical_tile_26_0_to_tile_25_0_2;
	wire vertical_tile_26_0_to_tile_25_0_3;

	wire vertical_tile_25_1_to_tile_26_1_0;
	wire vertical_tile_25_1_to_tile_26_1_1;
	wire vertical_tile_25_1_to_tile_26_1_2;
	wire vertical_tile_25_1_to_tile_26_1_3;
	wire vertical_tile_26_1_to_tile_25_1_0;
	wire vertical_tile_26_1_to_tile_25_1_1;
	wire vertical_tile_26_1_to_tile_25_1_2;
	wire vertical_tile_26_1_to_tile_25_1_3;

	wire vertical_tile_25_2_to_tile_26_2_0;
	wire vertical_tile_25_2_to_tile_26_2_1;
	wire vertical_tile_25_2_to_tile_26_2_2;
	wire vertical_tile_25_2_to_tile_26_2_3;
	wire vertical_tile_26_2_to_tile_25_2_0;
	wire vertical_tile_26_2_to_tile_25_2_1;
	wire vertical_tile_26_2_to_tile_25_2_2;
	wire vertical_tile_26_2_to_tile_25_2_3;

	wire vertical_tile_25_3_to_tile_26_3_0;
	wire vertical_tile_25_3_to_tile_26_3_1;
	wire vertical_tile_25_3_to_tile_26_3_2;
	wire vertical_tile_25_3_to_tile_26_3_3;
	wire vertical_tile_26_3_to_tile_25_3_0;
	wire vertical_tile_26_3_to_tile_25_3_1;
	wire vertical_tile_26_3_to_tile_25_3_2;
	wire vertical_tile_26_3_to_tile_25_3_3;

	wire vertical_tile_25_4_to_tile_26_4_0;
	wire vertical_tile_25_4_to_tile_26_4_1;
	wire vertical_tile_25_4_to_tile_26_4_2;
	wire vertical_tile_25_4_to_tile_26_4_3;
	wire vertical_tile_26_4_to_tile_25_4_0;
	wire vertical_tile_26_4_to_tile_25_4_1;
	wire vertical_tile_26_4_to_tile_25_4_2;
	wire vertical_tile_26_4_to_tile_25_4_3;

	wire vertical_tile_25_5_to_tile_26_5_0;
	wire vertical_tile_25_5_to_tile_26_5_1;
	wire vertical_tile_25_5_to_tile_26_5_2;
	wire vertical_tile_25_5_to_tile_26_5_3;
	wire vertical_tile_26_5_to_tile_25_5_0;
	wire vertical_tile_26_5_to_tile_25_5_1;
	wire vertical_tile_26_5_to_tile_25_5_2;
	wire vertical_tile_26_5_to_tile_25_5_3;

	wire vertical_tile_25_6_to_tile_26_6_0;
	wire vertical_tile_25_6_to_tile_26_6_1;
	wire vertical_tile_25_6_to_tile_26_6_2;
	wire vertical_tile_25_6_to_tile_26_6_3;
	wire vertical_tile_26_6_to_tile_25_6_0;
	wire vertical_tile_26_6_to_tile_25_6_1;
	wire vertical_tile_26_6_to_tile_25_6_2;
	wire vertical_tile_26_6_to_tile_25_6_3;

	wire vertical_tile_25_7_to_tile_26_7_0;
	wire vertical_tile_25_7_to_tile_26_7_1;
	wire vertical_tile_25_7_to_tile_26_7_2;
	wire vertical_tile_25_7_to_tile_26_7_3;
	wire vertical_tile_26_7_to_tile_25_7_0;
	wire vertical_tile_26_7_to_tile_25_7_1;
	wire vertical_tile_26_7_to_tile_25_7_2;
	wire vertical_tile_26_7_to_tile_25_7_3;

	wire vertical_tile_25_8_to_tile_26_8_0;
	wire vertical_tile_25_8_to_tile_26_8_1;
	wire vertical_tile_25_8_to_tile_26_8_2;
	wire vertical_tile_25_8_to_tile_26_8_3;
	wire vertical_tile_26_8_to_tile_25_8_0;
	wire vertical_tile_26_8_to_tile_25_8_1;
	wire vertical_tile_26_8_to_tile_25_8_2;
	wire vertical_tile_26_8_to_tile_25_8_3;

	wire vertical_tile_25_9_to_tile_26_9_0;
	wire vertical_tile_25_9_to_tile_26_9_1;
	wire vertical_tile_25_9_to_tile_26_9_2;
	wire vertical_tile_25_9_to_tile_26_9_3;
	wire vertical_tile_26_9_to_tile_25_9_0;
	wire vertical_tile_26_9_to_tile_25_9_1;
	wire vertical_tile_26_9_to_tile_25_9_2;
	wire vertical_tile_26_9_to_tile_25_9_3;

	wire vertical_tile_25_10_to_tile_26_10_0;
	wire vertical_tile_25_10_to_tile_26_10_1;
	wire vertical_tile_25_10_to_tile_26_10_2;
	wire vertical_tile_25_10_to_tile_26_10_3;
	wire vertical_tile_26_10_to_tile_25_10_0;
	wire vertical_tile_26_10_to_tile_25_10_1;
	wire vertical_tile_26_10_to_tile_25_10_2;
	wire vertical_tile_26_10_to_tile_25_10_3;

	wire vertical_tile_25_11_to_tile_26_11_0;
	wire vertical_tile_25_11_to_tile_26_11_1;
	wire vertical_tile_25_11_to_tile_26_11_2;
	wire vertical_tile_25_11_to_tile_26_11_3;
	wire vertical_tile_26_11_to_tile_25_11_0;
	wire vertical_tile_26_11_to_tile_25_11_1;
	wire vertical_tile_26_11_to_tile_25_11_2;
	wire vertical_tile_26_11_to_tile_25_11_3;

	wire vertical_tile_25_12_to_tile_26_12_0;
	wire vertical_tile_25_12_to_tile_26_12_1;
	wire vertical_tile_25_12_to_tile_26_12_2;
	wire vertical_tile_25_12_to_tile_26_12_3;
	wire vertical_tile_26_12_to_tile_25_12_0;
	wire vertical_tile_26_12_to_tile_25_12_1;
	wire vertical_tile_26_12_to_tile_25_12_2;
	wire vertical_tile_26_12_to_tile_25_12_3;

	wire vertical_tile_25_13_to_tile_26_13_0;
	wire vertical_tile_25_13_to_tile_26_13_1;
	wire vertical_tile_25_13_to_tile_26_13_2;
	wire vertical_tile_25_13_to_tile_26_13_3;
	wire vertical_tile_26_13_to_tile_25_13_0;
	wire vertical_tile_26_13_to_tile_25_13_1;
	wire vertical_tile_26_13_to_tile_25_13_2;
	wire vertical_tile_26_13_to_tile_25_13_3;

	wire vertical_tile_25_14_to_tile_26_14_0;
	wire vertical_tile_25_14_to_tile_26_14_1;
	wire vertical_tile_25_14_to_tile_26_14_2;
	wire vertical_tile_25_14_to_tile_26_14_3;
	wire vertical_tile_26_14_to_tile_25_14_0;
	wire vertical_tile_26_14_to_tile_25_14_1;
	wire vertical_tile_26_14_to_tile_25_14_2;
	wire vertical_tile_26_14_to_tile_25_14_3;

	wire vertical_tile_25_15_to_tile_26_15_0;
	wire vertical_tile_25_15_to_tile_26_15_1;
	wire vertical_tile_25_15_to_tile_26_15_2;
	wire vertical_tile_25_15_to_tile_26_15_3;
	wire vertical_tile_26_15_to_tile_25_15_0;
	wire vertical_tile_26_15_to_tile_25_15_1;
	wire vertical_tile_26_15_to_tile_25_15_2;
	wire vertical_tile_26_15_to_tile_25_15_3;

	wire vertical_tile_25_16_to_tile_26_16_0;
	wire vertical_tile_25_16_to_tile_26_16_1;
	wire vertical_tile_25_16_to_tile_26_16_2;
	wire vertical_tile_25_16_to_tile_26_16_3;
	wire vertical_tile_26_16_to_tile_25_16_0;
	wire vertical_tile_26_16_to_tile_25_16_1;
	wire vertical_tile_26_16_to_tile_25_16_2;
	wire vertical_tile_26_16_to_tile_25_16_3;

	wire vertical_tile_25_17_to_tile_26_17_0;
	wire vertical_tile_25_17_to_tile_26_17_1;
	wire vertical_tile_25_17_to_tile_26_17_2;
	wire vertical_tile_25_17_to_tile_26_17_3;
	wire vertical_tile_26_17_to_tile_25_17_0;
	wire vertical_tile_26_17_to_tile_25_17_1;
	wire vertical_tile_26_17_to_tile_25_17_2;
	wire vertical_tile_26_17_to_tile_25_17_3;

	wire vertical_tile_25_18_to_tile_26_18_0;
	wire vertical_tile_25_18_to_tile_26_18_1;
	wire vertical_tile_25_18_to_tile_26_18_2;
	wire vertical_tile_25_18_to_tile_26_18_3;
	wire vertical_tile_26_18_to_tile_25_18_0;
	wire vertical_tile_26_18_to_tile_25_18_1;
	wire vertical_tile_26_18_to_tile_25_18_2;
	wire vertical_tile_26_18_to_tile_25_18_3;

	wire vertical_tile_25_19_to_tile_26_19_0;
	wire vertical_tile_25_19_to_tile_26_19_1;
	wire vertical_tile_25_19_to_tile_26_19_2;
	wire vertical_tile_25_19_to_tile_26_19_3;
	wire vertical_tile_26_19_to_tile_25_19_0;
	wire vertical_tile_26_19_to_tile_25_19_1;
	wire vertical_tile_26_19_to_tile_25_19_2;
	wire vertical_tile_26_19_to_tile_25_19_3;

	wire vertical_tile_25_20_to_tile_26_20_0;
	wire vertical_tile_25_20_to_tile_26_20_1;
	wire vertical_tile_25_20_to_tile_26_20_2;
	wire vertical_tile_25_20_to_tile_26_20_3;
	wire vertical_tile_26_20_to_tile_25_20_0;
	wire vertical_tile_26_20_to_tile_25_20_1;
	wire vertical_tile_26_20_to_tile_25_20_2;
	wire vertical_tile_26_20_to_tile_25_20_3;

	wire vertical_tile_25_21_to_tile_26_21_0;
	wire vertical_tile_25_21_to_tile_26_21_1;
	wire vertical_tile_25_21_to_tile_26_21_2;
	wire vertical_tile_25_21_to_tile_26_21_3;
	wire vertical_tile_26_21_to_tile_25_21_0;
	wire vertical_tile_26_21_to_tile_25_21_1;
	wire vertical_tile_26_21_to_tile_25_21_2;
	wire vertical_tile_26_21_to_tile_25_21_3;

	wire vertical_tile_25_22_to_tile_26_22_0;
	wire vertical_tile_25_22_to_tile_26_22_1;
	wire vertical_tile_25_22_to_tile_26_22_2;
	wire vertical_tile_25_22_to_tile_26_22_3;
	wire vertical_tile_26_22_to_tile_25_22_0;
	wire vertical_tile_26_22_to_tile_25_22_1;
	wire vertical_tile_26_22_to_tile_25_22_2;
	wire vertical_tile_26_22_to_tile_25_22_3;

	wire vertical_tile_25_23_to_tile_26_23_0;
	wire vertical_tile_25_23_to_tile_26_23_1;
	wire vertical_tile_25_23_to_tile_26_23_2;
	wire vertical_tile_25_23_to_tile_26_23_3;
	wire vertical_tile_26_23_to_tile_25_23_0;
	wire vertical_tile_26_23_to_tile_25_23_1;
	wire vertical_tile_26_23_to_tile_25_23_2;
	wire vertical_tile_26_23_to_tile_25_23_3;

	wire vertical_tile_25_24_to_tile_26_24_0;
	wire vertical_tile_25_24_to_tile_26_24_1;
	wire vertical_tile_25_24_to_tile_26_24_2;
	wire vertical_tile_25_24_to_tile_26_24_3;
	wire vertical_tile_26_24_to_tile_25_24_0;
	wire vertical_tile_26_24_to_tile_25_24_1;
	wire vertical_tile_26_24_to_tile_25_24_2;
	wire vertical_tile_26_24_to_tile_25_24_3;

	wire vertical_tile_25_25_to_tile_26_25_0;
	wire vertical_tile_25_25_to_tile_26_25_1;
	wire vertical_tile_25_25_to_tile_26_25_2;
	wire vertical_tile_25_25_to_tile_26_25_3;
	wire vertical_tile_26_25_to_tile_25_25_0;
	wire vertical_tile_26_25_to_tile_25_25_1;
	wire vertical_tile_26_25_to_tile_25_25_2;
	wire vertical_tile_26_25_to_tile_25_25_3;

	wire vertical_tile_25_26_to_tile_26_26_0;
	wire vertical_tile_25_26_to_tile_26_26_1;
	wire vertical_tile_25_26_to_tile_26_26_2;
	wire vertical_tile_25_26_to_tile_26_26_3;
	wire vertical_tile_26_26_to_tile_25_26_0;
	wire vertical_tile_26_26_to_tile_25_26_1;
	wire vertical_tile_26_26_to_tile_25_26_2;
	wire vertical_tile_26_26_to_tile_25_26_3;

	wire vertical_tile_25_27_to_tile_26_27_0;
	wire vertical_tile_25_27_to_tile_26_27_1;
	wire vertical_tile_25_27_to_tile_26_27_2;
	wire vertical_tile_25_27_to_tile_26_27_3;
	wire vertical_tile_26_27_to_tile_25_27_0;
	wire vertical_tile_26_27_to_tile_25_27_1;
	wire vertical_tile_26_27_to_tile_25_27_2;
	wire vertical_tile_26_27_to_tile_25_27_3;

	wire vertical_tile_25_28_to_tile_26_28_0;
	wire vertical_tile_25_28_to_tile_26_28_1;
	wire vertical_tile_25_28_to_tile_26_28_2;
	wire vertical_tile_25_28_to_tile_26_28_3;
	wire vertical_tile_26_28_to_tile_25_28_0;
	wire vertical_tile_26_28_to_tile_25_28_1;
	wire vertical_tile_26_28_to_tile_25_28_2;
	wire vertical_tile_26_28_to_tile_25_28_3;

	wire vertical_tile_25_29_to_tile_26_29_0;
	wire vertical_tile_25_29_to_tile_26_29_1;
	wire vertical_tile_25_29_to_tile_26_29_2;
	wire vertical_tile_25_29_to_tile_26_29_3;
	wire vertical_tile_26_29_to_tile_25_29_0;
	wire vertical_tile_26_29_to_tile_25_29_1;
	wire vertical_tile_26_29_to_tile_25_29_2;
	wire vertical_tile_26_29_to_tile_25_29_3;

	wire vertical_tile_25_30_to_tile_26_30_0;
	wire vertical_tile_25_30_to_tile_26_30_1;
	wire vertical_tile_25_30_to_tile_26_30_2;
	wire vertical_tile_25_30_to_tile_26_30_3;
	wire vertical_tile_26_30_to_tile_25_30_0;
	wire vertical_tile_26_30_to_tile_25_30_1;
	wire vertical_tile_26_30_to_tile_25_30_2;
	wire vertical_tile_26_30_to_tile_25_30_3;

	wire vertical_tile_25_31_to_tile_26_31_0;
	wire vertical_tile_25_31_to_tile_26_31_1;
	wire vertical_tile_25_31_to_tile_26_31_2;
	wire vertical_tile_25_31_to_tile_26_31_3;
	wire vertical_tile_26_31_to_tile_25_31_0;
	wire vertical_tile_26_31_to_tile_25_31_1;
	wire vertical_tile_26_31_to_tile_25_31_2;
	wire vertical_tile_26_31_to_tile_25_31_3;

	wire vertical_tile_26_0_to_tile_27_0_0;
	wire vertical_tile_26_0_to_tile_27_0_1;
	wire vertical_tile_26_0_to_tile_27_0_2;
	wire vertical_tile_26_0_to_tile_27_0_3;
	wire vertical_tile_27_0_to_tile_26_0_0;
	wire vertical_tile_27_0_to_tile_26_0_1;
	wire vertical_tile_27_0_to_tile_26_0_2;
	wire vertical_tile_27_0_to_tile_26_0_3;

	wire vertical_tile_26_1_to_tile_27_1_0;
	wire vertical_tile_26_1_to_tile_27_1_1;
	wire vertical_tile_26_1_to_tile_27_1_2;
	wire vertical_tile_26_1_to_tile_27_1_3;
	wire vertical_tile_27_1_to_tile_26_1_0;
	wire vertical_tile_27_1_to_tile_26_1_1;
	wire vertical_tile_27_1_to_tile_26_1_2;
	wire vertical_tile_27_1_to_tile_26_1_3;

	wire vertical_tile_26_2_to_tile_27_2_0;
	wire vertical_tile_26_2_to_tile_27_2_1;
	wire vertical_tile_26_2_to_tile_27_2_2;
	wire vertical_tile_26_2_to_tile_27_2_3;
	wire vertical_tile_27_2_to_tile_26_2_0;
	wire vertical_tile_27_2_to_tile_26_2_1;
	wire vertical_tile_27_2_to_tile_26_2_2;
	wire vertical_tile_27_2_to_tile_26_2_3;

	wire vertical_tile_26_3_to_tile_27_3_0;
	wire vertical_tile_26_3_to_tile_27_3_1;
	wire vertical_tile_26_3_to_tile_27_3_2;
	wire vertical_tile_26_3_to_tile_27_3_3;
	wire vertical_tile_27_3_to_tile_26_3_0;
	wire vertical_tile_27_3_to_tile_26_3_1;
	wire vertical_tile_27_3_to_tile_26_3_2;
	wire vertical_tile_27_3_to_tile_26_3_3;

	wire vertical_tile_26_4_to_tile_27_4_0;
	wire vertical_tile_26_4_to_tile_27_4_1;
	wire vertical_tile_26_4_to_tile_27_4_2;
	wire vertical_tile_26_4_to_tile_27_4_3;
	wire vertical_tile_27_4_to_tile_26_4_0;
	wire vertical_tile_27_4_to_tile_26_4_1;
	wire vertical_tile_27_4_to_tile_26_4_2;
	wire vertical_tile_27_4_to_tile_26_4_3;

	wire vertical_tile_26_5_to_tile_27_5_0;
	wire vertical_tile_26_5_to_tile_27_5_1;
	wire vertical_tile_26_5_to_tile_27_5_2;
	wire vertical_tile_26_5_to_tile_27_5_3;
	wire vertical_tile_27_5_to_tile_26_5_0;
	wire vertical_tile_27_5_to_tile_26_5_1;
	wire vertical_tile_27_5_to_tile_26_5_2;
	wire vertical_tile_27_5_to_tile_26_5_3;

	wire vertical_tile_26_6_to_tile_27_6_0;
	wire vertical_tile_26_6_to_tile_27_6_1;
	wire vertical_tile_26_6_to_tile_27_6_2;
	wire vertical_tile_26_6_to_tile_27_6_3;
	wire vertical_tile_27_6_to_tile_26_6_0;
	wire vertical_tile_27_6_to_tile_26_6_1;
	wire vertical_tile_27_6_to_tile_26_6_2;
	wire vertical_tile_27_6_to_tile_26_6_3;

	wire vertical_tile_26_7_to_tile_27_7_0;
	wire vertical_tile_26_7_to_tile_27_7_1;
	wire vertical_tile_26_7_to_tile_27_7_2;
	wire vertical_tile_26_7_to_tile_27_7_3;
	wire vertical_tile_27_7_to_tile_26_7_0;
	wire vertical_tile_27_7_to_tile_26_7_1;
	wire vertical_tile_27_7_to_tile_26_7_2;
	wire vertical_tile_27_7_to_tile_26_7_3;

	wire vertical_tile_26_8_to_tile_27_8_0;
	wire vertical_tile_26_8_to_tile_27_8_1;
	wire vertical_tile_26_8_to_tile_27_8_2;
	wire vertical_tile_26_8_to_tile_27_8_3;
	wire vertical_tile_27_8_to_tile_26_8_0;
	wire vertical_tile_27_8_to_tile_26_8_1;
	wire vertical_tile_27_8_to_tile_26_8_2;
	wire vertical_tile_27_8_to_tile_26_8_3;

	wire vertical_tile_26_9_to_tile_27_9_0;
	wire vertical_tile_26_9_to_tile_27_9_1;
	wire vertical_tile_26_9_to_tile_27_9_2;
	wire vertical_tile_26_9_to_tile_27_9_3;
	wire vertical_tile_27_9_to_tile_26_9_0;
	wire vertical_tile_27_9_to_tile_26_9_1;
	wire vertical_tile_27_9_to_tile_26_9_2;
	wire vertical_tile_27_9_to_tile_26_9_3;

	wire vertical_tile_26_10_to_tile_27_10_0;
	wire vertical_tile_26_10_to_tile_27_10_1;
	wire vertical_tile_26_10_to_tile_27_10_2;
	wire vertical_tile_26_10_to_tile_27_10_3;
	wire vertical_tile_27_10_to_tile_26_10_0;
	wire vertical_tile_27_10_to_tile_26_10_1;
	wire vertical_tile_27_10_to_tile_26_10_2;
	wire vertical_tile_27_10_to_tile_26_10_3;

	wire vertical_tile_26_11_to_tile_27_11_0;
	wire vertical_tile_26_11_to_tile_27_11_1;
	wire vertical_tile_26_11_to_tile_27_11_2;
	wire vertical_tile_26_11_to_tile_27_11_3;
	wire vertical_tile_27_11_to_tile_26_11_0;
	wire vertical_tile_27_11_to_tile_26_11_1;
	wire vertical_tile_27_11_to_tile_26_11_2;
	wire vertical_tile_27_11_to_tile_26_11_3;

	wire vertical_tile_26_12_to_tile_27_12_0;
	wire vertical_tile_26_12_to_tile_27_12_1;
	wire vertical_tile_26_12_to_tile_27_12_2;
	wire vertical_tile_26_12_to_tile_27_12_3;
	wire vertical_tile_27_12_to_tile_26_12_0;
	wire vertical_tile_27_12_to_tile_26_12_1;
	wire vertical_tile_27_12_to_tile_26_12_2;
	wire vertical_tile_27_12_to_tile_26_12_3;

	wire vertical_tile_26_13_to_tile_27_13_0;
	wire vertical_tile_26_13_to_tile_27_13_1;
	wire vertical_tile_26_13_to_tile_27_13_2;
	wire vertical_tile_26_13_to_tile_27_13_3;
	wire vertical_tile_27_13_to_tile_26_13_0;
	wire vertical_tile_27_13_to_tile_26_13_1;
	wire vertical_tile_27_13_to_tile_26_13_2;
	wire vertical_tile_27_13_to_tile_26_13_3;

	wire vertical_tile_26_14_to_tile_27_14_0;
	wire vertical_tile_26_14_to_tile_27_14_1;
	wire vertical_tile_26_14_to_tile_27_14_2;
	wire vertical_tile_26_14_to_tile_27_14_3;
	wire vertical_tile_27_14_to_tile_26_14_0;
	wire vertical_tile_27_14_to_tile_26_14_1;
	wire vertical_tile_27_14_to_tile_26_14_2;
	wire vertical_tile_27_14_to_tile_26_14_3;

	wire vertical_tile_26_15_to_tile_27_15_0;
	wire vertical_tile_26_15_to_tile_27_15_1;
	wire vertical_tile_26_15_to_tile_27_15_2;
	wire vertical_tile_26_15_to_tile_27_15_3;
	wire vertical_tile_27_15_to_tile_26_15_0;
	wire vertical_tile_27_15_to_tile_26_15_1;
	wire vertical_tile_27_15_to_tile_26_15_2;
	wire vertical_tile_27_15_to_tile_26_15_3;

	wire vertical_tile_26_16_to_tile_27_16_0;
	wire vertical_tile_26_16_to_tile_27_16_1;
	wire vertical_tile_26_16_to_tile_27_16_2;
	wire vertical_tile_26_16_to_tile_27_16_3;
	wire vertical_tile_27_16_to_tile_26_16_0;
	wire vertical_tile_27_16_to_tile_26_16_1;
	wire vertical_tile_27_16_to_tile_26_16_2;
	wire vertical_tile_27_16_to_tile_26_16_3;

	wire vertical_tile_26_17_to_tile_27_17_0;
	wire vertical_tile_26_17_to_tile_27_17_1;
	wire vertical_tile_26_17_to_tile_27_17_2;
	wire vertical_tile_26_17_to_tile_27_17_3;
	wire vertical_tile_27_17_to_tile_26_17_0;
	wire vertical_tile_27_17_to_tile_26_17_1;
	wire vertical_tile_27_17_to_tile_26_17_2;
	wire vertical_tile_27_17_to_tile_26_17_3;

	wire vertical_tile_26_18_to_tile_27_18_0;
	wire vertical_tile_26_18_to_tile_27_18_1;
	wire vertical_tile_26_18_to_tile_27_18_2;
	wire vertical_tile_26_18_to_tile_27_18_3;
	wire vertical_tile_27_18_to_tile_26_18_0;
	wire vertical_tile_27_18_to_tile_26_18_1;
	wire vertical_tile_27_18_to_tile_26_18_2;
	wire vertical_tile_27_18_to_tile_26_18_3;

	wire vertical_tile_26_19_to_tile_27_19_0;
	wire vertical_tile_26_19_to_tile_27_19_1;
	wire vertical_tile_26_19_to_tile_27_19_2;
	wire vertical_tile_26_19_to_tile_27_19_3;
	wire vertical_tile_27_19_to_tile_26_19_0;
	wire vertical_tile_27_19_to_tile_26_19_1;
	wire vertical_tile_27_19_to_tile_26_19_2;
	wire vertical_tile_27_19_to_tile_26_19_3;

	wire vertical_tile_26_20_to_tile_27_20_0;
	wire vertical_tile_26_20_to_tile_27_20_1;
	wire vertical_tile_26_20_to_tile_27_20_2;
	wire vertical_tile_26_20_to_tile_27_20_3;
	wire vertical_tile_27_20_to_tile_26_20_0;
	wire vertical_tile_27_20_to_tile_26_20_1;
	wire vertical_tile_27_20_to_tile_26_20_2;
	wire vertical_tile_27_20_to_tile_26_20_3;

	wire vertical_tile_26_21_to_tile_27_21_0;
	wire vertical_tile_26_21_to_tile_27_21_1;
	wire vertical_tile_26_21_to_tile_27_21_2;
	wire vertical_tile_26_21_to_tile_27_21_3;
	wire vertical_tile_27_21_to_tile_26_21_0;
	wire vertical_tile_27_21_to_tile_26_21_1;
	wire vertical_tile_27_21_to_tile_26_21_2;
	wire vertical_tile_27_21_to_tile_26_21_3;

	wire vertical_tile_26_22_to_tile_27_22_0;
	wire vertical_tile_26_22_to_tile_27_22_1;
	wire vertical_tile_26_22_to_tile_27_22_2;
	wire vertical_tile_26_22_to_tile_27_22_3;
	wire vertical_tile_27_22_to_tile_26_22_0;
	wire vertical_tile_27_22_to_tile_26_22_1;
	wire vertical_tile_27_22_to_tile_26_22_2;
	wire vertical_tile_27_22_to_tile_26_22_3;

	wire vertical_tile_26_23_to_tile_27_23_0;
	wire vertical_tile_26_23_to_tile_27_23_1;
	wire vertical_tile_26_23_to_tile_27_23_2;
	wire vertical_tile_26_23_to_tile_27_23_3;
	wire vertical_tile_27_23_to_tile_26_23_0;
	wire vertical_tile_27_23_to_tile_26_23_1;
	wire vertical_tile_27_23_to_tile_26_23_2;
	wire vertical_tile_27_23_to_tile_26_23_3;

	wire vertical_tile_26_24_to_tile_27_24_0;
	wire vertical_tile_26_24_to_tile_27_24_1;
	wire vertical_tile_26_24_to_tile_27_24_2;
	wire vertical_tile_26_24_to_tile_27_24_3;
	wire vertical_tile_27_24_to_tile_26_24_0;
	wire vertical_tile_27_24_to_tile_26_24_1;
	wire vertical_tile_27_24_to_tile_26_24_2;
	wire vertical_tile_27_24_to_tile_26_24_3;

	wire vertical_tile_26_25_to_tile_27_25_0;
	wire vertical_tile_26_25_to_tile_27_25_1;
	wire vertical_tile_26_25_to_tile_27_25_2;
	wire vertical_tile_26_25_to_tile_27_25_3;
	wire vertical_tile_27_25_to_tile_26_25_0;
	wire vertical_tile_27_25_to_tile_26_25_1;
	wire vertical_tile_27_25_to_tile_26_25_2;
	wire vertical_tile_27_25_to_tile_26_25_3;

	wire vertical_tile_26_26_to_tile_27_26_0;
	wire vertical_tile_26_26_to_tile_27_26_1;
	wire vertical_tile_26_26_to_tile_27_26_2;
	wire vertical_tile_26_26_to_tile_27_26_3;
	wire vertical_tile_27_26_to_tile_26_26_0;
	wire vertical_tile_27_26_to_tile_26_26_1;
	wire vertical_tile_27_26_to_tile_26_26_2;
	wire vertical_tile_27_26_to_tile_26_26_3;

	wire vertical_tile_26_27_to_tile_27_27_0;
	wire vertical_tile_26_27_to_tile_27_27_1;
	wire vertical_tile_26_27_to_tile_27_27_2;
	wire vertical_tile_26_27_to_tile_27_27_3;
	wire vertical_tile_27_27_to_tile_26_27_0;
	wire vertical_tile_27_27_to_tile_26_27_1;
	wire vertical_tile_27_27_to_tile_26_27_2;
	wire vertical_tile_27_27_to_tile_26_27_3;

	wire vertical_tile_26_28_to_tile_27_28_0;
	wire vertical_tile_26_28_to_tile_27_28_1;
	wire vertical_tile_26_28_to_tile_27_28_2;
	wire vertical_tile_26_28_to_tile_27_28_3;
	wire vertical_tile_27_28_to_tile_26_28_0;
	wire vertical_tile_27_28_to_tile_26_28_1;
	wire vertical_tile_27_28_to_tile_26_28_2;
	wire vertical_tile_27_28_to_tile_26_28_3;

	wire vertical_tile_26_29_to_tile_27_29_0;
	wire vertical_tile_26_29_to_tile_27_29_1;
	wire vertical_tile_26_29_to_tile_27_29_2;
	wire vertical_tile_26_29_to_tile_27_29_3;
	wire vertical_tile_27_29_to_tile_26_29_0;
	wire vertical_tile_27_29_to_tile_26_29_1;
	wire vertical_tile_27_29_to_tile_26_29_2;
	wire vertical_tile_27_29_to_tile_26_29_3;

	wire vertical_tile_26_30_to_tile_27_30_0;
	wire vertical_tile_26_30_to_tile_27_30_1;
	wire vertical_tile_26_30_to_tile_27_30_2;
	wire vertical_tile_26_30_to_tile_27_30_3;
	wire vertical_tile_27_30_to_tile_26_30_0;
	wire vertical_tile_27_30_to_tile_26_30_1;
	wire vertical_tile_27_30_to_tile_26_30_2;
	wire vertical_tile_27_30_to_tile_26_30_3;

	wire vertical_tile_26_31_to_tile_27_31_0;
	wire vertical_tile_26_31_to_tile_27_31_1;
	wire vertical_tile_26_31_to_tile_27_31_2;
	wire vertical_tile_26_31_to_tile_27_31_3;
	wire vertical_tile_27_31_to_tile_26_31_0;
	wire vertical_tile_27_31_to_tile_26_31_1;
	wire vertical_tile_27_31_to_tile_26_31_2;
	wire vertical_tile_27_31_to_tile_26_31_3;

	wire vertical_tile_27_0_to_tile_28_0_0;
	wire vertical_tile_27_0_to_tile_28_0_1;
	wire vertical_tile_27_0_to_tile_28_0_2;
	wire vertical_tile_27_0_to_tile_28_0_3;
	wire vertical_tile_28_0_to_tile_27_0_0;
	wire vertical_tile_28_0_to_tile_27_0_1;
	wire vertical_tile_28_0_to_tile_27_0_2;
	wire vertical_tile_28_0_to_tile_27_0_3;

	wire vertical_tile_27_1_to_tile_28_1_0;
	wire vertical_tile_27_1_to_tile_28_1_1;
	wire vertical_tile_27_1_to_tile_28_1_2;
	wire vertical_tile_27_1_to_tile_28_1_3;
	wire vertical_tile_28_1_to_tile_27_1_0;
	wire vertical_tile_28_1_to_tile_27_1_1;
	wire vertical_tile_28_1_to_tile_27_1_2;
	wire vertical_tile_28_1_to_tile_27_1_3;

	wire vertical_tile_27_2_to_tile_28_2_0;
	wire vertical_tile_27_2_to_tile_28_2_1;
	wire vertical_tile_27_2_to_tile_28_2_2;
	wire vertical_tile_27_2_to_tile_28_2_3;
	wire vertical_tile_28_2_to_tile_27_2_0;
	wire vertical_tile_28_2_to_tile_27_2_1;
	wire vertical_tile_28_2_to_tile_27_2_2;
	wire vertical_tile_28_2_to_tile_27_2_3;

	wire vertical_tile_27_3_to_tile_28_3_0;
	wire vertical_tile_27_3_to_tile_28_3_1;
	wire vertical_tile_27_3_to_tile_28_3_2;
	wire vertical_tile_27_3_to_tile_28_3_3;
	wire vertical_tile_28_3_to_tile_27_3_0;
	wire vertical_tile_28_3_to_tile_27_3_1;
	wire vertical_tile_28_3_to_tile_27_3_2;
	wire vertical_tile_28_3_to_tile_27_3_3;

	wire vertical_tile_27_4_to_tile_28_4_0;
	wire vertical_tile_27_4_to_tile_28_4_1;
	wire vertical_tile_27_4_to_tile_28_4_2;
	wire vertical_tile_27_4_to_tile_28_4_3;
	wire vertical_tile_28_4_to_tile_27_4_0;
	wire vertical_tile_28_4_to_tile_27_4_1;
	wire vertical_tile_28_4_to_tile_27_4_2;
	wire vertical_tile_28_4_to_tile_27_4_3;

	wire vertical_tile_27_5_to_tile_28_5_0;
	wire vertical_tile_27_5_to_tile_28_5_1;
	wire vertical_tile_27_5_to_tile_28_5_2;
	wire vertical_tile_27_5_to_tile_28_5_3;
	wire vertical_tile_28_5_to_tile_27_5_0;
	wire vertical_tile_28_5_to_tile_27_5_1;
	wire vertical_tile_28_5_to_tile_27_5_2;
	wire vertical_tile_28_5_to_tile_27_5_3;

	wire vertical_tile_27_6_to_tile_28_6_0;
	wire vertical_tile_27_6_to_tile_28_6_1;
	wire vertical_tile_27_6_to_tile_28_6_2;
	wire vertical_tile_27_6_to_tile_28_6_3;
	wire vertical_tile_28_6_to_tile_27_6_0;
	wire vertical_tile_28_6_to_tile_27_6_1;
	wire vertical_tile_28_6_to_tile_27_6_2;
	wire vertical_tile_28_6_to_tile_27_6_3;

	wire vertical_tile_27_7_to_tile_28_7_0;
	wire vertical_tile_27_7_to_tile_28_7_1;
	wire vertical_tile_27_7_to_tile_28_7_2;
	wire vertical_tile_27_7_to_tile_28_7_3;
	wire vertical_tile_28_7_to_tile_27_7_0;
	wire vertical_tile_28_7_to_tile_27_7_1;
	wire vertical_tile_28_7_to_tile_27_7_2;
	wire vertical_tile_28_7_to_tile_27_7_3;

	wire vertical_tile_27_8_to_tile_28_8_0;
	wire vertical_tile_27_8_to_tile_28_8_1;
	wire vertical_tile_27_8_to_tile_28_8_2;
	wire vertical_tile_27_8_to_tile_28_8_3;
	wire vertical_tile_28_8_to_tile_27_8_0;
	wire vertical_tile_28_8_to_tile_27_8_1;
	wire vertical_tile_28_8_to_tile_27_8_2;
	wire vertical_tile_28_8_to_tile_27_8_3;

	wire vertical_tile_27_9_to_tile_28_9_0;
	wire vertical_tile_27_9_to_tile_28_9_1;
	wire vertical_tile_27_9_to_tile_28_9_2;
	wire vertical_tile_27_9_to_tile_28_9_3;
	wire vertical_tile_28_9_to_tile_27_9_0;
	wire vertical_tile_28_9_to_tile_27_9_1;
	wire vertical_tile_28_9_to_tile_27_9_2;
	wire vertical_tile_28_9_to_tile_27_9_3;

	wire vertical_tile_27_10_to_tile_28_10_0;
	wire vertical_tile_27_10_to_tile_28_10_1;
	wire vertical_tile_27_10_to_tile_28_10_2;
	wire vertical_tile_27_10_to_tile_28_10_3;
	wire vertical_tile_28_10_to_tile_27_10_0;
	wire vertical_tile_28_10_to_tile_27_10_1;
	wire vertical_tile_28_10_to_tile_27_10_2;
	wire vertical_tile_28_10_to_tile_27_10_3;

	wire vertical_tile_27_11_to_tile_28_11_0;
	wire vertical_tile_27_11_to_tile_28_11_1;
	wire vertical_tile_27_11_to_tile_28_11_2;
	wire vertical_tile_27_11_to_tile_28_11_3;
	wire vertical_tile_28_11_to_tile_27_11_0;
	wire vertical_tile_28_11_to_tile_27_11_1;
	wire vertical_tile_28_11_to_tile_27_11_2;
	wire vertical_tile_28_11_to_tile_27_11_3;

	wire vertical_tile_27_12_to_tile_28_12_0;
	wire vertical_tile_27_12_to_tile_28_12_1;
	wire vertical_tile_27_12_to_tile_28_12_2;
	wire vertical_tile_27_12_to_tile_28_12_3;
	wire vertical_tile_28_12_to_tile_27_12_0;
	wire vertical_tile_28_12_to_tile_27_12_1;
	wire vertical_tile_28_12_to_tile_27_12_2;
	wire vertical_tile_28_12_to_tile_27_12_3;

	wire vertical_tile_27_13_to_tile_28_13_0;
	wire vertical_tile_27_13_to_tile_28_13_1;
	wire vertical_tile_27_13_to_tile_28_13_2;
	wire vertical_tile_27_13_to_tile_28_13_3;
	wire vertical_tile_28_13_to_tile_27_13_0;
	wire vertical_tile_28_13_to_tile_27_13_1;
	wire vertical_tile_28_13_to_tile_27_13_2;
	wire vertical_tile_28_13_to_tile_27_13_3;

	wire vertical_tile_27_14_to_tile_28_14_0;
	wire vertical_tile_27_14_to_tile_28_14_1;
	wire vertical_tile_27_14_to_tile_28_14_2;
	wire vertical_tile_27_14_to_tile_28_14_3;
	wire vertical_tile_28_14_to_tile_27_14_0;
	wire vertical_tile_28_14_to_tile_27_14_1;
	wire vertical_tile_28_14_to_tile_27_14_2;
	wire vertical_tile_28_14_to_tile_27_14_3;

	wire vertical_tile_27_15_to_tile_28_15_0;
	wire vertical_tile_27_15_to_tile_28_15_1;
	wire vertical_tile_27_15_to_tile_28_15_2;
	wire vertical_tile_27_15_to_tile_28_15_3;
	wire vertical_tile_28_15_to_tile_27_15_0;
	wire vertical_tile_28_15_to_tile_27_15_1;
	wire vertical_tile_28_15_to_tile_27_15_2;
	wire vertical_tile_28_15_to_tile_27_15_3;

	wire vertical_tile_27_16_to_tile_28_16_0;
	wire vertical_tile_27_16_to_tile_28_16_1;
	wire vertical_tile_27_16_to_tile_28_16_2;
	wire vertical_tile_27_16_to_tile_28_16_3;
	wire vertical_tile_28_16_to_tile_27_16_0;
	wire vertical_tile_28_16_to_tile_27_16_1;
	wire vertical_tile_28_16_to_tile_27_16_2;
	wire vertical_tile_28_16_to_tile_27_16_3;

	wire vertical_tile_27_17_to_tile_28_17_0;
	wire vertical_tile_27_17_to_tile_28_17_1;
	wire vertical_tile_27_17_to_tile_28_17_2;
	wire vertical_tile_27_17_to_tile_28_17_3;
	wire vertical_tile_28_17_to_tile_27_17_0;
	wire vertical_tile_28_17_to_tile_27_17_1;
	wire vertical_tile_28_17_to_tile_27_17_2;
	wire vertical_tile_28_17_to_tile_27_17_3;

	wire vertical_tile_27_18_to_tile_28_18_0;
	wire vertical_tile_27_18_to_tile_28_18_1;
	wire vertical_tile_27_18_to_tile_28_18_2;
	wire vertical_tile_27_18_to_tile_28_18_3;
	wire vertical_tile_28_18_to_tile_27_18_0;
	wire vertical_tile_28_18_to_tile_27_18_1;
	wire vertical_tile_28_18_to_tile_27_18_2;
	wire vertical_tile_28_18_to_tile_27_18_3;

	wire vertical_tile_27_19_to_tile_28_19_0;
	wire vertical_tile_27_19_to_tile_28_19_1;
	wire vertical_tile_27_19_to_tile_28_19_2;
	wire vertical_tile_27_19_to_tile_28_19_3;
	wire vertical_tile_28_19_to_tile_27_19_0;
	wire vertical_tile_28_19_to_tile_27_19_1;
	wire vertical_tile_28_19_to_tile_27_19_2;
	wire vertical_tile_28_19_to_tile_27_19_3;

	wire vertical_tile_27_20_to_tile_28_20_0;
	wire vertical_tile_27_20_to_tile_28_20_1;
	wire vertical_tile_27_20_to_tile_28_20_2;
	wire vertical_tile_27_20_to_tile_28_20_3;
	wire vertical_tile_28_20_to_tile_27_20_0;
	wire vertical_tile_28_20_to_tile_27_20_1;
	wire vertical_tile_28_20_to_tile_27_20_2;
	wire vertical_tile_28_20_to_tile_27_20_3;

	wire vertical_tile_27_21_to_tile_28_21_0;
	wire vertical_tile_27_21_to_tile_28_21_1;
	wire vertical_tile_27_21_to_tile_28_21_2;
	wire vertical_tile_27_21_to_tile_28_21_3;
	wire vertical_tile_28_21_to_tile_27_21_0;
	wire vertical_tile_28_21_to_tile_27_21_1;
	wire vertical_tile_28_21_to_tile_27_21_2;
	wire vertical_tile_28_21_to_tile_27_21_3;

	wire vertical_tile_27_22_to_tile_28_22_0;
	wire vertical_tile_27_22_to_tile_28_22_1;
	wire vertical_tile_27_22_to_tile_28_22_2;
	wire vertical_tile_27_22_to_tile_28_22_3;
	wire vertical_tile_28_22_to_tile_27_22_0;
	wire vertical_tile_28_22_to_tile_27_22_1;
	wire vertical_tile_28_22_to_tile_27_22_2;
	wire vertical_tile_28_22_to_tile_27_22_3;

	wire vertical_tile_27_23_to_tile_28_23_0;
	wire vertical_tile_27_23_to_tile_28_23_1;
	wire vertical_tile_27_23_to_tile_28_23_2;
	wire vertical_tile_27_23_to_tile_28_23_3;
	wire vertical_tile_28_23_to_tile_27_23_0;
	wire vertical_tile_28_23_to_tile_27_23_1;
	wire vertical_tile_28_23_to_tile_27_23_2;
	wire vertical_tile_28_23_to_tile_27_23_3;

	wire vertical_tile_27_24_to_tile_28_24_0;
	wire vertical_tile_27_24_to_tile_28_24_1;
	wire vertical_tile_27_24_to_tile_28_24_2;
	wire vertical_tile_27_24_to_tile_28_24_3;
	wire vertical_tile_28_24_to_tile_27_24_0;
	wire vertical_tile_28_24_to_tile_27_24_1;
	wire vertical_tile_28_24_to_tile_27_24_2;
	wire vertical_tile_28_24_to_tile_27_24_3;

	wire vertical_tile_27_25_to_tile_28_25_0;
	wire vertical_tile_27_25_to_tile_28_25_1;
	wire vertical_tile_27_25_to_tile_28_25_2;
	wire vertical_tile_27_25_to_tile_28_25_3;
	wire vertical_tile_28_25_to_tile_27_25_0;
	wire vertical_tile_28_25_to_tile_27_25_1;
	wire vertical_tile_28_25_to_tile_27_25_2;
	wire vertical_tile_28_25_to_tile_27_25_3;

	wire vertical_tile_27_26_to_tile_28_26_0;
	wire vertical_tile_27_26_to_tile_28_26_1;
	wire vertical_tile_27_26_to_tile_28_26_2;
	wire vertical_tile_27_26_to_tile_28_26_3;
	wire vertical_tile_28_26_to_tile_27_26_0;
	wire vertical_tile_28_26_to_tile_27_26_1;
	wire vertical_tile_28_26_to_tile_27_26_2;
	wire vertical_tile_28_26_to_tile_27_26_3;

	wire vertical_tile_27_27_to_tile_28_27_0;
	wire vertical_tile_27_27_to_tile_28_27_1;
	wire vertical_tile_27_27_to_tile_28_27_2;
	wire vertical_tile_27_27_to_tile_28_27_3;
	wire vertical_tile_28_27_to_tile_27_27_0;
	wire vertical_tile_28_27_to_tile_27_27_1;
	wire vertical_tile_28_27_to_tile_27_27_2;
	wire vertical_tile_28_27_to_tile_27_27_3;

	wire vertical_tile_27_28_to_tile_28_28_0;
	wire vertical_tile_27_28_to_tile_28_28_1;
	wire vertical_tile_27_28_to_tile_28_28_2;
	wire vertical_tile_27_28_to_tile_28_28_3;
	wire vertical_tile_28_28_to_tile_27_28_0;
	wire vertical_tile_28_28_to_tile_27_28_1;
	wire vertical_tile_28_28_to_tile_27_28_2;
	wire vertical_tile_28_28_to_tile_27_28_3;

	wire vertical_tile_27_29_to_tile_28_29_0;
	wire vertical_tile_27_29_to_tile_28_29_1;
	wire vertical_tile_27_29_to_tile_28_29_2;
	wire vertical_tile_27_29_to_tile_28_29_3;
	wire vertical_tile_28_29_to_tile_27_29_0;
	wire vertical_tile_28_29_to_tile_27_29_1;
	wire vertical_tile_28_29_to_tile_27_29_2;
	wire vertical_tile_28_29_to_tile_27_29_3;

	wire vertical_tile_27_30_to_tile_28_30_0;
	wire vertical_tile_27_30_to_tile_28_30_1;
	wire vertical_tile_27_30_to_tile_28_30_2;
	wire vertical_tile_27_30_to_tile_28_30_3;
	wire vertical_tile_28_30_to_tile_27_30_0;
	wire vertical_tile_28_30_to_tile_27_30_1;
	wire vertical_tile_28_30_to_tile_27_30_2;
	wire vertical_tile_28_30_to_tile_27_30_3;

	wire vertical_tile_27_31_to_tile_28_31_0;
	wire vertical_tile_27_31_to_tile_28_31_1;
	wire vertical_tile_27_31_to_tile_28_31_2;
	wire vertical_tile_27_31_to_tile_28_31_3;
	wire vertical_tile_28_31_to_tile_27_31_0;
	wire vertical_tile_28_31_to_tile_27_31_1;
	wire vertical_tile_28_31_to_tile_27_31_2;
	wire vertical_tile_28_31_to_tile_27_31_3;

	wire vertical_tile_28_0_to_tile_29_0_0;
	wire vertical_tile_28_0_to_tile_29_0_1;
	wire vertical_tile_28_0_to_tile_29_0_2;
	wire vertical_tile_28_0_to_tile_29_0_3;
	wire vertical_tile_29_0_to_tile_28_0_0;
	wire vertical_tile_29_0_to_tile_28_0_1;
	wire vertical_tile_29_0_to_tile_28_0_2;
	wire vertical_tile_29_0_to_tile_28_0_3;

	wire vertical_tile_28_1_to_tile_29_1_0;
	wire vertical_tile_28_1_to_tile_29_1_1;
	wire vertical_tile_28_1_to_tile_29_1_2;
	wire vertical_tile_28_1_to_tile_29_1_3;
	wire vertical_tile_29_1_to_tile_28_1_0;
	wire vertical_tile_29_1_to_tile_28_1_1;
	wire vertical_tile_29_1_to_tile_28_1_2;
	wire vertical_tile_29_1_to_tile_28_1_3;

	wire vertical_tile_28_2_to_tile_29_2_0;
	wire vertical_tile_28_2_to_tile_29_2_1;
	wire vertical_tile_28_2_to_tile_29_2_2;
	wire vertical_tile_28_2_to_tile_29_2_3;
	wire vertical_tile_29_2_to_tile_28_2_0;
	wire vertical_tile_29_2_to_tile_28_2_1;
	wire vertical_tile_29_2_to_tile_28_2_2;
	wire vertical_tile_29_2_to_tile_28_2_3;

	wire vertical_tile_28_3_to_tile_29_3_0;
	wire vertical_tile_28_3_to_tile_29_3_1;
	wire vertical_tile_28_3_to_tile_29_3_2;
	wire vertical_tile_28_3_to_tile_29_3_3;
	wire vertical_tile_29_3_to_tile_28_3_0;
	wire vertical_tile_29_3_to_tile_28_3_1;
	wire vertical_tile_29_3_to_tile_28_3_2;
	wire vertical_tile_29_3_to_tile_28_3_3;

	wire vertical_tile_28_4_to_tile_29_4_0;
	wire vertical_tile_28_4_to_tile_29_4_1;
	wire vertical_tile_28_4_to_tile_29_4_2;
	wire vertical_tile_28_4_to_tile_29_4_3;
	wire vertical_tile_29_4_to_tile_28_4_0;
	wire vertical_tile_29_4_to_tile_28_4_1;
	wire vertical_tile_29_4_to_tile_28_4_2;
	wire vertical_tile_29_4_to_tile_28_4_3;

	wire vertical_tile_28_5_to_tile_29_5_0;
	wire vertical_tile_28_5_to_tile_29_5_1;
	wire vertical_tile_28_5_to_tile_29_5_2;
	wire vertical_tile_28_5_to_tile_29_5_3;
	wire vertical_tile_29_5_to_tile_28_5_0;
	wire vertical_tile_29_5_to_tile_28_5_1;
	wire vertical_tile_29_5_to_tile_28_5_2;
	wire vertical_tile_29_5_to_tile_28_5_3;

	wire vertical_tile_28_6_to_tile_29_6_0;
	wire vertical_tile_28_6_to_tile_29_6_1;
	wire vertical_tile_28_6_to_tile_29_6_2;
	wire vertical_tile_28_6_to_tile_29_6_3;
	wire vertical_tile_29_6_to_tile_28_6_0;
	wire vertical_tile_29_6_to_tile_28_6_1;
	wire vertical_tile_29_6_to_tile_28_6_2;
	wire vertical_tile_29_6_to_tile_28_6_3;

	wire vertical_tile_28_7_to_tile_29_7_0;
	wire vertical_tile_28_7_to_tile_29_7_1;
	wire vertical_tile_28_7_to_tile_29_7_2;
	wire vertical_tile_28_7_to_tile_29_7_3;
	wire vertical_tile_29_7_to_tile_28_7_0;
	wire vertical_tile_29_7_to_tile_28_7_1;
	wire vertical_tile_29_7_to_tile_28_7_2;
	wire vertical_tile_29_7_to_tile_28_7_3;

	wire vertical_tile_28_8_to_tile_29_8_0;
	wire vertical_tile_28_8_to_tile_29_8_1;
	wire vertical_tile_28_8_to_tile_29_8_2;
	wire vertical_tile_28_8_to_tile_29_8_3;
	wire vertical_tile_29_8_to_tile_28_8_0;
	wire vertical_tile_29_8_to_tile_28_8_1;
	wire vertical_tile_29_8_to_tile_28_8_2;
	wire vertical_tile_29_8_to_tile_28_8_3;

	wire vertical_tile_28_9_to_tile_29_9_0;
	wire vertical_tile_28_9_to_tile_29_9_1;
	wire vertical_tile_28_9_to_tile_29_9_2;
	wire vertical_tile_28_9_to_tile_29_9_3;
	wire vertical_tile_29_9_to_tile_28_9_0;
	wire vertical_tile_29_9_to_tile_28_9_1;
	wire vertical_tile_29_9_to_tile_28_9_2;
	wire vertical_tile_29_9_to_tile_28_9_3;

	wire vertical_tile_28_10_to_tile_29_10_0;
	wire vertical_tile_28_10_to_tile_29_10_1;
	wire vertical_tile_28_10_to_tile_29_10_2;
	wire vertical_tile_28_10_to_tile_29_10_3;
	wire vertical_tile_29_10_to_tile_28_10_0;
	wire vertical_tile_29_10_to_tile_28_10_1;
	wire vertical_tile_29_10_to_tile_28_10_2;
	wire vertical_tile_29_10_to_tile_28_10_3;

	wire vertical_tile_28_11_to_tile_29_11_0;
	wire vertical_tile_28_11_to_tile_29_11_1;
	wire vertical_tile_28_11_to_tile_29_11_2;
	wire vertical_tile_28_11_to_tile_29_11_3;
	wire vertical_tile_29_11_to_tile_28_11_0;
	wire vertical_tile_29_11_to_tile_28_11_1;
	wire vertical_tile_29_11_to_tile_28_11_2;
	wire vertical_tile_29_11_to_tile_28_11_3;

	wire vertical_tile_28_12_to_tile_29_12_0;
	wire vertical_tile_28_12_to_tile_29_12_1;
	wire vertical_tile_28_12_to_tile_29_12_2;
	wire vertical_tile_28_12_to_tile_29_12_3;
	wire vertical_tile_29_12_to_tile_28_12_0;
	wire vertical_tile_29_12_to_tile_28_12_1;
	wire vertical_tile_29_12_to_tile_28_12_2;
	wire vertical_tile_29_12_to_tile_28_12_3;

	wire vertical_tile_28_13_to_tile_29_13_0;
	wire vertical_tile_28_13_to_tile_29_13_1;
	wire vertical_tile_28_13_to_tile_29_13_2;
	wire vertical_tile_28_13_to_tile_29_13_3;
	wire vertical_tile_29_13_to_tile_28_13_0;
	wire vertical_tile_29_13_to_tile_28_13_1;
	wire vertical_tile_29_13_to_tile_28_13_2;
	wire vertical_tile_29_13_to_tile_28_13_3;

	wire vertical_tile_28_14_to_tile_29_14_0;
	wire vertical_tile_28_14_to_tile_29_14_1;
	wire vertical_tile_28_14_to_tile_29_14_2;
	wire vertical_tile_28_14_to_tile_29_14_3;
	wire vertical_tile_29_14_to_tile_28_14_0;
	wire vertical_tile_29_14_to_tile_28_14_1;
	wire vertical_tile_29_14_to_tile_28_14_2;
	wire vertical_tile_29_14_to_tile_28_14_3;

	wire vertical_tile_28_15_to_tile_29_15_0;
	wire vertical_tile_28_15_to_tile_29_15_1;
	wire vertical_tile_28_15_to_tile_29_15_2;
	wire vertical_tile_28_15_to_tile_29_15_3;
	wire vertical_tile_29_15_to_tile_28_15_0;
	wire vertical_tile_29_15_to_tile_28_15_1;
	wire vertical_tile_29_15_to_tile_28_15_2;
	wire vertical_tile_29_15_to_tile_28_15_3;

	wire vertical_tile_28_16_to_tile_29_16_0;
	wire vertical_tile_28_16_to_tile_29_16_1;
	wire vertical_tile_28_16_to_tile_29_16_2;
	wire vertical_tile_28_16_to_tile_29_16_3;
	wire vertical_tile_29_16_to_tile_28_16_0;
	wire vertical_tile_29_16_to_tile_28_16_1;
	wire vertical_tile_29_16_to_tile_28_16_2;
	wire vertical_tile_29_16_to_tile_28_16_3;

	wire vertical_tile_28_17_to_tile_29_17_0;
	wire vertical_tile_28_17_to_tile_29_17_1;
	wire vertical_tile_28_17_to_tile_29_17_2;
	wire vertical_tile_28_17_to_tile_29_17_3;
	wire vertical_tile_29_17_to_tile_28_17_0;
	wire vertical_tile_29_17_to_tile_28_17_1;
	wire vertical_tile_29_17_to_tile_28_17_2;
	wire vertical_tile_29_17_to_tile_28_17_3;

	wire vertical_tile_28_18_to_tile_29_18_0;
	wire vertical_tile_28_18_to_tile_29_18_1;
	wire vertical_tile_28_18_to_tile_29_18_2;
	wire vertical_tile_28_18_to_tile_29_18_3;
	wire vertical_tile_29_18_to_tile_28_18_0;
	wire vertical_tile_29_18_to_tile_28_18_1;
	wire vertical_tile_29_18_to_tile_28_18_2;
	wire vertical_tile_29_18_to_tile_28_18_3;

	wire vertical_tile_28_19_to_tile_29_19_0;
	wire vertical_tile_28_19_to_tile_29_19_1;
	wire vertical_tile_28_19_to_tile_29_19_2;
	wire vertical_tile_28_19_to_tile_29_19_3;
	wire vertical_tile_29_19_to_tile_28_19_0;
	wire vertical_tile_29_19_to_tile_28_19_1;
	wire vertical_tile_29_19_to_tile_28_19_2;
	wire vertical_tile_29_19_to_tile_28_19_3;

	wire vertical_tile_28_20_to_tile_29_20_0;
	wire vertical_tile_28_20_to_tile_29_20_1;
	wire vertical_tile_28_20_to_tile_29_20_2;
	wire vertical_tile_28_20_to_tile_29_20_3;
	wire vertical_tile_29_20_to_tile_28_20_0;
	wire vertical_tile_29_20_to_tile_28_20_1;
	wire vertical_tile_29_20_to_tile_28_20_2;
	wire vertical_tile_29_20_to_tile_28_20_3;

	wire vertical_tile_28_21_to_tile_29_21_0;
	wire vertical_tile_28_21_to_tile_29_21_1;
	wire vertical_tile_28_21_to_tile_29_21_2;
	wire vertical_tile_28_21_to_tile_29_21_3;
	wire vertical_tile_29_21_to_tile_28_21_0;
	wire vertical_tile_29_21_to_tile_28_21_1;
	wire vertical_tile_29_21_to_tile_28_21_2;
	wire vertical_tile_29_21_to_tile_28_21_3;

	wire vertical_tile_28_22_to_tile_29_22_0;
	wire vertical_tile_28_22_to_tile_29_22_1;
	wire vertical_tile_28_22_to_tile_29_22_2;
	wire vertical_tile_28_22_to_tile_29_22_3;
	wire vertical_tile_29_22_to_tile_28_22_0;
	wire vertical_tile_29_22_to_tile_28_22_1;
	wire vertical_tile_29_22_to_tile_28_22_2;
	wire vertical_tile_29_22_to_tile_28_22_3;

	wire vertical_tile_28_23_to_tile_29_23_0;
	wire vertical_tile_28_23_to_tile_29_23_1;
	wire vertical_tile_28_23_to_tile_29_23_2;
	wire vertical_tile_28_23_to_tile_29_23_3;
	wire vertical_tile_29_23_to_tile_28_23_0;
	wire vertical_tile_29_23_to_tile_28_23_1;
	wire vertical_tile_29_23_to_tile_28_23_2;
	wire vertical_tile_29_23_to_tile_28_23_3;

	wire vertical_tile_28_24_to_tile_29_24_0;
	wire vertical_tile_28_24_to_tile_29_24_1;
	wire vertical_tile_28_24_to_tile_29_24_2;
	wire vertical_tile_28_24_to_tile_29_24_3;
	wire vertical_tile_29_24_to_tile_28_24_0;
	wire vertical_tile_29_24_to_tile_28_24_1;
	wire vertical_tile_29_24_to_tile_28_24_2;
	wire vertical_tile_29_24_to_tile_28_24_3;

	wire vertical_tile_28_25_to_tile_29_25_0;
	wire vertical_tile_28_25_to_tile_29_25_1;
	wire vertical_tile_28_25_to_tile_29_25_2;
	wire vertical_tile_28_25_to_tile_29_25_3;
	wire vertical_tile_29_25_to_tile_28_25_0;
	wire vertical_tile_29_25_to_tile_28_25_1;
	wire vertical_tile_29_25_to_tile_28_25_2;
	wire vertical_tile_29_25_to_tile_28_25_3;

	wire vertical_tile_28_26_to_tile_29_26_0;
	wire vertical_tile_28_26_to_tile_29_26_1;
	wire vertical_tile_28_26_to_tile_29_26_2;
	wire vertical_tile_28_26_to_tile_29_26_3;
	wire vertical_tile_29_26_to_tile_28_26_0;
	wire vertical_tile_29_26_to_tile_28_26_1;
	wire vertical_tile_29_26_to_tile_28_26_2;
	wire vertical_tile_29_26_to_tile_28_26_3;

	wire vertical_tile_28_27_to_tile_29_27_0;
	wire vertical_tile_28_27_to_tile_29_27_1;
	wire vertical_tile_28_27_to_tile_29_27_2;
	wire vertical_tile_28_27_to_tile_29_27_3;
	wire vertical_tile_29_27_to_tile_28_27_0;
	wire vertical_tile_29_27_to_tile_28_27_1;
	wire vertical_tile_29_27_to_tile_28_27_2;
	wire vertical_tile_29_27_to_tile_28_27_3;

	wire vertical_tile_28_28_to_tile_29_28_0;
	wire vertical_tile_28_28_to_tile_29_28_1;
	wire vertical_tile_28_28_to_tile_29_28_2;
	wire vertical_tile_28_28_to_tile_29_28_3;
	wire vertical_tile_29_28_to_tile_28_28_0;
	wire vertical_tile_29_28_to_tile_28_28_1;
	wire vertical_tile_29_28_to_tile_28_28_2;
	wire vertical_tile_29_28_to_tile_28_28_3;

	wire vertical_tile_28_29_to_tile_29_29_0;
	wire vertical_tile_28_29_to_tile_29_29_1;
	wire vertical_tile_28_29_to_tile_29_29_2;
	wire vertical_tile_28_29_to_tile_29_29_3;
	wire vertical_tile_29_29_to_tile_28_29_0;
	wire vertical_tile_29_29_to_tile_28_29_1;
	wire vertical_tile_29_29_to_tile_28_29_2;
	wire vertical_tile_29_29_to_tile_28_29_3;

	wire vertical_tile_28_30_to_tile_29_30_0;
	wire vertical_tile_28_30_to_tile_29_30_1;
	wire vertical_tile_28_30_to_tile_29_30_2;
	wire vertical_tile_28_30_to_tile_29_30_3;
	wire vertical_tile_29_30_to_tile_28_30_0;
	wire vertical_tile_29_30_to_tile_28_30_1;
	wire vertical_tile_29_30_to_tile_28_30_2;
	wire vertical_tile_29_30_to_tile_28_30_3;

	wire vertical_tile_28_31_to_tile_29_31_0;
	wire vertical_tile_28_31_to_tile_29_31_1;
	wire vertical_tile_28_31_to_tile_29_31_2;
	wire vertical_tile_28_31_to_tile_29_31_3;
	wire vertical_tile_29_31_to_tile_28_31_0;
	wire vertical_tile_29_31_to_tile_28_31_1;
	wire vertical_tile_29_31_to_tile_28_31_2;
	wire vertical_tile_29_31_to_tile_28_31_3;

	wire vertical_tile_29_0_to_tile_30_0_0;
	wire vertical_tile_29_0_to_tile_30_0_1;
	wire vertical_tile_29_0_to_tile_30_0_2;
	wire vertical_tile_29_0_to_tile_30_0_3;
	wire vertical_tile_30_0_to_tile_29_0_0;
	wire vertical_tile_30_0_to_tile_29_0_1;
	wire vertical_tile_30_0_to_tile_29_0_2;
	wire vertical_tile_30_0_to_tile_29_0_3;

	wire vertical_tile_29_1_to_tile_30_1_0;
	wire vertical_tile_29_1_to_tile_30_1_1;
	wire vertical_tile_29_1_to_tile_30_1_2;
	wire vertical_tile_29_1_to_tile_30_1_3;
	wire vertical_tile_30_1_to_tile_29_1_0;
	wire vertical_tile_30_1_to_tile_29_1_1;
	wire vertical_tile_30_1_to_tile_29_1_2;
	wire vertical_tile_30_1_to_tile_29_1_3;

	wire vertical_tile_29_2_to_tile_30_2_0;
	wire vertical_tile_29_2_to_tile_30_2_1;
	wire vertical_tile_29_2_to_tile_30_2_2;
	wire vertical_tile_29_2_to_tile_30_2_3;
	wire vertical_tile_30_2_to_tile_29_2_0;
	wire vertical_tile_30_2_to_tile_29_2_1;
	wire vertical_tile_30_2_to_tile_29_2_2;
	wire vertical_tile_30_2_to_tile_29_2_3;

	wire vertical_tile_29_3_to_tile_30_3_0;
	wire vertical_tile_29_3_to_tile_30_3_1;
	wire vertical_tile_29_3_to_tile_30_3_2;
	wire vertical_tile_29_3_to_tile_30_3_3;
	wire vertical_tile_30_3_to_tile_29_3_0;
	wire vertical_tile_30_3_to_tile_29_3_1;
	wire vertical_tile_30_3_to_tile_29_3_2;
	wire vertical_tile_30_3_to_tile_29_3_3;

	wire vertical_tile_29_4_to_tile_30_4_0;
	wire vertical_tile_29_4_to_tile_30_4_1;
	wire vertical_tile_29_4_to_tile_30_4_2;
	wire vertical_tile_29_4_to_tile_30_4_3;
	wire vertical_tile_30_4_to_tile_29_4_0;
	wire vertical_tile_30_4_to_tile_29_4_1;
	wire vertical_tile_30_4_to_tile_29_4_2;
	wire vertical_tile_30_4_to_tile_29_4_3;

	wire vertical_tile_29_5_to_tile_30_5_0;
	wire vertical_tile_29_5_to_tile_30_5_1;
	wire vertical_tile_29_5_to_tile_30_5_2;
	wire vertical_tile_29_5_to_tile_30_5_3;
	wire vertical_tile_30_5_to_tile_29_5_0;
	wire vertical_tile_30_5_to_tile_29_5_1;
	wire vertical_tile_30_5_to_tile_29_5_2;
	wire vertical_tile_30_5_to_tile_29_5_3;

	wire vertical_tile_29_6_to_tile_30_6_0;
	wire vertical_tile_29_6_to_tile_30_6_1;
	wire vertical_tile_29_6_to_tile_30_6_2;
	wire vertical_tile_29_6_to_tile_30_6_3;
	wire vertical_tile_30_6_to_tile_29_6_0;
	wire vertical_tile_30_6_to_tile_29_6_1;
	wire vertical_tile_30_6_to_tile_29_6_2;
	wire vertical_tile_30_6_to_tile_29_6_3;

	wire vertical_tile_29_7_to_tile_30_7_0;
	wire vertical_tile_29_7_to_tile_30_7_1;
	wire vertical_tile_29_7_to_tile_30_7_2;
	wire vertical_tile_29_7_to_tile_30_7_3;
	wire vertical_tile_30_7_to_tile_29_7_0;
	wire vertical_tile_30_7_to_tile_29_7_1;
	wire vertical_tile_30_7_to_tile_29_7_2;
	wire vertical_tile_30_7_to_tile_29_7_3;

	wire vertical_tile_29_8_to_tile_30_8_0;
	wire vertical_tile_29_8_to_tile_30_8_1;
	wire vertical_tile_29_8_to_tile_30_8_2;
	wire vertical_tile_29_8_to_tile_30_8_3;
	wire vertical_tile_30_8_to_tile_29_8_0;
	wire vertical_tile_30_8_to_tile_29_8_1;
	wire vertical_tile_30_8_to_tile_29_8_2;
	wire vertical_tile_30_8_to_tile_29_8_3;

	wire vertical_tile_29_9_to_tile_30_9_0;
	wire vertical_tile_29_9_to_tile_30_9_1;
	wire vertical_tile_29_9_to_tile_30_9_2;
	wire vertical_tile_29_9_to_tile_30_9_3;
	wire vertical_tile_30_9_to_tile_29_9_0;
	wire vertical_tile_30_9_to_tile_29_9_1;
	wire vertical_tile_30_9_to_tile_29_9_2;
	wire vertical_tile_30_9_to_tile_29_9_3;

	wire vertical_tile_29_10_to_tile_30_10_0;
	wire vertical_tile_29_10_to_tile_30_10_1;
	wire vertical_tile_29_10_to_tile_30_10_2;
	wire vertical_tile_29_10_to_tile_30_10_3;
	wire vertical_tile_30_10_to_tile_29_10_0;
	wire vertical_tile_30_10_to_tile_29_10_1;
	wire vertical_tile_30_10_to_tile_29_10_2;
	wire vertical_tile_30_10_to_tile_29_10_3;

	wire vertical_tile_29_11_to_tile_30_11_0;
	wire vertical_tile_29_11_to_tile_30_11_1;
	wire vertical_tile_29_11_to_tile_30_11_2;
	wire vertical_tile_29_11_to_tile_30_11_3;
	wire vertical_tile_30_11_to_tile_29_11_0;
	wire vertical_tile_30_11_to_tile_29_11_1;
	wire vertical_tile_30_11_to_tile_29_11_2;
	wire vertical_tile_30_11_to_tile_29_11_3;

	wire vertical_tile_29_12_to_tile_30_12_0;
	wire vertical_tile_29_12_to_tile_30_12_1;
	wire vertical_tile_29_12_to_tile_30_12_2;
	wire vertical_tile_29_12_to_tile_30_12_3;
	wire vertical_tile_30_12_to_tile_29_12_0;
	wire vertical_tile_30_12_to_tile_29_12_1;
	wire vertical_tile_30_12_to_tile_29_12_2;
	wire vertical_tile_30_12_to_tile_29_12_3;

	wire vertical_tile_29_13_to_tile_30_13_0;
	wire vertical_tile_29_13_to_tile_30_13_1;
	wire vertical_tile_29_13_to_tile_30_13_2;
	wire vertical_tile_29_13_to_tile_30_13_3;
	wire vertical_tile_30_13_to_tile_29_13_0;
	wire vertical_tile_30_13_to_tile_29_13_1;
	wire vertical_tile_30_13_to_tile_29_13_2;
	wire vertical_tile_30_13_to_tile_29_13_3;

	wire vertical_tile_29_14_to_tile_30_14_0;
	wire vertical_tile_29_14_to_tile_30_14_1;
	wire vertical_tile_29_14_to_tile_30_14_2;
	wire vertical_tile_29_14_to_tile_30_14_3;
	wire vertical_tile_30_14_to_tile_29_14_0;
	wire vertical_tile_30_14_to_tile_29_14_1;
	wire vertical_tile_30_14_to_tile_29_14_2;
	wire vertical_tile_30_14_to_tile_29_14_3;

	wire vertical_tile_29_15_to_tile_30_15_0;
	wire vertical_tile_29_15_to_tile_30_15_1;
	wire vertical_tile_29_15_to_tile_30_15_2;
	wire vertical_tile_29_15_to_tile_30_15_3;
	wire vertical_tile_30_15_to_tile_29_15_0;
	wire vertical_tile_30_15_to_tile_29_15_1;
	wire vertical_tile_30_15_to_tile_29_15_2;
	wire vertical_tile_30_15_to_tile_29_15_3;

	wire vertical_tile_29_16_to_tile_30_16_0;
	wire vertical_tile_29_16_to_tile_30_16_1;
	wire vertical_tile_29_16_to_tile_30_16_2;
	wire vertical_tile_29_16_to_tile_30_16_3;
	wire vertical_tile_30_16_to_tile_29_16_0;
	wire vertical_tile_30_16_to_tile_29_16_1;
	wire vertical_tile_30_16_to_tile_29_16_2;
	wire vertical_tile_30_16_to_tile_29_16_3;

	wire vertical_tile_29_17_to_tile_30_17_0;
	wire vertical_tile_29_17_to_tile_30_17_1;
	wire vertical_tile_29_17_to_tile_30_17_2;
	wire vertical_tile_29_17_to_tile_30_17_3;
	wire vertical_tile_30_17_to_tile_29_17_0;
	wire vertical_tile_30_17_to_tile_29_17_1;
	wire vertical_tile_30_17_to_tile_29_17_2;
	wire vertical_tile_30_17_to_tile_29_17_3;

	wire vertical_tile_29_18_to_tile_30_18_0;
	wire vertical_tile_29_18_to_tile_30_18_1;
	wire vertical_tile_29_18_to_tile_30_18_2;
	wire vertical_tile_29_18_to_tile_30_18_3;
	wire vertical_tile_30_18_to_tile_29_18_0;
	wire vertical_tile_30_18_to_tile_29_18_1;
	wire vertical_tile_30_18_to_tile_29_18_2;
	wire vertical_tile_30_18_to_tile_29_18_3;

	wire vertical_tile_29_19_to_tile_30_19_0;
	wire vertical_tile_29_19_to_tile_30_19_1;
	wire vertical_tile_29_19_to_tile_30_19_2;
	wire vertical_tile_29_19_to_tile_30_19_3;
	wire vertical_tile_30_19_to_tile_29_19_0;
	wire vertical_tile_30_19_to_tile_29_19_1;
	wire vertical_tile_30_19_to_tile_29_19_2;
	wire vertical_tile_30_19_to_tile_29_19_3;

	wire vertical_tile_29_20_to_tile_30_20_0;
	wire vertical_tile_29_20_to_tile_30_20_1;
	wire vertical_tile_29_20_to_tile_30_20_2;
	wire vertical_tile_29_20_to_tile_30_20_3;
	wire vertical_tile_30_20_to_tile_29_20_0;
	wire vertical_tile_30_20_to_tile_29_20_1;
	wire vertical_tile_30_20_to_tile_29_20_2;
	wire vertical_tile_30_20_to_tile_29_20_3;

	wire vertical_tile_29_21_to_tile_30_21_0;
	wire vertical_tile_29_21_to_tile_30_21_1;
	wire vertical_tile_29_21_to_tile_30_21_2;
	wire vertical_tile_29_21_to_tile_30_21_3;
	wire vertical_tile_30_21_to_tile_29_21_0;
	wire vertical_tile_30_21_to_tile_29_21_1;
	wire vertical_tile_30_21_to_tile_29_21_2;
	wire vertical_tile_30_21_to_tile_29_21_3;

	wire vertical_tile_29_22_to_tile_30_22_0;
	wire vertical_tile_29_22_to_tile_30_22_1;
	wire vertical_tile_29_22_to_tile_30_22_2;
	wire vertical_tile_29_22_to_tile_30_22_3;
	wire vertical_tile_30_22_to_tile_29_22_0;
	wire vertical_tile_30_22_to_tile_29_22_1;
	wire vertical_tile_30_22_to_tile_29_22_2;
	wire vertical_tile_30_22_to_tile_29_22_3;

	wire vertical_tile_29_23_to_tile_30_23_0;
	wire vertical_tile_29_23_to_tile_30_23_1;
	wire vertical_tile_29_23_to_tile_30_23_2;
	wire vertical_tile_29_23_to_tile_30_23_3;
	wire vertical_tile_30_23_to_tile_29_23_0;
	wire vertical_tile_30_23_to_tile_29_23_1;
	wire vertical_tile_30_23_to_tile_29_23_2;
	wire vertical_tile_30_23_to_tile_29_23_3;

	wire vertical_tile_29_24_to_tile_30_24_0;
	wire vertical_tile_29_24_to_tile_30_24_1;
	wire vertical_tile_29_24_to_tile_30_24_2;
	wire vertical_tile_29_24_to_tile_30_24_3;
	wire vertical_tile_30_24_to_tile_29_24_0;
	wire vertical_tile_30_24_to_tile_29_24_1;
	wire vertical_tile_30_24_to_tile_29_24_2;
	wire vertical_tile_30_24_to_tile_29_24_3;

	wire vertical_tile_29_25_to_tile_30_25_0;
	wire vertical_tile_29_25_to_tile_30_25_1;
	wire vertical_tile_29_25_to_tile_30_25_2;
	wire vertical_tile_29_25_to_tile_30_25_3;
	wire vertical_tile_30_25_to_tile_29_25_0;
	wire vertical_tile_30_25_to_tile_29_25_1;
	wire vertical_tile_30_25_to_tile_29_25_2;
	wire vertical_tile_30_25_to_tile_29_25_3;

	wire vertical_tile_29_26_to_tile_30_26_0;
	wire vertical_tile_29_26_to_tile_30_26_1;
	wire vertical_tile_29_26_to_tile_30_26_2;
	wire vertical_tile_29_26_to_tile_30_26_3;
	wire vertical_tile_30_26_to_tile_29_26_0;
	wire vertical_tile_30_26_to_tile_29_26_1;
	wire vertical_tile_30_26_to_tile_29_26_2;
	wire vertical_tile_30_26_to_tile_29_26_3;

	wire vertical_tile_29_27_to_tile_30_27_0;
	wire vertical_tile_29_27_to_tile_30_27_1;
	wire vertical_tile_29_27_to_tile_30_27_2;
	wire vertical_tile_29_27_to_tile_30_27_3;
	wire vertical_tile_30_27_to_tile_29_27_0;
	wire vertical_tile_30_27_to_tile_29_27_1;
	wire vertical_tile_30_27_to_tile_29_27_2;
	wire vertical_tile_30_27_to_tile_29_27_3;

	wire vertical_tile_29_28_to_tile_30_28_0;
	wire vertical_tile_29_28_to_tile_30_28_1;
	wire vertical_tile_29_28_to_tile_30_28_2;
	wire vertical_tile_29_28_to_tile_30_28_3;
	wire vertical_tile_30_28_to_tile_29_28_0;
	wire vertical_tile_30_28_to_tile_29_28_1;
	wire vertical_tile_30_28_to_tile_29_28_2;
	wire vertical_tile_30_28_to_tile_29_28_3;

	wire vertical_tile_29_29_to_tile_30_29_0;
	wire vertical_tile_29_29_to_tile_30_29_1;
	wire vertical_tile_29_29_to_tile_30_29_2;
	wire vertical_tile_29_29_to_tile_30_29_3;
	wire vertical_tile_30_29_to_tile_29_29_0;
	wire vertical_tile_30_29_to_tile_29_29_1;
	wire vertical_tile_30_29_to_tile_29_29_2;
	wire vertical_tile_30_29_to_tile_29_29_3;

	wire vertical_tile_29_30_to_tile_30_30_0;
	wire vertical_tile_29_30_to_tile_30_30_1;
	wire vertical_tile_29_30_to_tile_30_30_2;
	wire vertical_tile_29_30_to_tile_30_30_3;
	wire vertical_tile_30_30_to_tile_29_30_0;
	wire vertical_tile_30_30_to_tile_29_30_1;
	wire vertical_tile_30_30_to_tile_29_30_2;
	wire vertical_tile_30_30_to_tile_29_30_3;

	wire vertical_tile_29_31_to_tile_30_31_0;
	wire vertical_tile_29_31_to_tile_30_31_1;
	wire vertical_tile_29_31_to_tile_30_31_2;
	wire vertical_tile_29_31_to_tile_30_31_3;
	wire vertical_tile_30_31_to_tile_29_31_0;
	wire vertical_tile_30_31_to_tile_29_31_1;
	wire vertical_tile_30_31_to_tile_29_31_2;
	wire vertical_tile_30_31_to_tile_29_31_3;

	wire vertical_tile_30_0_to_tile_31_0_0;
	wire vertical_tile_30_0_to_tile_31_0_1;
	wire vertical_tile_30_0_to_tile_31_0_2;
	wire vertical_tile_30_0_to_tile_31_0_3;
	wire vertical_tile_31_0_to_tile_30_0_0;
	wire vertical_tile_31_0_to_tile_30_0_1;
	wire vertical_tile_31_0_to_tile_30_0_2;
	wire vertical_tile_31_0_to_tile_30_0_3;

	wire vertical_tile_30_1_to_tile_31_1_0;
	wire vertical_tile_30_1_to_tile_31_1_1;
	wire vertical_tile_30_1_to_tile_31_1_2;
	wire vertical_tile_30_1_to_tile_31_1_3;
	wire vertical_tile_31_1_to_tile_30_1_0;
	wire vertical_tile_31_1_to_tile_30_1_1;
	wire vertical_tile_31_1_to_tile_30_1_2;
	wire vertical_tile_31_1_to_tile_30_1_3;

	wire vertical_tile_30_2_to_tile_31_2_0;
	wire vertical_tile_30_2_to_tile_31_2_1;
	wire vertical_tile_30_2_to_tile_31_2_2;
	wire vertical_tile_30_2_to_tile_31_2_3;
	wire vertical_tile_31_2_to_tile_30_2_0;
	wire vertical_tile_31_2_to_tile_30_2_1;
	wire vertical_tile_31_2_to_tile_30_2_2;
	wire vertical_tile_31_2_to_tile_30_2_3;

	wire vertical_tile_30_3_to_tile_31_3_0;
	wire vertical_tile_30_3_to_tile_31_3_1;
	wire vertical_tile_30_3_to_tile_31_3_2;
	wire vertical_tile_30_3_to_tile_31_3_3;
	wire vertical_tile_31_3_to_tile_30_3_0;
	wire vertical_tile_31_3_to_tile_30_3_1;
	wire vertical_tile_31_3_to_tile_30_3_2;
	wire vertical_tile_31_3_to_tile_30_3_3;

	wire vertical_tile_30_4_to_tile_31_4_0;
	wire vertical_tile_30_4_to_tile_31_4_1;
	wire vertical_tile_30_4_to_tile_31_4_2;
	wire vertical_tile_30_4_to_tile_31_4_3;
	wire vertical_tile_31_4_to_tile_30_4_0;
	wire vertical_tile_31_4_to_tile_30_4_1;
	wire vertical_tile_31_4_to_tile_30_4_2;
	wire vertical_tile_31_4_to_tile_30_4_3;

	wire vertical_tile_30_5_to_tile_31_5_0;
	wire vertical_tile_30_5_to_tile_31_5_1;
	wire vertical_tile_30_5_to_tile_31_5_2;
	wire vertical_tile_30_5_to_tile_31_5_3;
	wire vertical_tile_31_5_to_tile_30_5_0;
	wire vertical_tile_31_5_to_tile_30_5_1;
	wire vertical_tile_31_5_to_tile_30_5_2;
	wire vertical_tile_31_5_to_tile_30_5_3;

	wire vertical_tile_30_6_to_tile_31_6_0;
	wire vertical_tile_30_6_to_tile_31_6_1;
	wire vertical_tile_30_6_to_tile_31_6_2;
	wire vertical_tile_30_6_to_tile_31_6_3;
	wire vertical_tile_31_6_to_tile_30_6_0;
	wire vertical_tile_31_6_to_tile_30_6_1;
	wire vertical_tile_31_6_to_tile_30_6_2;
	wire vertical_tile_31_6_to_tile_30_6_3;

	wire vertical_tile_30_7_to_tile_31_7_0;
	wire vertical_tile_30_7_to_tile_31_7_1;
	wire vertical_tile_30_7_to_tile_31_7_2;
	wire vertical_tile_30_7_to_tile_31_7_3;
	wire vertical_tile_31_7_to_tile_30_7_0;
	wire vertical_tile_31_7_to_tile_30_7_1;
	wire vertical_tile_31_7_to_tile_30_7_2;
	wire vertical_tile_31_7_to_tile_30_7_3;

	wire vertical_tile_30_8_to_tile_31_8_0;
	wire vertical_tile_30_8_to_tile_31_8_1;
	wire vertical_tile_30_8_to_tile_31_8_2;
	wire vertical_tile_30_8_to_tile_31_8_3;
	wire vertical_tile_31_8_to_tile_30_8_0;
	wire vertical_tile_31_8_to_tile_30_8_1;
	wire vertical_tile_31_8_to_tile_30_8_2;
	wire vertical_tile_31_8_to_tile_30_8_3;

	wire vertical_tile_30_9_to_tile_31_9_0;
	wire vertical_tile_30_9_to_tile_31_9_1;
	wire vertical_tile_30_9_to_tile_31_9_2;
	wire vertical_tile_30_9_to_tile_31_9_3;
	wire vertical_tile_31_9_to_tile_30_9_0;
	wire vertical_tile_31_9_to_tile_30_9_1;
	wire vertical_tile_31_9_to_tile_30_9_2;
	wire vertical_tile_31_9_to_tile_30_9_3;

	wire vertical_tile_30_10_to_tile_31_10_0;
	wire vertical_tile_30_10_to_tile_31_10_1;
	wire vertical_tile_30_10_to_tile_31_10_2;
	wire vertical_tile_30_10_to_tile_31_10_3;
	wire vertical_tile_31_10_to_tile_30_10_0;
	wire vertical_tile_31_10_to_tile_30_10_1;
	wire vertical_tile_31_10_to_tile_30_10_2;
	wire vertical_tile_31_10_to_tile_30_10_3;

	wire vertical_tile_30_11_to_tile_31_11_0;
	wire vertical_tile_30_11_to_tile_31_11_1;
	wire vertical_tile_30_11_to_tile_31_11_2;
	wire vertical_tile_30_11_to_tile_31_11_3;
	wire vertical_tile_31_11_to_tile_30_11_0;
	wire vertical_tile_31_11_to_tile_30_11_1;
	wire vertical_tile_31_11_to_tile_30_11_2;
	wire vertical_tile_31_11_to_tile_30_11_3;

	wire vertical_tile_30_12_to_tile_31_12_0;
	wire vertical_tile_30_12_to_tile_31_12_1;
	wire vertical_tile_30_12_to_tile_31_12_2;
	wire vertical_tile_30_12_to_tile_31_12_3;
	wire vertical_tile_31_12_to_tile_30_12_0;
	wire vertical_tile_31_12_to_tile_30_12_1;
	wire vertical_tile_31_12_to_tile_30_12_2;
	wire vertical_tile_31_12_to_tile_30_12_3;

	wire vertical_tile_30_13_to_tile_31_13_0;
	wire vertical_tile_30_13_to_tile_31_13_1;
	wire vertical_tile_30_13_to_tile_31_13_2;
	wire vertical_tile_30_13_to_tile_31_13_3;
	wire vertical_tile_31_13_to_tile_30_13_0;
	wire vertical_tile_31_13_to_tile_30_13_1;
	wire vertical_tile_31_13_to_tile_30_13_2;
	wire vertical_tile_31_13_to_tile_30_13_3;

	wire vertical_tile_30_14_to_tile_31_14_0;
	wire vertical_tile_30_14_to_tile_31_14_1;
	wire vertical_tile_30_14_to_tile_31_14_2;
	wire vertical_tile_30_14_to_tile_31_14_3;
	wire vertical_tile_31_14_to_tile_30_14_0;
	wire vertical_tile_31_14_to_tile_30_14_1;
	wire vertical_tile_31_14_to_tile_30_14_2;
	wire vertical_tile_31_14_to_tile_30_14_3;

	wire vertical_tile_30_15_to_tile_31_15_0;
	wire vertical_tile_30_15_to_tile_31_15_1;
	wire vertical_tile_30_15_to_tile_31_15_2;
	wire vertical_tile_30_15_to_tile_31_15_3;
	wire vertical_tile_31_15_to_tile_30_15_0;
	wire vertical_tile_31_15_to_tile_30_15_1;
	wire vertical_tile_31_15_to_tile_30_15_2;
	wire vertical_tile_31_15_to_tile_30_15_3;

	wire vertical_tile_30_16_to_tile_31_16_0;
	wire vertical_tile_30_16_to_tile_31_16_1;
	wire vertical_tile_30_16_to_tile_31_16_2;
	wire vertical_tile_30_16_to_tile_31_16_3;
	wire vertical_tile_31_16_to_tile_30_16_0;
	wire vertical_tile_31_16_to_tile_30_16_1;
	wire vertical_tile_31_16_to_tile_30_16_2;
	wire vertical_tile_31_16_to_tile_30_16_3;

	wire vertical_tile_30_17_to_tile_31_17_0;
	wire vertical_tile_30_17_to_tile_31_17_1;
	wire vertical_tile_30_17_to_tile_31_17_2;
	wire vertical_tile_30_17_to_tile_31_17_3;
	wire vertical_tile_31_17_to_tile_30_17_0;
	wire vertical_tile_31_17_to_tile_30_17_1;
	wire vertical_tile_31_17_to_tile_30_17_2;
	wire vertical_tile_31_17_to_tile_30_17_3;

	wire vertical_tile_30_18_to_tile_31_18_0;
	wire vertical_tile_30_18_to_tile_31_18_1;
	wire vertical_tile_30_18_to_tile_31_18_2;
	wire vertical_tile_30_18_to_tile_31_18_3;
	wire vertical_tile_31_18_to_tile_30_18_0;
	wire vertical_tile_31_18_to_tile_30_18_1;
	wire vertical_tile_31_18_to_tile_30_18_2;
	wire vertical_tile_31_18_to_tile_30_18_3;

	wire vertical_tile_30_19_to_tile_31_19_0;
	wire vertical_tile_30_19_to_tile_31_19_1;
	wire vertical_tile_30_19_to_tile_31_19_2;
	wire vertical_tile_30_19_to_tile_31_19_3;
	wire vertical_tile_31_19_to_tile_30_19_0;
	wire vertical_tile_31_19_to_tile_30_19_1;
	wire vertical_tile_31_19_to_tile_30_19_2;
	wire vertical_tile_31_19_to_tile_30_19_3;

	wire vertical_tile_30_20_to_tile_31_20_0;
	wire vertical_tile_30_20_to_tile_31_20_1;
	wire vertical_tile_30_20_to_tile_31_20_2;
	wire vertical_tile_30_20_to_tile_31_20_3;
	wire vertical_tile_31_20_to_tile_30_20_0;
	wire vertical_tile_31_20_to_tile_30_20_1;
	wire vertical_tile_31_20_to_tile_30_20_2;
	wire vertical_tile_31_20_to_tile_30_20_3;

	wire vertical_tile_30_21_to_tile_31_21_0;
	wire vertical_tile_30_21_to_tile_31_21_1;
	wire vertical_tile_30_21_to_tile_31_21_2;
	wire vertical_tile_30_21_to_tile_31_21_3;
	wire vertical_tile_31_21_to_tile_30_21_0;
	wire vertical_tile_31_21_to_tile_30_21_1;
	wire vertical_tile_31_21_to_tile_30_21_2;
	wire vertical_tile_31_21_to_tile_30_21_3;

	wire vertical_tile_30_22_to_tile_31_22_0;
	wire vertical_tile_30_22_to_tile_31_22_1;
	wire vertical_tile_30_22_to_tile_31_22_2;
	wire vertical_tile_30_22_to_tile_31_22_3;
	wire vertical_tile_31_22_to_tile_30_22_0;
	wire vertical_tile_31_22_to_tile_30_22_1;
	wire vertical_tile_31_22_to_tile_30_22_2;
	wire vertical_tile_31_22_to_tile_30_22_3;

	wire vertical_tile_30_23_to_tile_31_23_0;
	wire vertical_tile_30_23_to_tile_31_23_1;
	wire vertical_tile_30_23_to_tile_31_23_2;
	wire vertical_tile_30_23_to_tile_31_23_3;
	wire vertical_tile_31_23_to_tile_30_23_0;
	wire vertical_tile_31_23_to_tile_30_23_1;
	wire vertical_tile_31_23_to_tile_30_23_2;
	wire vertical_tile_31_23_to_tile_30_23_3;

	wire vertical_tile_30_24_to_tile_31_24_0;
	wire vertical_tile_30_24_to_tile_31_24_1;
	wire vertical_tile_30_24_to_tile_31_24_2;
	wire vertical_tile_30_24_to_tile_31_24_3;
	wire vertical_tile_31_24_to_tile_30_24_0;
	wire vertical_tile_31_24_to_tile_30_24_1;
	wire vertical_tile_31_24_to_tile_30_24_2;
	wire vertical_tile_31_24_to_tile_30_24_3;

	wire vertical_tile_30_25_to_tile_31_25_0;
	wire vertical_tile_30_25_to_tile_31_25_1;
	wire vertical_tile_30_25_to_tile_31_25_2;
	wire vertical_tile_30_25_to_tile_31_25_3;
	wire vertical_tile_31_25_to_tile_30_25_0;
	wire vertical_tile_31_25_to_tile_30_25_1;
	wire vertical_tile_31_25_to_tile_30_25_2;
	wire vertical_tile_31_25_to_tile_30_25_3;

	wire vertical_tile_30_26_to_tile_31_26_0;
	wire vertical_tile_30_26_to_tile_31_26_1;
	wire vertical_tile_30_26_to_tile_31_26_2;
	wire vertical_tile_30_26_to_tile_31_26_3;
	wire vertical_tile_31_26_to_tile_30_26_0;
	wire vertical_tile_31_26_to_tile_30_26_1;
	wire vertical_tile_31_26_to_tile_30_26_2;
	wire vertical_tile_31_26_to_tile_30_26_3;

	wire vertical_tile_30_27_to_tile_31_27_0;
	wire vertical_tile_30_27_to_tile_31_27_1;
	wire vertical_tile_30_27_to_tile_31_27_2;
	wire vertical_tile_30_27_to_tile_31_27_3;
	wire vertical_tile_31_27_to_tile_30_27_0;
	wire vertical_tile_31_27_to_tile_30_27_1;
	wire vertical_tile_31_27_to_tile_30_27_2;
	wire vertical_tile_31_27_to_tile_30_27_3;

	wire vertical_tile_30_28_to_tile_31_28_0;
	wire vertical_tile_30_28_to_tile_31_28_1;
	wire vertical_tile_30_28_to_tile_31_28_2;
	wire vertical_tile_30_28_to_tile_31_28_3;
	wire vertical_tile_31_28_to_tile_30_28_0;
	wire vertical_tile_31_28_to_tile_30_28_1;
	wire vertical_tile_31_28_to_tile_30_28_2;
	wire vertical_tile_31_28_to_tile_30_28_3;

	wire vertical_tile_30_29_to_tile_31_29_0;
	wire vertical_tile_30_29_to_tile_31_29_1;
	wire vertical_tile_30_29_to_tile_31_29_2;
	wire vertical_tile_30_29_to_tile_31_29_3;
	wire vertical_tile_31_29_to_tile_30_29_0;
	wire vertical_tile_31_29_to_tile_30_29_1;
	wire vertical_tile_31_29_to_tile_30_29_2;
	wire vertical_tile_31_29_to_tile_30_29_3;

	wire vertical_tile_30_30_to_tile_31_30_0;
	wire vertical_tile_30_30_to_tile_31_30_1;
	wire vertical_tile_30_30_to_tile_31_30_2;
	wire vertical_tile_30_30_to_tile_31_30_3;
	wire vertical_tile_31_30_to_tile_30_30_0;
	wire vertical_tile_31_30_to_tile_30_30_1;
	wire vertical_tile_31_30_to_tile_30_30_2;
	wire vertical_tile_31_30_to_tile_30_30_3;

	wire vertical_tile_30_31_to_tile_31_31_0;
	wire vertical_tile_30_31_to_tile_31_31_1;
	wire vertical_tile_30_31_to_tile_31_31_2;
	wire vertical_tile_30_31_to_tile_31_31_3;
	wire vertical_tile_31_31_to_tile_30_31_0;
	wire vertical_tile_31_31_to_tile_30_31_1;
	wire vertical_tile_31_31_to_tile_30_31_2;
	wire vertical_tile_31_31_to_tile_30_31_3;

	// Horizontal wires
	wire horizontal_tile_0_0_to_tile_0_1_0;
	wire horizontal_tile_0_0_to_tile_0_1_1;
	wire horizontal_tile_0_0_to_tile_0_1_2;
	wire horizontal_tile_0_0_to_tile_0_1_3;
	wire horizontal_tile_0_1_to_tile_0_0_0;
	wire horizontal_tile_0_1_to_tile_0_0_1;
	wire horizontal_tile_0_1_to_tile_0_0_2;
	wire horizontal_tile_0_1_to_tile_0_0_3;

	wire horizontal_tile_1_0_to_tile_1_1_0;
	wire horizontal_tile_1_0_to_tile_1_1_1;
	wire horizontal_tile_1_0_to_tile_1_1_2;
	wire horizontal_tile_1_0_to_tile_1_1_3;
	wire horizontal_tile_1_1_to_tile_1_0_0;
	wire horizontal_tile_1_1_to_tile_1_0_1;
	wire horizontal_tile_1_1_to_tile_1_0_2;
	wire horizontal_tile_1_1_to_tile_1_0_3;

	wire horizontal_tile_2_0_to_tile_2_1_0;
	wire horizontal_tile_2_0_to_tile_2_1_1;
	wire horizontal_tile_2_0_to_tile_2_1_2;
	wire horizontal_tile_2_0_to_tile_2_1_3;
	wire horizontal_tile_2_1_to_tile_2_0_0;
	wire horizontal_tile_2_1_to_tile_2_0_1;
	wire horizontal_tile_2_1_to_tile_2_0_2;
	wire horizontal_tile_2_1_to_tile_2_0_3;

	wire horizontal_tile_3_0_to_tile_3_1_0;
	wire horizontal_tile_3_0_to_tile_3_1_1;
	wire horizontal_tile_3_0_to_tile_3_1_2;
	wire horizontal_tile_3_0_to_tile_3_1_3;
	wire horizontal_tile_3_1_to_tile_3_0_0;
	wire horizontal_tile_3_1_to_tile_3_0_1;
	wire horizontal_tile_3_1_to_tile_3_0_2;
	wire horizontal_tile_3_1_to_tile_3_0_3;

	wire horizontal_tile_4_0_to_tile_4_1_0;
	wire horizontal_tile_4_0_to_tile_4_1_1;
	wire horizontal_tile_4_0_to_tile_4_1_2;
	wire horizontal_tile_4_0_to_tile_4_1_3;
	wire horizontal_tile_4_1_to_tile_4_0_0;
	wire horizontal_tile_4_1_to_tile_4_0_1;
	wire horizontal_tile_4_1_to_tile_4_0_2;
	wire horizontal_tile_4_1_to_tile_4_0_3;

	wire horizontal_tile_5_0_to_tile_5_1_0;
	wire horizontal_tile_5_0_to_tile_5_1_1;
	wire horizontal_tile_5_0_to_tile_5_1_2;
	wire horizontal_tile_5_0_to_tile_5_1_3;
	wire horizontal_tile_5_1_to_tile_5_0_0;
	wire horizontal_tile_5_1_to_tile_5_0_1;
	wire horizontal_tile_5_1_to_tile_5_0_2;
	wire horizontal_tile_5_1_to_tile_5_0_3;

	wire horizontal_tile_6_0_to_tile_6_1_0;
	wire horizontal_tile_6_0_to_tile_6_1_1;
	wire horizontal_tile_6_0_to_tile_6_1_2;
	wire horizontal_tile_6_0_to_tile_6_1_3;
	wire horizontal_tile_6_1_to_tile_6_0_0;
	wire horizontal_tile_6_1_to_tile_6_0_1;
	wire horizontal_tile_6_1_to_tile_6_0_2;
	wire horizontal_tile_6_1_to_tile_6_0_3;

	wire horizontal_tile_7_0_to_tile_7_1_0;
	wire horizontal_tile_7_0_to_tile_7_1_1;
	wire horizontal_tile_7_0_to_tile_7_1_2;
	wire horizontal_tile_7_0_to_tile_7_1_3;
	wire horizontal_tile_7_1_to_tile_7_0_0;
	wire horizontal_tile_7_1_to_tile_7_0_1;
	wire horizontal_tile_7_1_to_tile_7_0_2;
	wire horizontal_tile_7_1_to_tile_7_0_3;

	wire horizontal_tile_8_0_to_tile_8_1_0;
	wire horizontal_tile_8_0_to_tile_8_1_1;
	wire horizontal_tile_8_0_to_tile_8_1_2;
	wire horizontal_tile_8_0_to_tile_8_1_3;
	wire horizontal_tile_8_1_to_tile_8_0_0;
	wire horizontal_tile_8_1_to_tile_8_0_1;
	wire horizontal_tile_8_1_to_tile_8_0_2;
	wire horizontal_tile_8_1_to_tile_8_0_3;

	wire horizontal_tile_9_0_to_tile_9_1_0;
	wire horizontal_tile_9_0_to_tile_9_1_1;
	wire horizontal_tile_9_0_to_tile_9_1_2;
	wire horizontal_tile_9_0_to_tile_9_1_3;
	wire horizontal_tile_9_1_to_tile_9_0_0;
	wire horizontal_tile_9_1_to_tile_9_0_1;
	wire horizontal_tile_9_1_to_tile_9_0_2;
	wire horizontal_tile_9_1_to_tile_9_0_3;

	wire horizontal_tile_10_0_to_tile_10_1_0;
	wire horizontal_tile_10_0_to_tile_10_1_1;
	wire horizontal_tile_10_0_to_tile_10_1_2;
	wire horizontal_tile_10_0_to_tile_10_1_3;
	wire horizontal_tile_10_1_to_tile_10_0_0;
	wire horizontal_tile_10_1_to_tile_10_0_1;
	wire horizontal_tile_10_1_to_tile_10_0_2;
	wire horizontal_tile_10_1_to_tile_10_0_3;

	wire horizontal_tile_11_0_to_tile_11_1_0;
	wire horizontal_tile_11_0_to_tile_11_1_1;
	wire horizontal_tile_11_0_to_tile_11_1_2;
	wire horizontal_tile_11_0_to_tile_11_1_3;
	wire horizontal_tile_11_1_to_tile_11_0_0;
	wire horizontal_tile_11_1_to_tile_11_0_1;
	wire horizontal_tile_11_1_to_tile_11_0_2;
	wire horizontal_tile_11_1_to_tile_11_0_3;

	wire horizontal_tile_12_0_to_tile_12_1_0;
	wire horizontal_tile_12_0_to_tile_12_1_1;
	wire horizontal_tile_12_0_to_tile_12_1_2;
	wire horizontal_tile_12_0_to_tile_12_1_3;
	wire horizontal_tile_12_1_to_tile_12_0_0;
	wire horizontal_tile_12_1_to_tile_12_0_1;
	wire horizontal_tile_12_1_to_tile_12_0_2;
	wire horizontal_tile_12_1_to_tile_12_0_3;

	wire horizontal_tile_13_0_to_tile_13_1_0;
	wire horizontal_tile_13_0_to_tile_13_1_1;
	wire horizontal_tile_13_0_to_tile_13_1_2;
	wire horizontal_tile_13_0_to_tile_13_1_3;
	wire horizontal_tile_13_1_to_tile_13_0_0;
	wire horizontal_tile_13_1_to_tile_13_0_1;
	wire horizontal_tile_13_1_to_tile_13_0_2;
	wire horizontal_tile_13_1_to_tile_13_0_3;

	wire horizontal_tile_14_0_to_tile_14_1_0;
	wire horizontal_tile_14_0_to_tile_14_1_1;
	wire horizontal_tile_14_0_to_tile_14_1_2;
	wire horizontal_tile_14_0_to_tile_14_1_3;
	wire horizontal_tile_14_1_to_tile_14_0_0;
	wire horizontal_tile_14_1_to_tile_14_0_1;
	wire horizontal_tile_14_1_to_tile_14_0_2;
	wire horizontal_tile_14_1_to_tile_14_0_3;

	wire horizontal_tile_15_0_to_tile_15_1_0;
	wire horizontal_tile_15_0_to_tile_15_1_1;
	wire horizontal_tile_15_0_to_tile_15_1_2;
	wire horizontal_tile_15_0_to_tile_15_1_3;
	wire horizontal_tile_15_1_to_tile_15_0_0;
	wire horizontal_tile_15_1_to_tile_15_0_1;
	wire horizontal_tile_15_1_to_tile_15_0_2;
	wire horizontal_tile_15_1_to_tile_15_0_3;

	wire horizontal_tile_16_0_to_tile_16_1_0;
	wire horizontal_tile_16_0_to_tile_16_1_1;
	wire horizontal_tile_16_0_to_tile_16_1_2;
	wire horizontal_tile_16_0_to_tile_16_1_3;
	wire horizontal_tile_16_1_to_tile_16_0_0;
	wire horizontal_tile_16_1_to_tile_16_0_1;
	wire horizontal_tile_16_1_to_tile_16_0_2;
	wire horizontal_tile_16_1_to_tile_16_0_3;

	wire horizontal_tile_17_0_to_tile_17_1_0;
	wire horizontal_tile_17_0_to_tile_17_1_1;
	wire horizontal_tile_17_0_to_tile_17_1_2;
	wire horizontal_tile_17_0_to_tile_17_1_3;
	wire horizontal_tile_17_1_to_tile_17_0_0;
	wire horizontal_tile_17_1_to_tile_17_0_1;
	wire horizontal_tile_17_1_to_tile_17_0_2;
	wire horizontal_tile_17_1_to_tile_17_0_3;

	wire horizontal_tile_18_0_to_tile_18_1_0;
	wire horizontal_tile_18_0_to_tile_18_1_1;
	wire horizontal_tile_18_0_to_tile_18_1_2;
	wire horizontal_tile_18_0_to_tile_18_1_3;
	wire horizontal_tile_18_1_to_tile_18_0_0;
	wire horizontal_tile_18_1_to_tile_18_0_1;
	wire horizontal_tile_18_1_to_tile_18_0_2;
	wire horizontal_tile_18_1_to_tile_18_0_3;

	wire horizontal_tile_19_0_to_tile_19_1_0;
	wire horizontal_tile_19_0_to_tile_19_1_1;
	wire horizontal_tile_19_0_to_tile_19_1_2;
	wire horizontal_tile_19_0_to_tile_19_1_3;
	wire horizontal_tile_19_1_to_tile_19_0_0;
	wire horizontal_tile_19_1_to_tile_19_0_1;
	wire horizontal_tile_19_1_to_tile_19_0_2;
	wire horizontal_tile_19_1_to_tile_19_0_3;

	wire horizontal_tile_20_0_to_tile_20_1_0;
	wire horizontal_tile_20_0_to_tile_20_1_1;
	wire horizontal_tile_20_0_to_tile_20_1_2;
	wire horizontal_tile_20_0_to_tile_20_1_3;
	wire horizontal_tile_20_1_to_tile_20_0_0;
	wire horizontal_tile_20_1_to_tile_20_0_1;
	wire horizontal_tile_20_1_to_tile_20_0_2;
	wire horizontal_tile_20_1_to_tile_20_0_3;

	wire horizontal_tile_21_0_to_tile_21_1_0;
	wire horizontal_tile_21_0_to_tile_21_1_1;
	wire horizontal_tile_21_0_to_tile_21_1_2;
	wire horizontal_tile_21_0_to_tile_21_1_3;
	wire horizontal_tile_21_1_to_tile_21_0_0;
	wire horizontal_tile_21_1_to_tile_21_0_1;
	wire horizontal_tile_21_1_to_tile_21_0_2;
	wire horizontal_tile_21_1_to_tile_21_0_3;

	wire horizontal_tile_22_0_to_tile_22_1_0;
	wire horizontal_tile_22_0_to_tile_22_1_1;
	wire horizontal_tile_22_0_to_tile_22_1_2;
	wire horizontal_tile_22_0_to_tile_22_1_3;
	wire horizontal_tile_22_1_to_tile_22_0_0;
	wire horizontal_tile_22_1_to_tile_22_0_1;
	wire horizontal_tile_22_1_to_tile_22_0_2;
	wire horizontal_tile_22_1_to_tile_22_0_3;

	wire horizontal_tile_23_0_to_tile_23_1_0;
	wire horizontal_tile_23_0_to_tile_23_1_1;
	wire horizontal_tile_23_0_to_tile_23_1_2;
	wire horizontal_tile_23_0_to_tile_23_1_3;
	wire horizontal_tile_23_1_to_tile_23_0_0;
	wire horizontal_tile_23_1_to_tile_23_0_1;
	wire horizontal_tile_23_1_to_tile_23_0_2;
	wire horizontal_tile_23_1_to_tile_23_0_3;

	wire horizontal_tile_24_0_to_tile_24_1_0;
	wire horizontal_tile_24_0_to_tile_24_1_1;
	wire horizontal_tile_24_0_to_tile_24_1_2;
	wire horizontal_tile_24_0_to_tile_24_1_3;
	wire horizontal_tile_24_1_to_tile_24_0_0;
	wire horizontal_tile_24_1_to_tile_24_0_1;
	wire horizontal_tile_24_1_to_tile_24_0_2;
	wire horizontal_tile_24_1_to_tile_24_0_3;

	wire horizontal_tile_25_0_to_tile_25_1_0;
	wire horizontal_tile_25_0_to_tile_25_1_1;
	wire horizontal_tile_25_0_to_tile_25_1_2;
	wire horizontal_tile_25_0_to_tile_25_1_3;
	wire horizontal_tile_25_1_to_tile_25_0_0;
	wire horizontal_tile_25_1_to_tile_25_0_1;
	wire horizontal_tile_25_1_to_tile_25_0_2;
	wire horizontal_tile_25_1_to_tile_25_0_3;

	wire horizontal_tile_26_0_to_tile_26_1_0;
	wire horizontal_tile_26_0_to_tile_26_1_1;
	wire horizontal_tile_26_0_to_tile_26_1_2;
	wire horizontal_tile_26_0_to_tile_26_1_3;
	wire horizontal_tile_26_1_to_tile_26_0_0;
	wire horizontal_tile_26_1_to_tile_26_0_1;
	wire horizontal_tile_26_1_to_tile_26_0_2;
	wire horizontal_tile_26_1_to_tile_26_0_3;

	wire horizontal_tile_27_0_to_tile_27_1_0;
	wire horizontal_tile_27_0_to_tile_27_1_1;
	wire horizontal_tile_27_0_to_tile_27_1_2;
	wire horizontal_tile_27_0_to_tile_27_1_3;
	wire horizontal_tile_27_1_to_tile_27_0_0;
	wire horizontal_tile_27_1_to_tile_27_0_1;
	wire horizontal_tile_27_1_to_tile_27_0_2;
	wire horizontal_tile_27_1_to_tile_27_0_3;

	wire horizontal_tile_28_0_to_tile_28_1_0;
	wire horizontal_tile_28_0_to_tile_28_1_1;
	wire horizontal_tile_28_0_to_tile_28_1_2;
	wire horizontal_tile_28_0_to_tile_28_1_3;
	wire horizontal_tile_28_1_to_tile_28_0_0;
	wire horizontal_tile_28_1_to_tile_28_0_1;
	wire horizontal_tile_28_1_to_tile_28_0_2;
	wire horizontal_tile_28_1_to_tile_28_0_3;

	wire horizontal_tile_29_0_to_tile_29_1_0;
	wire horizontal_tile_29_0_to_tile_29_1_1;
	wire horizontal_tile_29_0_to_tile_29_1_2;
	wire horizontal_tile_29_0_to_tile_29_1_3;
	wire horizontal_tile_29_1_to_tile_29_0_0;
	wire horizontal_tile_29_1_to_tile_29_0_1;
	wire horizontal_tile_29_1_to_tile_29_0_2;
	wire horizontal_tile_29_1_to_tile_29_0_3;

	wire horizontal_tile_30_0_to_tile_30_1_0;
	wire horizontal_tile_30_0_to_tile_30_1_1;
	wire horizontal_tile_30_0_to_tile_30_1_2;
	wire horizontal_tile_30_0_to_tile_30_1_3;
	wire horizontal_tile_30_1_to_tile_30_0_0;
	wire horizontal_tile_30_1_to_tile_30_0_1;
	wire horizontal_tile_30_1_to_tile_30_0_2;
	wire horizontal_tile_30_1_to_tile_30_0_3;

	wire horizontal_tile_31_0_to_tile_31_1_0;
	wire horizontal_tile_31_0_to_tile_31_1_1;
	wire horizontal_tile_31_0_to_tile_31_1_2;
	wire horizontal_tile_31_0_to_tile_31_1_3;
	wire horizontal_tile_31_1_to_tile_31_0_0;
	wire horizontal_tile_31_1_to_tile_31_0_1;
	wire horizontal_tile_31_1_to_tile_31_0_2;
	wire horizontal_tile_31_1_to_tile_31_0_3;

	wire horizontal_tile_0_1_to_tile_0_2_0;
	wire horizontal_tile_0_1_to_tile_0_2_1;
	wire horizontal_tile_0_1_to_tile_0_2_2;
	wire horizontal_tile_0_1_to_tile_0_2_3;
	wire horizontal_tile_0_2_to_tile_0_1_0;
	wire horizontal_tile_0_2_to_tile_0_1_1;
	wire horizontal_tile_0_2_to_tile_0_1_2;
	wire horizontal_tile_0_2_to_tile_0_1_3;

	wire horizontal_tile_1_1_to_tile_1_2_0;
	wire horizontal_tile_1_1_to_tile_1_2_1;
	wire horizontal_tile_1_1_to_tile_1_2_2;
	wire horizontal_tile_1_1_to_tile_1_2_3;
	wire horizontal_tile_1_2_to_tile_1_1_0;
	wire horizontal_tile_1_2_to_tile_1_1_1;
	wire horizontal_tile_1_2_to_tile_1_1_2;
	wire horizontal_tile_1_2_to_tile_1_1_3;

	wire horizontal_tile_2_1_to_tile_2_2_0;
	wire horizontal_tile_2_1_to_tile_2_2_1;
	wire horizontal_tile_2_1_to_tile_2_2_2;
	wire horizontal_tile_2_1_to_tile_2_2_3;
	wire horizontal_tile_2_2_to_tile_2_1_0;
	wire horizontal_tile_2_2_to_tile_2_1_1;
	wire horizontal_tile_2_2_to_tile_2_1_2;
	wire horizontal_tile_2_2_to_tile_2_1_3;

	wire horizontal_tile_3_1_to_tile_3_2_0;
	wire horizontal_tile_3_1_to_tile_3_2_1;
	wire horizontal_tile_3_1_to_tile_3_2_2;
	wire horizontal_tile_3_1_to_tile_3_2_3;
	wire horizontal_tile_3_2_to_tile_3_1_0;
	wire horizontal_tile_3_2_to_tile_3_1_1;
	wire horizontal_tile_3_2_to_tile_3_1_2;
	wire horizontal_tile_3_2_to_tile_3_1_3;

	wire horizontal_tile_4_1_to_tile_4_2_0;
	wire horizontal_tile_4_1_to_tile_4_2_1;
	wire horizontal_tile_4_1_to_tile_4_2_2;
	wire horizontal_tile_4_1_to_tile_4_2_3;
	wire horizontal_tile_4_2_to_tile_4_1_0;
	wire horizontal_tile_4_2_to_tile_4_1_1;
	wire horizontal_tile_4_2_to_tile_4_1_2;
	wire horizontal_tile_4_2_to_tile_4_1_3;

	wire horizontal_tile_5_1_to_tile_5_2_0;
	wire horizontal_tile_5_1_to_tile_5_2_1;
	wire horizontal_tile_5_1_to_tile_5_2_2;
	wire horizontal_tile_5_1_to_tile_5_2_3;
	wire horizontal_tile_5_2_to_tile_5_1_0;
	wire horizontal_tile_5_2_to_tile_5_1_1;
	wire horizontal_tile_5_2_to_tile_5_1_2;
	wire horizontal_tile_5_2_to_tile_5_1_3;

	wire horizontal_tile_6_1_to_tile_6_2_0;
	wire horizontal_tile_6_1_to_tile_6_2_1;
	wire horizontal_tile_6_1_to_tile_6_2_2;
	wire horizontal_tile_6_1_to_tile_6_2_3;
	wire horizontal_tile_6_2_to_tile_6_1_0;
	wire horizontal_tile_6_2_to_tile_6_1_1;
	wire horizontal_tile_6_2_to_tile_6_1_2;
	wire horizontal_tile_6_2_to_tile_6_1_3;

	wire horizontal_tile_7_1_to_tile_7_2_0;
	wire horizontal_tile_7_1_to_tile_7_2_1;
	wire horizontal_tile_7_1_to_tile_7_2_2;
	wire horizontal_tile_7_1_to_tile_7_2_3;
	wire horizontal_tile_7_2_to_tile_7_1_0;
	wire horizontal_tile_7_2_to_tile_7_1_1;
	wire horizontal_tile_7_2_to_tile_7_1_2;
	wire horizontal_tile_7_2_to_tile_7_1_3;

	wire horizontal_tile_8_1_to_tile_8_2_0;
	wire horizontal_tile_8_1_to_tile_8_2_1;
	wire horizontal_tile_8_1_to_tile_8_2_2;
	wire horizontal_tile_8_1_to_tile_8_2_3;
	wire horizontal_tile_8_2_to_tile_8_1_0;
	wire horizontal_tile_8_2_to_tile_8_1_1;
	wire horizontal_tile_8_2_to_tile_8_1_2;
	wire horizontal_tile_8_2_to_tile_8_1_3;

	wire horizontal_tile_9_1_to_tile_9_2_0;
	wire horizontal_tile_9_1_to_tile_9_2_1;
	wire horizontal_tile_9_1_to_tile_9_2_2;
	wire horizontal_tile_9_1_to_tile_9_2_3;
	wire horizontal_tile_9_2_to_tile_9_1_0;
	wire horizontal_tile_9_2_to_tile_9_1_1;
	wire horizontal_tile_9_2_to_tile_9_1_2;
	wire horizontal_tile_9_2_to_tile_9_1_3;

	wire horizontal_tile_10_1_to_tile_10_2_0;
	wire horizontal_tile_10_1_to_tile_10_2_1;
	wire horizontal_tile_10_1_to_tile_10_2_2;
	wire horizontal_tile_10_1_to_tile_10_2_3;
	wire horizontal_tile_10_2_to_tile_10_1_0;
	wire horizontal_tile_10_2_to_tile_10_1_1;
	wire horizontal_tile_10_2_to_tile_10_1_2;
	wire horizontal_tile_10_2_to_tile_10_1_3;

	wire horizontal_tile_11_1_to_tile_11_2_0;
	wire horizontal_tile_11_1_to_tile_11_2_1;
	wire horizontal_tile_11_1_to_tile_11_2_2;
	wire horizontal_tile_11_1_to_tile_11_2_3;
	wire horizontal_tile_11_2_to_tile_11_1_0;
	wire horizontal_tile_11_2_to_tile_11_1_1;
	wire horizontal_tile_11_2_to_tile_11_1_2;
	wire horizontal_tile_11_2_to_tile_11_1_3;

	wire horizontal_tile_12_1_to_tile_12_2_0;
	wire horizontal_tile_12_1_to_tile_12_2_1;
	wire horizontal_tile_12_1_to_tile_12_2_2;
	wire horizontal_tile_12_1_to_tile_12_2_3;
	wire horizontal_tile_12_2_to_tile_12_1_0;
	wire horizontal_tile_12_2_to_tile_12_1_1;
	wire horizontal_tile_12_2_to_tile_12_1_2;
	wire horizontal_tile_12_2_to_tile_12_1_3;

	wire horizontal_tile_13_1_to_tile_13_2_0;
	wire horizontal_tile_13_1_to_tile_13_2_1;
	wire horizontal_tile_13_1_to_tile_13_2_2;
	wire horizontal_tile_13_1_to_tile_13_2_3;
	wire horizontal_tile_13_2_to_tile_13_1_0;
	wire horizontal_tile_13_2_to_tile_13_1_1;
	wire horizontal_tile_13_2_to_tile_13_1_2;
	wire horizontal_tile_13_2_to_tile_13_1_3;

	wire horizontal_tile_14_1_to_tile_14_2_0;
	wire horizontal_tile_14_1_to_tile_14_2_1;
	wire horizontal_tile_14_1_to_tile_14_2_2;
	wire horizontal_tile_14_1_to_tile_14_2_3;
	wire horizontal_tile_14_2_to_tile_14_1_0;
	wire horizontal_tile_14_2_to_tile_14_1_1;
	wire horizontal_tile_14_2_to_tile_14_1_2;
	wire horizontal_tile_14_2_to_tile_14_1_3;

	wire horizontal_tile_15_1_to_tile_15_2_0;
	wire horizontal_tile_15_1_to_tile_15_2_1;
	wire horizontal_tile_15_1_to_tile_15_2_2;
	wire horizontal_tile_15_1_to_tile_15_2_3;
	wire horizontal_tile_15_2_to_tile_15_1_0;
	wire horizontal_tile_15_2_to_tile_15_1_1;
	wire horizontal_tile_15_2_to_tile_15_1_2;
	wire horizontal_tile_15_2_to_tile_15_1_3;

	wire horizontal_tile_16_1_to_tile_16_2_0;
	wire horizontal_tile_16_1_to_tile_16_2_1;
	wire horizontal_tile_16_1_to_tile_16_2_2;
	wire horizontal_tile_16_1_to_tile_16_2_3;
	wire horizontal_tile_16_2_to_tile_16_1_0;
	wire horizontal_tile_16_2_to_tile_16_1_1;
	wire horizontal_tile_16_2_to_tile_16_1_2;
	wire horizontal_tile_16_2_to_tile_16_1_3;

	wire horizontal_tile_17_1_to_tile_17_2_0;
	wire horizontal_tile_17_1_to_tile_17_2_1;
	wire horizontal_tile_17_1_to_tile_17_2_2;
	wire horizontal_tile_17_1_to_tile_17_2_3;
	wire horizontal_tile_17_2_to_tile_17_1_0;
	wire horizontal_tile_17_2_to_tile_17_1_1;
	wire horizontal_tile_17_2_to_tile_17_1_2;
	wire horizontal_tile_17_2_to_tile_17_1_3;

	wire horizontal_tile_18_1_to_tile_18_2_0;
	wire horizontal_tile_18_1_to_tile_18_2_1;
	wire horizontal_tile_18_1_to_tile_18_2_2;
	wire horizontal_tile_18_1_to_tile_18_2_3;
	wire horizontal_tile_18_2_to_tile_18_1_0;
	wire horizontal_tile_18_2_to_tile_18_1_1;
	wire horizontal_tile_18_2_to_tile_18_1_2;
	wire horizontal_tile_18_2_to_tile_18_1_3;

	wire horizontal_tile_19_1_to_tile_19_2_0;
	wire horizontal_tile_19_1_to_tile_19_2_1;
	wire horizontal_tile_19_1_to_tile_19_2_2;
	wire horizontal_tile_19_1_to_tile_19_2_3;
	wire horizontal_tile_19_2_to_tile_19_1_0;
	wire horizontal_tile_19_2_to_tile_19_1_1;
	wire horizontal_tile_19_2_to_tile_19_1_2;
	wire horizontal_tile_19_2_to_tile_19_1_3;

	wire horizontal_tile_20_1_to_tile_20_2_0;
	wire horizontal_tile_20_1_to_tile_20_2_1;
	wire horizontal_tile_20_1_to_tile_20_2_2;
	wire horizontal_tile_20_1_to_tile_20_2_3;
	wire horizontal_tile_20_2_to_tile_20_1_0;
	wire horizontal_tile_20_2_to_tile_20_1_1;
	wire horizontal_tile_20_2_to_tile_20_1_2;
	wire horizontal_tile_20_2_to_tile_20_1_3;

	wire horizontal_tile_21_1_to_tile_21_2_0;
	wire horizontal_tile_21_1_to_tile_21_2_1;
	wire horizontal_tile_21_1_to_tile_21_2_2;
	wire horizontal_tile_21_1_to_tile_21_2_3;
	wire horizontal_tile_21_2_to_tile_21_1_0;
	wire horizontal_tile_21_2_to_tile_21_1_1;
	wire horizontal_tile_21_2_to_tile_21_1_2;
	wire horizontal_tile_21_2_to_tile_21_1_3;

	wire horizontal_tile_22_1_to_tile_22_2_0;
	wire horizontal_tile_22_1_to_tile_22_2_1;
	wire horizontal_tile_22_1_to_tile_22_2_2;
	wire horizontal_tile_22_1_to_tile_22_2_3;
	wire horizontal_tile_22_2_to_tile_22_1_0;
	wire horizontal_tile_22_2_to_tile_22_1_1;
	wire horizontal_tile_22_2_to_tile_22_1_2;
	wire horizontal_tile_22_2_to_tile_22_1_3;

	wire horizontal_tile_23_1_to_tile_23_2_0;
	wire horizontal_tile_23_1_to_tile_23_2_1;
	wire horizontal_tile_23_1_to_tile_23_2_2;
	wire horizontal_tile_23_1_to_tile_23_2_3;
	wire horizontal_tile_23_2_to_tile_23_1_0;
	wire horizontal_tile_23_2_to_tile_23_1_1;
	wire horizontal_tile_23_2_to_tile_23_1_2;
	wire horizontal_tile_23_2_to_tile_23_1_3;

	wire horizontal_tile_24_1_to_tile_24_2_0;
	wire horizontal_tile_24_1_to_tile_24_2_1;
	wire horizontal_tile_24_1_to_tile_24_2_2;
	wire horizontal_tile_24_1_to_tile_24_2_3;
	wire horizontal_tile_24_2_to_tile_24_1_0;
	wire horizontal_tile_24_2_to_tile_24_1_1;
	wire horizontal_tile_24_2_to_tile_24_1_2;
	wire horizontal_tile_24_2_to_tile_24_1_3;

	wire horizontal_tile_25_1_to_tile_25_2_0;
	wire horizontal_tile_25_1_to_tile_25_2_1;
	wire horizontal_tile_25_1_to_tile_25_2_2;
	wire horizontal_tile_25_1_to_tile_25_2_3;
	wire horizontal_tile_25_2_to_tile_25_1_0;
	wire horizontal_tile_25_2_to_tile_25_1_1;
	wire horizontal_tile_25_2_to_tile_25_1_2;
	wire horizontal_tile_25_2_to_tile_25_1_3;

	wire horizontal_tile_26_1_to_tile_26_2_0;
	wire horizontal_tile_26_1_to_tile_26_2_1;
	wire horizontal_tile_26_1_to_tile_26_2_2;
	wire horizontal_tile_26_1_to_tile_26_2_3;
	wire horizontal_tile_26_2_to_tile_26_1_0;
	wire horizontal_tile_26_2_to_tile_26_1_1;
	wire horizontal_tile_26_2_to_tile_26_1_2;
	wire horizontal_tile_26_2_to_tile_26_1_3;

	wire horizontal_tile_27_1_to_tile_27_2_0;
	wire horizontal_tile_27_1_to_tile_27_2_1;
	wire horizontal_tile_27_1_to_tile_27_2_2;
	wire horizontal_tile_27_1_to_tile_27_2_3;
	wire horizontal_tile_27_2_to_tile_27_1_0;
	wire horizontal_tile_27_2_to_tile_27_1_1;
	wire horizontal_tile_27_2_to_tile_27_1_2;
	wire horizontal_tile_27_2_to_tile_27_1_3;

	wire horizontal_tile_28_1_to_tile_28_2_0;
	wire horizontal_tile_28_1_to_tile_28_2_1;
	wire horizontal_tile_28_1_to_tile_28_2_2;
	wire horizontal_tile_28_1_to_tile_28_2_3;
	wire horizontal_tile_28_2_to_tile_28_1_0;
	wire horizontal_tile_28_2_to_tile_28_1_1;
	wire horizontal_tile_28_2_to_tile_28_1_2;
	wire horizontal_tile_28_2_to_tile_28_1_3;

	wire horizontal_tile_29_1_to_tile_29_2_0;
	wire horizontal_tile_29_1_to_tile_29_2_1;
	wire horizontal_tile_29_1_to_tile_29_2_2;
	wire horizontal_tile_29_1_to_tile_29_2_3;
	wire horizontal_tile_29_2_to_tile_29_1_0;
	wire horizontal_tile_29_2_to_tile_29_1_1;
	wire horizontal_tile_29_2_to_tile_29_1_2;
	wire horizontal_tile_29_2_to_tile_29_1_3;

	wire horizontal_tile_30_1_to_tile_30_2_0;
	wire horizontal_tile_30_1_to_tile_30_2_1;
	wire horizontal_tile_30_1_to_tile_30_2_2;
	wire horizontal_tile_30_1_to_tile_30_2_3;
	wire horizontal_tile_30_2_to_tile_30_1_0;
	wire horizontal_tile_30_2_to_tile_30_1_1;
	wire horizontal_tile_30_2_to_tile_30_1_2;
	wire horizontal_tile_30_2_to_tile_30_1_3;

	wire horizontal_tile_31_1_to_tile_31_2_0;
	wire horizontal_tile_31_1_to_tile_31_2_1;
	wire horizontal_tile_31_1_to_tile_31_2_2;
	wire horizontal_tile_31_1_to_tile_31_2_3;
	wire horizontal_tile_31_2_to_tile_31_1_0;
	wire horizontal_tile_31_2_to_tile_31_1_1;
	wire horizontal_tile_31_2_to_tile_31_1_2;
	wire horizontal_tile_31_2_to_tile_31_1_3;

	wire horizontal_tile_0_2_to_tile_0_3_0;
	wire horizontal_tile_0_2_to_tile_0_3_1;
	wire horizontal_tile_0_2_to_tile_0_3_2;
	wire horizontal_tile_0_2_to_tile_0_3_3;
	wire horizontal_tile_0_3_to_tile_0_2_0;
	wire horizontal_tile_0_3_to_tile_0_2_1;
	wire horizontal_tile_0_3_to_tile_0_2_2;
	wire horizontal_tile_0_3_to_tile_0_2_3;

	wire horizontal_tile_1_2_to_tile_1_3_0;
	wire horizontal_tile_1_2_to_tile_1_3_1;
	wire horizontal_tile_1_2_to_tile_1_3_2;
	wire horizontal_tile_1_2_to_tile_1_3_3;
	wire horizontal_tile_1_3_to_tile_1_2_0;
	wire horizontal_tile_1_3_to_tile_1_2_1;
	wire horizontal_tile_1_3_to_tile_1_2_2;
	wire horizontal_tile_1_3_to_tile_1_2_3;

	wire horizontal_tile_2_2_to_tile_2_3_0;
	wire horizontal_tile_2_2_to_tile_2_3_1;
	wire horizontal_tile_2_2_to_tile_2_3_2;
	wire horizontal_tile_2_2_to_tile_2_3_3;
	wire horizontal_tile_2_3_to_tile_2_2_0;
	wire horizontal_tile_2_3_to_tile_2_2_1;
	wire horizontal_tile_2_3_to_tile_2_2_2;
	wire horizontal_tile_2_3_to_tile_2_2_3;

	wire horizontal_tile_3_2_to_tile_3_3_0;
	wire horizontal_tile_3_2_to_tile_3_3_1;
	wire horizontal_tile_3_2_to_tile_3_3_2;
	wire horizontal_tile_3_2_to_tile_3_3_3;
	wire horizontal_tile_3_3_to_tile_3_2_0;
	wire horizontal_tile_3_3_to_tile_3_2_1;
	wire horizontal_tile_3_3_to_tile_3_2_2;
	wire horizontal_tile_3_3_to_tile_3_2_3;

	wire horizontal_tile_4_2_to_tile_4_3_0;
	wire horizontal_tile_4_2_to_tile_4_3_1;
	wire horizontal_tile_4_2_to_tile_4_3_2;
	wire horizontal_tile_4_2_to_tile_4_3_3;
	wire horizontal_tile_4_3_to_tile_4_2_0;
	wire horizontal_tile_4_3_to_tile_4_2_1;
	wire horizontal_tile_4_3_to_tile_4_2_2;
	wire horizontal_tile_4_3_to_tile_4_2_3;

	wire horizontal_tile_5_2_to_tile_5_3_0;
	wire horizontal_tile_5_2_to_tile_5_3_1;
	wire horizontal_tile_5_2_to_tile_5_3_2;
	wire horizontal_tile_5_2_to_tile_5_3_3;
	wire horizontal_tile_5_3_to_tile_5_2_0;
	wire horizontal_tile_5_3_to_tile_5_2_1;
	wire horizontal_tile_5_3_to_tile_5_2_2;
	wire horizontal_tile_5_3_to_tile_5_2_3;

	wire horizontal_tile_6_2_to_tile_6_3_0;
	wire horizontal_tile_6_2_to_tile_6_3_1;
	wire horizontal_tile_6_2_to_tile_6_3_2;
	wire horizontal_tile_6_2_to_tile_6_3_3;
	wire horizontal_tile_6_3_to_tile_6_2_0;
	wire horizontal_tile_6_3_to_tile_6_2_1;
	wire horizontal_tile_6_3_to_tile_6_2_2;
	wire horizontal_tile_6_3_to_tile_6_2_3;

	wire horizontal_tile_7_2_to_tile_7_3_0;
	wire horizontal_tile_7_2_to_tile_7_3_1;
	wire horizontal_tile_7_2_to_tile_7_3_2;
	wire horizontal_tile_7_2_to_tile_7_3_3;
	wire horizontal_tile_7_3_to_tile_7_2_0;
	wire horizontal_tile_7_3_to_tile_7_2_1;
	wire horizontal_tile_7_3_to_tile_7_2_2;
	wire horizontal_tile_7_3_to_tile_7_2_3;

	wire horizontal_tile_8_2_to_tile_8_3_0;
	wire horizontal_tile_8_2_to_tile_8_3_1;
	wire horizontal_tile_8_2_to_tile_8_3_2;
	wire horizontal_tile_8_2_to_tile_8_3_3;
	wire horizontal_tile_8_3_to_tile_8_2_0;
	wire horizontal_tile_8_3_to_tile_8_2_1;
	wire horizontal_tile_8_3_to_tile_8_2_2;
	wire horizontal_tile_8_3_to_tile_8_2_3;

	wire horizontal_tile_9_2_to_tile_9_3_0;
	wire horizontal_tile_9_2_to_tile_9_3_1;
	wire horizontal_tile_9_2_to_tile_9_3_2;
	wire horizontal_tile_9_2_to_tile_9_3_3;
	wire horizontal_tile_9_3_to_tile_9_2_0;
	wire horizontal_tile_9_3_to_tile_9_2_1;
	wire horizontal_tile_9_3_to_tile_9_2_2;
	wire horizontal_tile_9_3_to_tile_9_2_3;

	wire horizontal_tile_10_2_to_tile_10_3_0;
	wire horizontal_tile_10_2_to_tile_10_3_1;
	wire horizontal_tile_10_2_to_tile_10_3_2;
	wire horizontal_tile_10_2_to_tile_10_3_3;
	wire horizontal_tile_10_3_to_tile_10_2_0;
	wire horizontal_tile_10_3_to_tile_10_2_1;
	wire horizontal_tile_10_3_to_tile_10_2_2;
	wire horizontal_tile_10_3_to_tile_10_2_3;

	wire horizontal_tile_11_2_to_tile_11_3_0;
	wire horizontal_tile_11_2_to_tile_11_3_1;
	wire horizontal_tile_11_2_to_tile_11_3_2;
	wire horizontal_tile_11_2_to_tile_11_3_3;
	wire horizontal_tile_11_3_to_tile_11_2_0;
	wire horizontal_tile_11_3_to_tile_11_2_1;
	wire horizontal_tile_11_3_to_tile_11_2_2;
	wire horizontal_tile_11_3_to_tile_11_2_3;

	wire horizontal_tile_12_2_to_tile_12_3_0;
	wire horizontal_tile_12_2_to_tile_12_3_1;
	wire horizontal_tile_12_2_to_tile_12_3_2;
	wire horizontal_tile_12_2_to_tile_12_3_3;
	wire horizontal_tile_12_3_to_tile_12_2_0;
	wire horizontal_tile_12_3_to_tile_12_2_1;
	wire horizontal_tile_12_3_to_tile_12_2_2;
	wire horizontal_tile_12_3_to_tile_12_2_3;

	wire horizontal_tile_13_2_to_tile_13_3_0;
	wire horizontal_tile_13_2_to_tile_13_3_1;
	wire horizontal_tile_13_2_to_tile_13_3_2;
	wire horizontal_tile_13_2_to_tile_13_3_3;
	wire horizontal_tile_13_3_to_tile_13_2_0;
	wire horizontal_tile_13_3_to_tile_13_2_1;
	wire horizontal_tile_13_3_to_tile_13_2_2;
	wire horizontal_tile_13_3_to_tile_13_2_3;

	wire horizontal_tile_14_2_to_tile_14_3_0;
	wire horizontal_tile_14_2_to_tile_14_3_1;
	wire horizontal_tile_14_2_to_tile_14_3_2;
	wire horizontal_tile_14_2_to_tile_14_3_3;
	wire horizontal_tile_14_3_to_tile_14_2_0;
	wire horizontal_tile_14_3_to_tile_14_2_1;
	wire horizontal_tile_14_3_to_tile_14_2_2;
	wire horizontal_tile_14_3_to_tile_14_2_3;

	wire horizontal_tile_15_2_to_tile_15_3_0;
	wire horizontal_tile_15_2_to_tile_15_3_1;
	wire horizontal_tile_15_2_to_tile_15_3_2;
	wire horizontal_tile_15_2_to_tile_15_3_3;
	wire horizontal_tile_15_3_to_tile_15_2_0;
	wire horizontal_tile_15_3_to_tile_15_2_1;
	wire horizontal_tile_15_3_to_tile_15_2_2;
	wire horizontal_tile_15_3_to_tile_15_2_3;

	wire horizontal_tile_16_2_to_tile_16_3_0;
	wire horizontal_tile_16_2_to_tile_16_3_1;
	wire horizontal_tile_16_2_to_tile_16_3_2;
	wire horizontal_tile_16_2_to_tile_16_3_3;
	wire horizontal_tile_16_3_to_tile_16_2_0;
	wire horizontal_tile_16_3_to_tile_16_2_1;
	wire horizontal_tile_16_3_to_tile_16_2_2;
	wire horizontal_tile_16_3_to_tile_16_2_3;

	wire horizontal_tile_17_2_to_tile_17_3_0;
	wire horizontal_tile_17_2_to_tile_17_3_1;
	wire horizontal_tile_17_2_to_tile_17_3_2;
	wire horizontal_tile_17_2_to_tile_17_3_3;
	wire horizontal_tile_17_3_to_tile_17_2_0;
	wire horizontal_tile_17_3_to_tile_17_2_1;
	wire horizontal_tile_17_3_to_tile_17_2_2;
	wire horizontal_tile_17_3_to_tile_17_2_3;

	wire horizontal_tile_18_2_to_tile_18_3_0;
	wire horizontal_tile_18_2_to_tile_18_3_1;
	wire horizontal_tile_18_2_to_tile_18_3_2;
	wire horizontal_tile_18_2_to_tile_18_3_3;
	wire horizontal_tile_18_3_to_tile_18_2_0;
	wire horizontal_tile_18_3_to_tile_18_2_1;
	wire horizontal_tile_18_3_to_tile_18_2_2;
	wire horizontal_tile_18_3_to_tile_18_2_3;

	wire horizontal_tile_19_2_to_tile_19_3_0;
	wire horizontal_tile_19_2_to_tile_19_3_1;
	wire horizontal_tile_19_2_to_tile_19_3_2;
	wire horizontal_tile_19_2_to_tile_19_3_3;
	wire horizontal_tile_19_3_to_tile_19_2_0;
	wire horizontal_tile_19_3_to_tile_19_2_1;
	wire horizontal_tile_19_3_to_tile_19_2_2;
	wire horizontal_tile_19_3_to_tile_19_2_3;

	wire horizontal_tile_20_2_to_tile_20_3_0;
	wire horizontal_tile_20_2_to_tile_20_3_1;
	wire horizontal_tile_20_2_to_tile_20_3_2;
	wire horizontal_tile_20_2_to_tile_20_3_3;
	wire horizontal_tile_20_3_to_tile_20_2_0;
	wire horizontal_tile_20_3_to_tile_20_2_1;
	wire horizontal_tile_20_3_to_tile_20_2_2;
	wire horizontal_tile_20_3_to_tile_20_2_3;

	wire horizontal_tile_21_2_to_tile_21_3_0;
	wire horizontal_tile_21_2_to_tile_21_3_1;
	wire horizontal_tile_21_2_to_tile_21_3_2;
	wire horizontal_tile_21_2_to_tile_21_3_3;
	wire horizontal_tile_21_3_to_tile_21_2_0;
	wire horizontal_tile_21_3_to_tile_21_2_1;
	wire horizontal_tile_21_3_to_tile_21_2_2;
	wire horizontal_tile_21_3_to_tile_21_2_3;

	wire horizontal_tile_22_2_to_tile_22_3_0;
	wire horizontal_tile_22_2_to_tile_22_3_1;
	wire horizontal_tile_22_2_to_tile_22_3_2;
	wire horizontal_tile_22_2_to_tile_22_3_3;
	wire horizontal_tile_22_3_to_tile_22_2_0;
	wire horizontal_tile_22_3_to_tile_22_2_1;
	wire horizontal_tile_22_3_to_tile_22_2_2;
	wire horizontal_tile_22_3_to_tile_22_2_3;

	wire horizontal_tile_23_2_to_tile_23_3_0;
	wire horizontal_tile_23_2_to_tile_23_3_1;
	wire horizontal_tile_23_2_to_tile_23_3_2;
	wire horizontal_tile_23_2_to_tile_23_3_3;
	wire horizontal_tile_23_3_to_tile_23_2_0;
	wire horizontal_tile_23_3_to_tile_23_2_1;
	wire horizontal_tile_23_3_to_tile_23_2_2;
	wire horizontal_tile_23_3_to_tile_23_2_3;

	wire horizontal_tile_24_2_to_tile_24_3_0;
	wire horizontal_tile_24_2_to_tile_24_3_1;
	wire horizontal_tile_24_2_to_tile_24_3_2;
	wire horizontal_tile_24_2_to_tile_24_3_3;
	wire horizontal_tile_24_3_to_tile_24_2_0;
	wire horizontal_tile_24_3_to_tile_24_2_1;
	wire horizontal_tile_24_3_to_tile_24_2_2;
	wire horizontal_tile_24_3_to_tile_24_2_3;

	wire horizontal_tile_25_2_to_tile_25_3_0;
	wire horizontal_tile_25_2_to_tile_25_3_1;
	wire horizontal_tile_25_2_to_tile_25_3_2;
	wire horizontal_tile_25_2_to_tile_25_3_3;
	wire horizontal_tile_25_3_to_tile_25_2_0;
	wire horizontal_tile_25_3_to_tile_25_2_1;
	wire horizontal_tile_25_3_to_tile_25_2_2;
	wire horizontal_tile_25_3_to_tile_25_2_3;

	wire horizontal_tile_26_2_to_tile_26_3_0;
	wire horizontal_tile_26_2_to_tile_26_3_1;
	wire horizontal_tile_26_2_to_tile_26_3_2;
	wire horizontal_tile_26_2_to_tile_26_3_3;
	wire horizontal_tile_26_3_to_tile_26_2_0;
	wire horizontal_tile_26_3_to_tile_26_2_1;
	wire horizontal_tile_26_3_to_tile_26_2_2;
	wire horizontal_tile_26_3_to_tile_26_2_3;

	wire horizontal_tile_27_2_to_tile_27_3_0;
	wire horizontal_tile_27_2_to_tile_27_3_1;
	wire horizontal_tile_27_2_to_tile_27_3_2;
	wire horizontal_tile_27_2_to_tile_27_3_3;
	wire horizontal_tile_27_3_to_tile_27_2_0;
	wire horizontal_tile_27_3_to_tile_27_2_1;
	wire horizontal_tile_27_3_to_tile_27_2_2;
	wire horizontal_tile_27_3_to_tile_27_2_3;

	wire horizontal_tile_28_2_to_tile_28_3_0;
	wire horizontal_tile_28_2_to_tile_28_3_1;
	wire horizontal_tile_28_2_to_tile_28_3_2;
	wire horizontal_tile_28_2_to_tile_28_3_3;
	wire horizontal_tile_28_3_to_tile_28_2_0;
	wire horizontal_tile_28_3_to_tile_28_2_1;
	wire horizontal_tile_28_3_to_tile_28_2_2;
	wire horizontal_tile_28_3_to_tile_28_2_3;

	wire horizontal_tile_29_2_to_tile_29_3_0;
	wire horizontal_tile_29_2_to_tile_29_3_1;
	wire horizontal_tile_29_2_to_tile_29_3_2;
	wire horizontal_tile_29_2_to_tile_29_3_3;
	wire horizontal_tile_29_3_to_tile_29_2_0;
	wire horizontal_tile_29_3_to_tile_29_2_1;
	wire horizontal_tile_29_3_to_tile_29_2_2;
	wire horizontal_tile_29_3_to_tile_29_2_3;

	wire horizontal_tile_30_2_to_tile_30_3_0;
	wire horizontal_tile_30_2_to_tile_30_3_1;
	wire horizontal_tile_30_2_to_tile_30_3_2;
	wire horizontal_tile_30_2_to_tile_30_3_3;
	wire horizontal_tile_30_3_to_tile_30_2_0;
	wire horizontal_tile_30_3_to_tile_30_2_1;
	wire horizontal_tile_30_3_to_tile_30_2_2;
	wire horizontal_tile_30_3_to_tile_30_2_3;

	wire horizontal_tile_31_2_to_tile_31_3_0;
	wire horizontal_tile_31_2_to_tile_31_3_1;
	wire horizontal_tile_31_2_to_tile_31_3_2;
	wire horizontal_tile_31_2_to_tile_31_3_3;
	wire horizontal_tile_31_3_to_tile_31_2_0;
	wire horizontal_tile_31_3_to_tile_31_2_1;
	wire horizontal_tile_31_3_to_tile_31_2_2;
	wire horizontal_tile_31_3_to_tile_31_2_3;

	wire horizontal_tile_0_3_to_tile_0_4_0;
	wire horizontal_tile_0_3_to_tile_0_4_1;
	wire horizontal_tile_0_3_to_tile_0_4_2;
	wire horizontal_tile_0_3_to_tile_0_4_3;
	wire horizontal_tile_0_4_to_tile_0_3_0;
	wire horizontal_tile_0_4_to_tile_0_3_1;
	wire horizontal_tile_0_4_to_tile_0_3_2;
	wire horizontal_tile_0_4_to_tile_0_3_3;

	wire horizontal_tile_1_3_to_tile_1_4_0;
	wire horizontal_tile_1_3_to_tile_1_4_1;
	wire horizontal_tile_1_3_to_tile_1_4_2;
	wire horizontal_tile_1_3_to_tile_1_4_3;
	wire horizontal_tile_1_4_to_tile_1_3_0;
	wire horizontal_tile_1_4_to_tile_1_3_1;
	wire horizontal_tile_1_4_to_tile_1_3_2;
	wire horizontal_tile_1_4_to_tile_1_3_3;

	wire horizontal_tile_2_3_to_tile_2_4_0;
	wire horizontal_tile_2_3_to_tile_2_4_1;
	wire horizontal_tile_2_3_to_tile_2_4_2;
	wire horizontal_tile_2_3_to_tile_2_4_3;
	wire horizontal_tile_2_4_to_tile_2_3_0;
	wire horizontal_tile_2_4_to_tile_2_3_1;
	wire horizontal_tile_2_4_to_tile_2_3_2;
	wire horizontal_tile_2_4_to_tile_2_3_3;

	wire horizontal_tile_3_3_to_tile_3_4_0;
	wire horizontal_tile_3_3_to_tile_3_4_1;
	wire horizontal_tile_3_3_to_tile_3_4_2;
	wire horizontal_tile_3_3_to_tile_3_4_3;
	wire horizontal_tile_3_4_to_tile_3_3_0;
	wire horizontal_tile_3_4_to_tile_3_3_1;
	wire horizontal_tile_3_4_to_tile_3_3_2;
	wire horizontal_tile_3_4_to_tile_3_3_3;

	wire horizontal_tile_4_3_to_tile_4_4_0;
	wire horizontal_tile_4_3_to_tile_4_4_1;
	wire horizontal_tile_4_3_to_tile_4_4_2;
	wire horizontal_tile_4_3_to_tile_4_4_3;
	wire horizontal_tile_4_4_to_tile_4_3_0;
	wire horizontal_tile_4_4_to_tile_4_3_1;
	wire horizontal_tile_4_4_to_tile_4_3_2;
	wire horizontal_tile_4_4_to_tile_4_3_3;

	wire horizontal_tile_5_3_to_tile_5_4_0;
	wire horizontal_tile_5_3_to_tile_5_4_1;
	wire horizontal_tile_5_3_to_tile_5_4_2;
	wire horizontal_tile_5_3_to_tile_5_4_3;
	wire horizontal_tile_5_4_to_tile_5_3_0;
	wire horizontal_tile_5_4_to_tile_5_3_1;
	wire horizontal_tile_5_4_to_tile_5_3_2;
	wire horizontal_tile_5_4_to_tile_5_3_3;

	wire horizontal_tile_6_3_to_tile_6_4_0;
	wire horizontal_tile_6_3_to_tile_6_4_1;
	wire horizontal_tile_6_3_to_tile_6_4_2;
	wire horizontal_tile_6_3_to_tile_6_4_3;
	wire horizontal_tile_6_4_to_tile_6_3_0;
	wire horizontal_tile_6_4_to_tile_6_3_1;
	wire horizontal_tile_6_4_to_tile_6_3_2;
	wire horizontal_tile_6_4_to_tile_6_3_3;

	wire horizontal_tile_7_3_to_tile_7_4_0;
	wire horizontal_tile_7_3_to_tile_7_4_1;
	wire horizontal_tile_7_3_to_tile_7_4_2;
	wire horizontal_tile_7_3_to_tile_7_4_3;
	wire horizontal_tile_7_4_to_tile_7_3_0;
	wire horizontal_tile_7_4_to_tile_7_3_1;
	wire horizontal_tile_7_4_to_tile_7_3_2;
	wire horizontal_tile_7_4_to_tile_7_3_3;

	wire horizontal_tile_8_3_to_tile_8_4_0;
	wire horizontal_tile_8_3_to_tile_8_4_1;
	wire horizontal_tile_8_3_to_tile_8_4_2;
	wire horizontal_tile_8_3_to_tile_8_4_3;
	wire horizontal_tile_8_4_to_tile_8_3_0;
	wire horizontal_tile_8_4_to_tile_8_3_1;
	wire horizontal_tile_8_4_to_tile_8_3_2;
	wire horizontal_tile_8_4_to_tile_8_3_3;

	wire horizontal_tile_9_3_to_tile_9_4_0;
	wire horizontal_tile_9_3_to_tile_9_4_1;
	wire horizontal_tile_9_3_to_tile_9_4_2;
	wire horizontal_tile_9_3_to_tile_9_4_3;
	wire horizontal_tile_9_4_to_tile_9_3_0;
	wire horizontal_tile_9_4_to_tile_9_3_1;
	wire horizontal_tile_9_4_to_tile_9_3_2;
	wire horizontal_tile_9_4_to_tile_9_3_3;

	wire horizontal_tile_10_3_to_tile_10_4_0;
	wire horizontal_tile_10_3_to_tile_10_4_1;
	wire horizontal_tile_10_3_to_tile_10_4_2;
	wire horizontal_tile_10_3_to_tile_10_4_3;
	wire horizontal_tile_10_4_to_tile_10_3_0;
	wire horizontal_tile_10_4_to_tile_10_3_1;
	wire horizontal_tile_10_4_to_tile_10_3_2;
	wire horizontal_tile_10_4_to_tile_10_3_3;

	wire horizontal_tile_11_3_to_tile_11_4_0;
	wire horizontal_tile_11_3_to_tile_11_4_1;
	wire horizontal_tile_11_3_to_tile_11_4_2;
	wire horizontal_tile_11_3_to_tile_11_4_3;
	wire horizontal_tile_11_4_to_tile_11_3_0;
	wire horizontal_tile_11_4_to_tile_11_3_1;
	wire horizontal_tile_11_4_to_tile_11_3_2;
	wire horizontal_tile_11_4_to_tile_11_3_3;

	wire horizontal_tile_12_3_to_tile_12_4_0;
	wire horizontal_tile_12_3_to_tile_12_4_1;
	wire horizontal_tile_12_3_to_tile_12_4_2;
	wire horizontal_tile_12_3_to_tile_12_4_3;
	wire horizontal_tile_12_4_to_tile_12_3_0;
	wire horizontal_tile_12_4_to_tile_12_3_1;
	wire horizontal_tile_12_4_to_tile_12_3_2;
	wire horizontal_tile_12_4_to_tile_12_3_3;

	wire horizontal_tile_13_3_to_tile_13_4_0;
	wire horizontal_tile_13_3_to_tile_13_4_1;
	wire horizontal_tile_13_3_to_tile_13_4_2;
	wire horizontal_tile_13_3_to_tile_13_4_3;
	wire horizontal_tile_13_4_to_tile_13_3_0;
	wire horizontal_tile_13_4_to_tile_13_3_1;
	wire horizontal_tile_13_4_to_tile_13_3_2;
	wire horizontal_tile_13_4_to_tile_13_3_3;

	wire horizontal_tile_14_3_to_tile_14_4_0;
	wire horizontal_tile_14_3_to_tile_14_4_1;
	wire horizontal_tile_14_3_to_tile_14_4_2;
	wire horizontal_tile_14_3_to_tile_14_4_3;
	wire horizontal_tile_14_4_to_tile_14_3_0;
	wire horizontal_tile_14_4_to_tile_14_3_1;
	wire horizontal_tile_14_4_to_tile_14_3_2;
	wire horizontal_tile_14_4_to_tile_14_3_3;

	wire horizontal_tile_15_3_to_tile_15_4_0;
	wire horizontal_tile_15_3_to_tile_15_4_1;
	wire horizontal_tile_15_3_to_tile_15_4_2;
	wire horizontal_tile_15_3_to_tile_15_4_3;
	wire horizontal_tile_15_4_to_tile_15_3_0;
	wire horizontal_tile_15_4_to_tile_15_3_1;
	wire horizontal_tile_15_4_to_tile_15_3_2;
	wire horizontal_tile_15_4_to_tile_15_3_3;

	wire horizontal_tile_16_3_to_tile_16_4_0;
	wire horizontal_tile_16_3_to_tile_16_4_1;
	wire horizontal_tile_16_3_to_tile_16_4_2;
	wire horizontal_tile_16_3_to_tile_16_4_3;
	wire horizontal_tile_16_4_to_tile_16_3_0;
	wire horizontal_tile_16_4_to_tile_16_3_1;
	wire horizontal_tile_16_4_to_tile_16_3_2;
	wire horizontal_tile_16_4_to_tile_16_3_3;

	wire horizontal_tile_17_3_to_tile_17_4_0;
	wire horizontal_tile_17_3_to_tile_17_4_1;
	wire horizontal_tile_17_3_to_tile_17_4_2;
	wire horizontal_tile_17_3_to_tile_17_4_3;
	wire horizontal_tile_17_4_to_tile_17_3_0;
	wire horizontal_tile_17_4_to_tile_17_3_1;
	wire horizontal_tile_17_4_to_tile_17_3_2;
	wire horizontal_tile_17_4_to_tile_17_3_3;

	wire horizontal_tile_18_3_to_tile_18_4_0;
	wire horizontal_tile_18_3_to_tile_18_4_1;
	wire horizontal_tile_18_3_to_tile_18_4_2;
	wire horizontal_tile_18_3_to_tile_18_4_3;
	wire horizontal_tile_18_4_to_tile_18_3_0;
	wire horizontal_tile_18_4_to_tile_18_3_1;
	wire horizontal_tile_18_4_to_tile_18_3_2;
	wire horizontal_tile_18_4_to_tile_18_3_3;

	wire horizontal_tile_19_3_to_tile_19_4_0;
	wire horizontal_tile_19_3_to_tile_19_4_1;
	wire horizontal_tile_19_3_to_tile_19_4_2;
	wire horizontal_tile_19_3_to_tile_19_4_3;
	wire horizontal_tile_19_4_to_tile_19_3_0;
	wire horizontal_tile_19_4_to_tile_19_3_1;
	wire horizontal_tile_19_4_to_tile_19_3_2;
	wire horizontal_tile_19_4_to_tile_19_3_3;

	wire horizontal_tile_20_3_to_tile_20_4_0;
	wire horizontal_tile_20_3_to_tile_20_4_1;
	wire horizontal_tile_20_3_to_tile_20_4_2;
	wire horizontal_tile_20_3_to_tile_20_4_3;
	wire horizontal_tile_20_4_to_tile_20_3_0;
	wire horizontal_tile_20_4_to_tile_20_3_1;
	wire horizontal_tile_20_4_to_tile_20_3_2;
	wire horizontal_tile_20_4_to_tile_20_3_3;

	wire horizontal_tile_21_3_to_tile_21_4_0;
	wire horizontal_tile_21_3_to_tile_21_4_1;
	wire horizontal_tile_21_3_to_tile_21_4_2;
	wire horizontal_tile_21_3_to_tile_21_4_3;
	wire horizontal_tile_21_4_to_tile_21_3_0;
	wire horizontal_tile_21_4_to_tile_21_3_1;
	wire horizontal_tile_21_4_to_tile_21_3_2;
	wire horizontal_tile_21_4_to_tile_21_3_3;

	wire horizontal_tile_22_3_to_tile_22_4_0;
	wire horizontal_tile_22_3_to_tile_22_4_1;
	wire horizontal_tile_22_3_to_tile_22_4_2;
	wire horizontal_tile_22_3_to_tile_22_4_3;
	wire horizontal_tile_22_4_to_tile_22_3_0;
	wire horizontal_tile_22_4_to_tile_22_3_1;
	wire horizontal_tile_22_4_to_tile_22_3_2;
	wire horizontal_tile_22_4_to_tile_22_3_3;

	wire horizontal_tile_23_3_to_tile_23_4_0;
	wire horizontal_tile_23_3_to_tile_23_4_1;
	wire horizontal_tile_23_3_to_tile_23_4_2;
	wire horizontal_tile_23_3_to_tile_23_4_3;
	wire horizontal_tile_23_4_to_tile_23_3_0;
	wire horizontal_tile_23_4_to_tile_23_3_1;
	wire horizontal_tile_23_4_to_tile_23_3_2;
	wire horizontal_tile_23_4_to_tile_23_3_3;

	wire horizontal_tile_24_3_to_tile_24_4_0;
	wire horizontal_tile_24_3_to_tile_24_4_1;
	wire horizontal_tile_24_3_to_tile_24_4_2;
	wire horizontal_tile_24_3_to_tile_24_4_3;
	wire horizontal_tile_24_4_to_tile_24_3_0;
	wire horizontal_tile_24_4_to_tile_24_3_1;
	wire horizontal_tile_24_4_to_tile_24_3_2;
	wire horizontal_tile_24_4_to_tile_24_3_3;

	wire horizontal_tile_25_3_to_tile_25_4_0;
	wire horizontal_tile_25_3_to_tile_25_4_1;
	wire horizontal_tile_25_3_to_tile_25_4_2;
	wire horizontal_tile_25_3_to_tile_25_4_3;
	wire horizontal_tile_25_4_to_tile_25_3_0;
	wire horizontal_tile_25_4_to_tile_25_3_1;
	wire horizontal_tile_25_4_to_tile_25_3_2;
	wire horizontal_tile_25_4_to_tile_25_3_3;

	wire horizontal_tile_26_3_to_tile_26_4_0;
	wire horizontal_tile_26_3_to_tile_26_4_1;
	wire horizontal_tile_26_3_to_tile_26_4_2;
	wire horizontal_tile_26_3_to_tile_26_4_3;
	wire horizontal_tile_26_4_to_tile_26_3_0;
	wire horizontal_tile_26_4_to_tile_26_3_1;
	wire horizontal_tile_26_4_to_tile_26_3_2;
	wire horizontal_tile_26_4_to_tile_26_3_3;

	wire horizontal_tile_27_3_to_tile_27_4_0;
	wire horizontal_tile_27_3_to_tile_27_4_1;
	wire horizontal_tile_27_3_to_tile_27_4_2;
	wire horizontal_tile_27_3_to_tile_27_4_3;
	wire horizontal_tile_27_4_to_tile_27_3_0;
	wire horizontal_tile_27_4_to_tile_27_3_1;
	wire horizontal_tile_27_4_to_tile_27_3_2;
	wire horizontal_tile_27_4_to_tile_27_3_3;

	wire horizontal_tile_28_3_to_tile_28_4_0;
	wire horizontal_tile_28_3_to_tile_28_4_1;
	wire horizontal_tile_28_3_to_tile_28_4_2;
	wire horizontal_tile_28_3_to_tile_28_4_3;
	wire horizontal_tile_28_4_to_tile_28_3_0;
	wire horizontal_tile_28_4_to_tile_28_3_1;
	wire horizontal_tile_28_4_to_tile_28_3_2;
	wire horizontal_tile_28_4_to_tile_28_3_3;

	wire horizontal_tile_29_3_to_tile_29_4_0;
	wire horizontal_tile_29_3_to_tile_29_4_1;
	wire horizontal_tile_29_3_to_tile_29_4_2;
	wire horizontal_tile_29_3_to_tile_29_4_3;
	wire horizontal_tile_29_4_to_tile_29_3_0;
	wire horizontal_tile_29_4_to_tile_29_3_1;
	wire horizontal_tile_29_4_to_tile_29_3_2;
	wire horizontal_tile_29_4_to_tile_29_3_3;

	wire horizontal_tile_30_3_to_tile_30_4_0;
	wire horizontal_tile_30_3_to_tile_30_4_1;
	wire horizontal_tile_30_3_to_tile_30_4_2;
	wire horizontal_tile_30_3_to_tile_30_4_3;
	wire horizontal_tile_30_4_to_tile_30_3_0;
	wire horizontal_tile_30_4_to_tile_30_3_1;
	wire horizontal_tile_30_4_to_tile_30_3_2;
	wire horizontal_tile_30_4_to_tile_30_3_3;

	wire horizontal_tile_31_3_to_tile_31_4_0;
	wire horizontal_tile_31_3_to_tile_31_4_1;
	wire horizontal_tile_31_3_to_tile_31_4_2;
	wire horizontal_tile_31_3_to_tile_31_4_3;
	wire horizontal_tile_31_4_to_tile_31_3_0;
	wire horizontal_tile_31_4_to_tile_31_3_1;
	wire horizontal_tile_31_4_to_tile_31_3_2;
	wire horizontal_tile_31_4_to_tile_31_3_3;

	wire horizontal_tile_0_4_to_tile_0_5_0;
	wire horizontal_tile_0_4_to_tile_0_5_1;
	wire horizontal_tile_0_4_to_tile_0_5_2;
	wire horizontal_tile_0_4_to_tile_0_5_3;
	wire horizontal_tile_0_5_to_tile_0_4_0;
	wire horizontal_tile_0_5_to_tile_0_4_1;
	wire horizontal_tile_0_5_to_tile_0_4_2;
	wire horizontal_tile_0_5_to_tile_0_4_3;

	wire horizontal_tile_1_4_to_tile_1_5_0;
	wire horizontal_tile_1_4_to_tile_1_5_1;
	wire horizontal_tile_1_4_to_tile_1_5_2;
	wire horizontal_tile_1_4_to_tile_1_5_3;
	wire horizontal_tile_1_5_to_tile_1_4_0;
	wire horizontal_tile_1_5_to_tile_1_4_1;
	wire horizontal_tile_1_5_to_tile_1_4_2;
	wire horizontal_tile_1_5_to_tile_1_4_3;

	wire horizontal_tile_2_4_to_tile_2_5_0;
	wire horizontal_tile_2_4_to_tile_2_5_1;
	wire horizontal_tile_2_4_to_tile_2_5_2;
	wire horizontal_tile_2_4_to_tile_2_5_3;
	wire horizontal_tile_2_5_to_tile_2_4_0;
	wire horizontal_tile_2_5_to_tile_2_4_1;
	wire horizontal_tile_2_5_to_tile_2_4_2;
	wire horizontal_tile_2_5_to_tile_2_4_3;

	wire horizontal_tile_3_4_to_tile_3_5_0;
	wire horizontal_tile_3_4_to_tile_3_5_1;
	wire horizontal_tile_3_4_to_tile_3_5_2;
	wire horizontal_tile_3_4_to_tile_3_5_3;
	wire horizontal_tile_3_5_to_tile_3_4_0;
	wire horizontal_tile_3_5_to_tile_3_4_1;
	wire horizontal_tile_3_5_to_tile_3_4_2;
	wire horizontal_tile_3_5_to_tile_3_4_3;

	wire horizontal_tile_4_4_to_tile_4_5_0;
	wire horizontal_tile_4_4_to_tile_4_5_1;
	wire horizontal_tile_4_4_to_tile_4_5_2;
	wire horizontal_tile_4_4_to_tile_4_5_3;
	wire horizontal_tile_4_5_to_tile_4_4_0;
	wire horizontal_tile_4_5_to_tile_4_4_1;
	wire horizontal_tile_4_5_to_tile_4_4_2;
	wire horizontal_tile_4_5_to_tile_4_4_3;

	wire horizontal_tile_5_4_to_tile_5_5_0;
	wire horizontal_tile_5_4_to_tile_5_5_1;
	wire horizontal_tile_5_4_to_tile_5_5_2;
	wire horizontal_tile_5_4_to_tile_5_5_3;
	wire horizontal_tile_5_5_to_tile_5_4_0;
	wire horizontal_tile_5_5_to_tile_5_4_1;
	wire horizontal_tile_5_5_to_tile_5_4_2;
	wire horizontal_tile_5_5_to_tile_5_4_3;

	wire horizontal_tile_6_4_to_tile_6_5_0;
	wire horizontal_tile_6_4_to_tile_6_5_1;
	wire horizontal_tile_6_4_to_tile_6_5_2;
	wire horizontal_tile_6_4_to_tile_6_5_3;
	wire horizontal_tile_6_5_to_tile_6_4_0;
	wire horizontal_tile_6_5_to_tile_6_4_1;
	wire horizontal_tile_6_5_to_tile_6_4_2;
	wire horizontal_tile_6_5_to_tile_6_4_3;

	wire horizontal_tile_7_4_to_tile_7_5_0;
	wire horizontal_tile_7_4_to_tile_7_5_1;
	wire horizontal_tile_7_4_to_tile_7_5_2;
	wire horizontal_tile_7_4_to_tile_7_5_3;
	wire horizontal_tile_7_5_to_tile_7_4_0;
	wire horizontal_tile_7_5_to_tile_7_4_1;
	wire horizontal_tile_7_5_to_tile_7_4_2;
	wire horizontal_tile_7_5_to_tile_7_4_3;

	wire horizontal_tile_8_4_to_tile_8_5_0;
	wire horizontal_tile_8_4_to_tile_8_5_1;
	wire horizontal_tile_8_4_to_tile_8_5_2;
	wire horizontal_tile_8_4_to_tile_8_5_3;
	wire horizontal_tile_8_5_to_tile_8_4_0;
	wire horizontal_tile_8_5_to_tile_8_4_1;
	wire horizontal_tile_8_5_to_tile_8_4_2;
	wire horizontal_tile_8_5_to_tile_8_4_3;

	wire horizontal_tile_9_4_to_tile_9_5_0;
	wire horizontal_tile_9_4_to_tile_9_5_1;
	wire horizontal_tile_9_4_to_tile_9_5_2;
	wire horizontal_tile_9_4_to_tile_9_5_3;
	wire horizontal_tile_9_5_to_tile_9_4_0;
	wire horizontal_tile_9_5_to_tile_9_4_1;
	wire horizontal_tile_9_5_to_tile_9_4_2;
	wire horizontal_tile_9_5_to_tile_9_4_3;

	wire horizontal_tile_10_4_to_tile_10_5_0;
	wire horizontal_tile_10_4_to_tile_10_5_1;
	wire horizontal_tile_10_4_to_tile_10_5_2;
	wire horizontal_tile_10_4_to_tile_10_5_3;
	wire horizontal_tile_10_5_to_tile_10_4_0;
	wire horizontal_tile_10_5_to_tile_10_4_1;
	wire horizontal_tile_10_5_to_tile_10_4_2;
	wire horizontal_tile_10_5_to_tile_10_4_3;

	wire horizontal_tile_11_4_to_tile_11_5_0;
	wire horizontal_tile_11_4_to_tile_11_5_1;
	wire horizontal_tile_11_4_to_tile_11_5_2;
	wire horizontal_tile_11_4_to_tile_11_5_3;
	wire horizontal_tile_11_5_to_tile_11_4_0;
	wire horizontal_tile_11_5_to_tile_11_4_1;
	wire horizontal_tile_11_5_to_tile_11_4_2;
	wire horizontal_tile_11_5_to_tile_11_4_3;

	wire horizontal_tile_12_4_to_tile_12_5_0;
	wire horizontal_tile_12_4_to_tile_12_5_1;
	wire horizontal_tile_12_4_to_tile_12_5_2;
	wire horizontal_tile_12_4_to_tile_12_5_3;
	wire horizontal_tile_12_5_to_tile_12_4_0;
	wire horizontal_tile_12_5_to_tile_12_4_1;
	wire horizontal_tile_12_5_to_tile_12_4_2;
	wire horizontal_tile_12_5_to_tile_12_4_3;

	wire horizontal_tile_13_4_to_tile_13_5_0;
	wire horizontal_tile_13_4_to_tile_13_5_1;
	wire horizontal_tile_13_4_to_tile_13_5_2;
	wire horizontal_tile_13_4_to_tile_13_5_3;
	wire horizontal_tile_13_5_to_tile_13_4_0;
	wire horizontal_tile_13_5_to_tile_13_4_1;
	wire horizontal_tile_13_5_to_tile_13_4_2;
	wire horizontal_tile_13_5_to_tile_13_4_3;

	wire horizontal_tile_14_4_to_tile_14_5_0;
	wire horizontal_tile_14_4_to_tile_14_5_1;
	wire horizontal_tile_14_4_to_tile_14_5_2;
	wire horizontal_tile_14_4_to_tile_14_5_3;
	wire horizontal_tile_14_5_to_tile_14_4_0;
	wire horizontal_tile_14_5_to_tile_14_4_1;
	wire horizontal_tile_14_5_to_tile_14_4_2;
	wire horizontal_tile_14_5_to_tile_14_4_3;

	wire horizontal_tile_15_4_to_tile_15_5_0;
	wire horizontal_tile_15_4_to_tile_15_5_1;
	wire horizontal_tile_15_4_to_tile_15_5_2;
	wire horizontal_tile_15_4_to_tile_15_5_3;
	wire horizontal_tile_15_5_to_tile_15_4_0;
	wire horizontal_tile_15_5_to_tile_15_4_1;
	wire horizontal_tile_15_5_to_tile_15_4_2;
	wire horizontal_tile_15_5_to_tile_15_4_3;

	wire horizontal_tile_16_4_to_tile_16_5_0;
	wire horizontal_tile_16_4_to_tile_16_5_1;
	wire horizontal_tile_16_4_to_tile_16_5_2;
	wire horizontal_tile_16_4_to_tile_16_5_3;
	wire horizontal_tile_16_5_to_tile_16_4_0;
	wire horizontal_tile_16_5_to_tile_16_4_1;
	wire horizontal_tile_16_5_to_tile_16_4_2;
	wire horizontal_tile_16_5_to_tile_16_4_3;

	wire horizontal_tile_17_4_to_tile_17_5_0;
	wire horizontal_tile_17_4_to_tile_17_5_1;
	wire horizontal_tile_17_4_to_tile_17_5_2;
	wire horizontal_tile_17_4_to_tile_17_5_3;
	wire horizontal_tile_17_5_to_tile_17_4_0;
	wire horizontal_tile_17_5_to_tile_17_4_1;
	wire horizontal_tile_17_5_to_tile_17_4_2;
	wire horizontal_tile_17_5_to_tile_17_4_3;

	wire horizontal_tile_18_4_to_tile_18_5_0;
	wire horizontal_tile_18_4_to_tile_18_5_1;
	wire horizontal_tile_18_4_to_tile_18_5_2;
	wire horizontal_tile_18_4_to_tile_18_5_3;
	wire horizontal_tile_18_5_to_tile_18_4_0;
	wire horizontal_tile_18_5_to_tile_18_4_1;
	wire horizontal_tile_18_5_to_tile_18_4_2;
	wire horizontal_tile_18_5_to_tile_18_4_3;

	wire horizontal_tile_19_4_to_tile_19_5_0;
	wire horizontal_tile_19_4_to_tile_19_5_1;
	wire horizontal_tile_19_4_to_tile_19_5_2;
	wire horizontal_tile_19_4_to_tile_19_5_3;
	wire horizontal_tile_19_5_to_tile_19_4_0;
	wire horizontal_tile_19_5_to_tile_19_4_1;
	wire horizontal_tile_19_5_to_tile_19_4_2;
	wire horizontal_tile_19_5_to_tile_19_4_3;

	wire horizontal_tile_20_4_to_tile_20_5_0;
	wire horizontal_tile_20_4_to_tile_20_5_1;
	wire horizontal_tile_20_4_to_tile_20_5_2;
	wire horizontal_tile_20_4_to_tile_20_5_3;
	wire horizontal_tile_20_5_to_tile_20_4_0;
	wire horizontal_tile_20_5_to_tile_20_4_1;
	wire horizontal_tile_20_5_to_tile_20_4_2;
	wire horizontal_tile_20_5_to_tile_20_4_3;

	wire horizontal_tile_21_4_to_tile_21_5_0;
	wire horizontal_tile_21_4_to_tile_21_5_1;
	wire horizontal_tile_21_4_to_tile_21_5_2;
	wire horizontal_tile_21_4_to_tile_21_5_3;
	wire horizontal_tile_21_5_to_tile_21_4_0;
	wire horizontal_tile_21_5_to_tile_21_4_1;
	wire horizontal_tile_21_5_to_tile_21_4_2;
	wire horizontal_tile_21_5_to_tile_21_4_3;

	wire horizontal_tile_22_4_to_tile_22_5_0;
	wire horizontal_tile_22_4_to_tile_22_5_1;
	wire horizontal_tile_22_4_to_tile_22_5_2;
	wire horizontal_tile_22_4_to_tile_22_5_3;
	wire horizontal_tile_22_5_to_tile_22_4_0;
	wire horizontal_tile_22_5_to_tile_22_4_1;
	wire horizontal_tile_22_5_to_tile_22_4_2;
	wire horizontal_tile_22_5_to_tile_22_4_3;

	wire horizontal_tile_23_4_to_tile_23_5_0;
	wire horizontal_tile_23_4_to_tile_23_5_1;
	wire horizontal_tile_23_4_to_tile_23_5_2;
	wire horizontal_tile_23_4_to_tile_23_5_3;
	wire horizontal_tile_23_5_to_tile_23_4_0;
	wire horizontal_tile_23_5_to_tile_23_4_1;
	wire horizontal_tile_23_5_to_tile_23_4_2;
	wire horizontal_tile_23_5_to_tile_23_4_3;

	wire horizontal_tile_24_4_to_tile_24_5_0;
	wire horizontal_tile_24_4_to_tile_24_5_1;
	wire horizontal_tile_24_4_to_tile_24_5_2;
	wire horizontal_tile_24_4_to_tile_24_5_3;
	wire horizontal_tile_24_5_to_tile_24_4_0;
	wire horizontal_tile_24_5_to_tile_24_4_1;
	wire horizontal_tile_24_5_to_tile_24_4_2;
	wire horizontal_tile_24_5_to_tile_24_4_3;

	wire horizontal_tile_25_4_to_tile_25_5_0;
	wire horizontal_tile_25_4_to_tile_25_5_1;
	wire horizontal_tile_25_4_to_tile_25_5_2;
	wire horizontal_tile_25_4_to_tile_25_5_3;
	wire horizontal_tile_25_5_to_tile_25_4_0;
	wire horizontal_tile_25_5_to_tile_25_4_1;
	wire horizontal_tile_25_5_to_tile_25_4_2;
	wire horizontal_tile_25_5_to_tile_25_4_3;

	wire horizontal_tile_26_4_to_tile_26_5_0;
	wire horizontal_tile_26_4_to_tile_26_5_1;
	wire horizontal_tile_26_4_to_tile_26_5_2;
	wire horizontal_tile_26_4_to_tile_26_5_3;
	wire horizontal_tile_26_5_to_tile_26_4_0;
	wire horizontal_tile_26_5_to_tile_26_4_1;
	wire horizontal_tile_26_5_to_tile_26_4_2;
	wire horizontal_tile_26_5_to_tile_26_4_3;

	wire horizontal_tile_27_4_to_tile_27_5_0;
	wire horizontal_tile_27_4_to_tile_27_5_1;
	wire horizontal_tile_27_4_to_tile_27_5_2;
	wire horizontal_tile_27_4_to_tile_27_5_3;
	wire horizontal_tile_27_5_to_tile_27_4_0;
	wire horizontal_tile_27_5_to_tile_27_4_1;
	wire horizontal_tile_27_5_to_tile_27_4_2;
	wire horizontal_tile_27_5_to_tile_27_4_3;

	wire horizontal_tile_28_4_to_tile_28_5_0;
	wire horizontal_tile_28_4_to_tile_28_5_1;
	wire horizontal_tile_28_4_to_tile_28_5_2;
	wire horizontal_tile_28_4_to_tile_28_5_3;
	wire horizontal_tile_28_5_to_tile_28_4_0;
	wire horizontal_tile_28_5_to_tile_28_4_1;
	wire horizontal_tile_28_5_to_tile_28_4_2;
	wire horizontal_tile_28_5_to_tile_28_4_3;

	wire horizontal_tile_29_4_to_tile_29_5_0;
	wire horizontal_tile_29_4_to_tile_29_5_1;
	wire horizontal_tile_29_4_to_tile_29_5_2;
	wire horizontal_tile_29_4_to_tile_29_5_3;
	wire horizontal_tile_29_5_to_tile_29_4_0;
	wire horizontal_tile_29_5_to_tile_29_4_1;
	wire horizontal_tile_29_5_to_tile_29_4_2;
	wire horizontal_tile_29_5_to_tile_29_4_3;

	wire horizontal_tile_30_4_to_tile_30_5_0;
	wire horizontal_tile_30_4_to_tile_30_5_1;
	wire horizontal_tile_30_4_to_tile_30_5_2;
	wire horizontal_tile_30_4_to_tile_30_5_3;
	wire horizontal_tile_30_5_to_tile_30_4_0;
	wire horizontal_tile_30_5_to_tile_30_4_1;
	wire horizontal_tile_30_5_to_tile_30_4_2;
	wire horizontal_tile_30_5_to_tile_30_4_3;

	wire horizontal_tile_31_4_to_tile_31_5_0;
	wire horizontal_tile_31_4_to_tile_31_5_1;
	wire horizontal_tile_31_4_to_tile_31_5_2;
	wire horizontal_tile_31_4_to_tile_31_5_3;
	wire horizontal_tile_31_5_to_tile_31_4_0;
	wire horizontal_tile_31_5_to_tile_31_4_1;
	wire horizontal_tile_31_5_to_tile_31_4_2;
	wire horizontal_tile_31_5_to_tile_31_4_3;

	wire horizontal_tile_0_5_to_tile_0_6_0;
	wire horizontal_tile_0_5_to_tile_0_6_1;
	wire horizontal_tile_0_5_to_tile_0_6_2;
	wire horizontal_tile_0_5_to_tile_0_6_3;
	wire horizontal_tile_0_6_to_tile_0_5_0;
	wire horizontal_tile_0_6_to_tile_0_5_1;
	wire horizontal_tile_0_6_to_tile_0_5_2;
	wire horizontal_tile_0_6_to_tile_0_5_3;

	wire horizontal_tile_1_5_to_tile_1_6_0;
	wire horizontal_tile_1_5_to_tile_1_6_1;
	wire horizontal_tile_1_5_to_tile_1_6_2;
	wire horizontal_tile_1_5_to_tile_1_6_3;
	wire horizontal_tile_1_6_to_tile_1_5_0;
	wire horizontal_tile_1_6_to_tile_1_5_1;
	wire horizontal_tile_1_6_to_tile_1_5_2;
	wire horizontal_tile_1_6_to_tile_1_5_3;

	wire horizontal_tile_2_5_to_tile_2_6_0;
	wire horizontal_tile_2_5_to_tile_2_6_1;
	wire horizontal_tile_2_5_to_tile_2_6_2;
	wire horizontal_tile_2_5_to_tile_2_6_3;
	wire horizontal_tile_2_6_to_tile_2_5_0;
	wire horizontal_tile_2_6_to_tile_2_5_1;
	wire horizontal_tile_2_6_to_tile_2_5_2;
	wire horizontal_tile_2_6_to_tile_2_5_3;

	wire horizontal_tile_3_5_to_tile_3_6_0;
	wire horizontal_tile_3_5_to_tile_3_6_1;
	wire horizontal_tile_3_5_to_tile_3_6_2;
	wire horizontal_tile_3_5_to_tile_3_6_3;
	wire horizontal_tile_3_6_to_tile_3_5_0;
	wire horizontal_tile_3_6_to_tile_3_5_1;
	wire horizontal_tile_3_6_to_tile_3_5_2;
	wire horizontal_tile_3_6_to_tile_3_5_3;

	wire horizontal_tile_4_5_to_tile_4_6_0;
	wire horizontal_tile_4_5_to_tile_4_6_1;
	wire horizontal_tile_4_5_to_tile_4_6_2;
	wire horizontal_tile_4_5_to_tile_4_6_3;
	wire horizontal_tile_4_6_to_tile_4_5_0;
	wire horizontal_tile_4_6_to_tile_4_5_1;
	wire horizontal_tile_4_6_to_tile_4_5_2;
	wire horizontal_tile_4_6_to_tile_4_5_3;

	wire horizontal_tile_5_5_to_tile_5_6_0;
	wire horizontal_tile_5_5_to_tile_5_6_1;
	wire horizontal_tile_5_5_to_tile_5_6_2;
	wire horizontal_tile_5_5_to_tile_5_6_3;
	wire horizontal_tile_5_6_to_tile_5_5_0;
	wire horizontal_tile_5_6_to_tile_5_5_1;
	wire horizontal_tile_5_6_to_tile_5_5_2;
	wire horizontal_tile_5_6_to_tile_5_5_3;

	wire horizontal_tile_6_5_to_tile_6_6_0;
	wire horizontal_tile_6_5_to_tile_6_6_1;
	wire horizontal_tile_6_5_to_tile_6_6_2;
	wire horizontal_tile_6_5_to_tile_6_6_3;
	wire horizontal_tile_6_6_to_tile_6_5_0;
	wire horizontal_tile_6_6_to_tile_6_5_1;
	wire horizontal_tile_6_6_to_tile_6_5_2;
	wire horizontal_tile_6_6_to_tile_6_5_3;

	wire horizontal_tile_7_5_to_tile_7_6_0;
	wire horizontal_tile_7_5_to_tile_7_6_1;
	wire horizontal_tile_7_5_to_tile_7_6_2;
	wire horizontal_tile_7_5_to_tile_7_6_3;
	wire horizontal_tile_7_6_to_tile_7_5_0;
	wire horizontal_tile_7_6_to_tile_7_5_1;
	wire horizontal_tile_7_6_to_tile_7_5_2;
	wire horizontal_tile_7_6_to_tile_7_5_3;

	wire horizontal_tile_8_5_to_tile_8_6_0;
	wire horizontal_tile_8_5_to_tile_8_6_1;
	wire horizontal_tile_8_5_to_tile_8_6_2;
	wire horizontal_tile_8_5_to_tile_8_6_3;
	wire horizontal_tile_8_6_to_tile_8_5_0;
	wire horizontal_tile_8_6_to_tile_8_5_1;
	wire horizontal_tile_8_6_to_tile_8_5_2;
	wire horizontal_tile_8_6_to_tile_8_5_3;

	wire horizontal_tile_9_5_to_tile_9_6_0;
	wire horizontal_tile_9_5_to_tile_9_6_1;
	wire horizontal_tile_9_5_to_tile_9_6_2;
	wire horizontal_tile_9_5_to_tile_9_6_3;
	wire horizontal_tile_9_6_to_tile_9_5_0;
	wire horizontal_tile_9_6_to_tile_9_5_1;
	wire horizontal_tile_9_6_to_tile_9_5_2;
	wire horizontal_tile_9_6_to_tile_9_5_3;

	wire horizontal_tile_10_5_to_tile_10_6_0;
	wire horizontal_tile_10_5_to_tile_10_6_1;
	wire horizontal_tile_10_5_to_tile_10_6_2;
	wire horizontal_tile_10_5_to_tile_10_6_3;
	wire horizontal_tile_10_6_to_tile_10_5_0;
	wire horizontal_tile_10_6_to_tile_10_5_1;
	wire horizontal_tile_10_6_to_tile_10_5_2;
	wire horizontal_tile_10_6_to_tile_10_5_3;

	wire horizontal_tile_11_5_to_tile_11_6_0;
	wire horizontal_tile_11_5_to_tile_11_6_1;
	wire horizontal_tile_11_5_to_tile_11_6_2;
	wire horizontal_tile_11_5_to_tile_11_6_3;
	wire horizontal_tile_11_6_to_tile_11_5_0;
	wire horizontal_tile_11_6_to_tile_11_5_1;
	wire horizontal_tile_11_6_to_tile_11_5_2;
	wire horizontal_tile_11_6_to_tile_11_5_3;

	wire horizontal_tile_12_5_to_tile_12_6_0;
	wire horizontal_tile_12_5_to_tile_12_6_1;
	wire horizontal_tile_12_5_to_tile_12_6_2;
	wire horizontal_tile_12_5_to_tile_12_6_3;
	wire horizontal_tile_12_6_to_tile_12_5_0;
	wire horizontal_tile_12_6_to_tile_12_5_1;
	wire horizontal_tile_12_6_to_tile_12_5_2;
	wire horizontal_tile_12_6_to_tile_12_5_3;

	wire horizontal_tile_13_5_to_tile_13_6_0;
	wire horizontal_tile_13_5_to_tile_13_6_1;
	wire horizontal_tile_13_5_to_tile_13_6_2;
	wire horizontal_tile_13_5_to_tile_13_6_3;
	wire horizontal_tile_13_6_to_tile_13_5_0;
	wire horizontal_tile_13_6_to_tile_13_5_1;
	wire horizontal_tile_13_6_to_tile_13_5_2;
	wire horizontal_tile_13_6_to_tile_13_5_3;

	wire horizontal_tile_14_5_to_tile_14_6_0;
	wire horizontal_tile_14_5_to_tile_14_6_1;
	wire horizontal_tile_14_5_to_tile_14_6_2;
	wire horizontal_tile_14_5_to_tile_14_6_3;
	wire horizontal_tile_14_6_to_tile_14_5_0;
	wire horizontal_tile_14_6_to_tile_14_5_1;
	wire horizontal_tile_14_6_to_tile_14_5_2;
	wire horizontal_tile_14_6_to_tile_14_5_3;

	wire horizontal_tile_15_5_to_tile_15_6_0;
	wire horizontal_tile_15_5_to_tile_15_6_1;
	wire horizontal_tile_15_5_to_tile_15_6_2;
	wire horizontal_tile_15_5_to_tile_15_6_3;
	wire horizontal_tile_15_6_to_tile_15_5_0;
	wire horizontal_tile_15_6_to_tile_15_5_1;
	wire horizontal_tile_15_6_to_tile_15_5_2;
	wire horizontal_tile_15_6_to_tile_15_5_3;

	wire horizontal_tile_16_5_to_tile_16_6_0;
	wire horizontal_tile_16_5_to_tile_16_6_1;
	wire horizontal_tile_16_5_to_tile_16_6_2;
	wire horizontal_tile_16_5_to_tile_16_6_3;
	wire horizontal_tile_16_6_to_tile_16_5_0;
	wire horizontal_tile_16_6_to_tile_16_5_1;
	wire horizontal_tile_16_6_to_tile_16_5_2;
	wire horizontal_tile_16_6_to_tile_16_5_3;

	wire horizontal_tile_17_5_to_tile_17_6_0;
	wire horizontal_tile_17_5_to_tile_17_6_1;
	wire horizontal_tile_17_5_to_tile_17_6_2;
	wire horizontal_tile_17_5_to_tile_17_6_3;
	wire horizontal_tile_17_6_to_tile_17_5_0;
	wire horizontal_tile_17_6_to_tile_17_5_1;
	wire horizontal_tile_17_6_to_tile_17_5_2;
	wire horizontal_tile_17_6_to_tile_17_5_3;

	wire horizontal_tile_18_5_to_tile_18_6_0;
	wire horizontal_tile_18_5_to_tile_18_6_1;
	wire horizontal_tile_18_5_to_tile_18_6_2;
	wire horizontal_tile_18_5_to_tile_18_6_3;
	wire horizontal_tile_18_6_to_tile_18_5_0;
	wire horizontal_tile_18_6_to_tile_18_5_1;
	wire horizontal_tile_18_6_to_tile_18_5_2;
	wire horizontal_tile_18_6_to_tile_18_5_3;

	wire horizontal_tile_19_5_to_tile_19_6_0;
	wire horizontal_tile_19_5_to_tile_19_6_1;
	wire horizontal_tile_19_5_to_tile_19_6_2;
	wire horizontal_tile_19_5_to_tile_19_6_3;
	wire horizontal_tile_19_6_to_tile_19_5_0;
	wire horizontal_tile_19_6_to_tile_19_5_1;
	wire horizontal_tile_19_6_to_tile_19_5_2;
	wire horizontal_tile_19_6_to_tile_19_5_3;

	wire horizontal_tile_20_5_to_tile_20_6_0;
	wire horizontal_tile_20_5_to_tile_20_6_1;
	wire horizontal_tile_20_5_to_tile_20_6_2;
	wire horizontal_tile_20_5_to_tile_20_6_3;
	wire horizontal_tile_20_6_to_tile_20_5_0;
	wire horizontal_tile_20_6_to_tile_20_5_1;
	wire horizontal_tile_20_6_to_tile_20_5_2;
	wire horizontal_tile_20_6_to_tile_20_5_3;

	wire horizontal_tile_21_5_to_tile_21_6_0;
	wire horizontal_tile_21_5_to_tile_21_6_1;
	wire horizontal_tile_21_5_to_tile_21_6_2;
	wire horizontal_tile_21_5_to_tile_21_6_3;
	wire horizontal_tile_21_6_to_tile_21_5_0;
	wire horizontal_tile_21_6_to_tile_21_5_1;
	wire horizontal_tile_21_6_to_tile_21_5_2;
	wire horizontal_tile_21_6_to_tile_21_5_3;

	wire horizontal_tile_22_5_to_tile_22_6_0;
	wire horizontal_tile_22_5_to_tile_22_6_1;
	wire horizontal_tile_22_5_to_tile_22_6_2;
	wire horizontal_tile_22_5_to_tile_22_6_3;
	wire horizontal_tile_22_6_to_tile_22_5_0;
	wire horizontal_tile_22_6_to_tile_22_5_1;
	wire horizontal_tile_22_6_to_tile_22_5_2;
	wire horizontal_tile_22_6_to_tile_22_5_3;

	wire horizontal_tile_23_5_to_tile_23_6_0;
	wire horizontal_tile_23_5_to_tile_23_6_1;
	wire horizontal_tile_23_5_to_tile_23_6_2;
	wire horizontal_tile_23_5_to_tile_23_6_3;
	wire horizontal_tile_23_6_to_tile_23_5_0;
	wire horizontal_tile_23_6_to_tile_23_5_1;
	wire horizontal_tile_23_6_to_tile_23_5_2;
	wire horizontal_tile_23_6_to_tile_23_5_3;

	wire horizontal_tile_24_5_to_tile_24_6_0;
	wire horizontal_tile_24_5_to_tile_24_6_1;
	wire horizontal_tile_24_5_to_tile_24_6_2;
	wire horizontal_tile_24_5_to_tile_24_6_3;
	wire horizontal_tile_24_6_to_tile_24_5_0;
	wire horizontal_tile_24_6_to_tile_24_5_1;
	wire horizontal_tile_24_6_to_tile_24_5_2;
	wire horizontal_tile_24_6_to_tile_24_5_3;

	wire horizontal_tile_25_5_to_tile_25_6_0;
	wire horizontal_tile_25_5_to_tile_25_6_1;
	wire horizontal_tile_25_5_to_tile_25_6_2;
	wire horizontal_tile_25_5_to_tile_25_6_3;
	wire horizontal_tile_25_6_to_tile_25_5_0;
	wire horizontal_tile_25_6_to_tile_25_5_1;
	wire horizontal_tile_25_6_to_tile_25_5_2;
	wire horizontal_tile_25_6_to_tile_25_5_3;

	wire horizontal_tile_26_5_to_tile_26_6_0;
	wire horizontal_tile_26_5_to_tile_26_6_1;
	wire horizontal_tile_26_5_to_tile_26_6_2;
	wire horizontal_tile_26_5_to_tile_26_6_3;
	wire horizontal_tile_26_6_to_tile_26_5_0;
	wire horizontal_tile_26_6_to_tile_26_5_1;
	wire horizontal_tile_26_6_to_tile_26_5_2;
	wire horizontal_tile_26_6_to_tile_26_5_3;

	wire horizontal_tile_27_5_to_tile_27_6_0;
	wire horizontal_tile_27_5_to_tile_27_6_1;
	wire horizontal_tile_27_5_to_tile_27_6_2;
	wire horizontal_tile_27_5_to_tile_27_6_3;
	wire horizontal_tile_27_6_to_tile_27_5_0;
	wire horizontal_tile_27_6_to_tile_27_5_1;
	wire horizontal_tile_27_6_to_tile_27_5_2;
	wire horizontal_tile_27_6_to_tile_27_5_3;

	wire horizontal_tile_28_5_to_tile_28_6_0;
	wire horizontal_tile_28_5_to_tile_28_6_1;
	wire horizontal_tile_28_5_to_tile_28_6_2;
	wire horizontal_tile_28_5_to_tile_28_6_3;
	wire horizontal_tile_28_6_to_tile_28_5_0;
	wire horizontal_tile_28_6_to_tile_28_5_1;
	wire horizontal_tile_28_6_to_tile_28_5_2;
	wire horizontal_tile_28_6_to_tile_28_5_3;

	wire horizontal_tile_29_5_to_tile_29_6_0;
	wire horizontal_tile_29_5_to_tile_29_6_1;
	wire horizontal_tile_29_5_to_tile_29_6_2;
	wire horizontal_tile_29_5_to_tile_29_6_3;
	wire horizontal_tile_29_6_to_tile_29_5_0;
	wire horizontal_tile_29_6_to_tile_29_5_1;
	wire horizontal_tile_29_6_to_tile_29_5_2;
	wire horizontal_tile_29_6_to_tile_29_5_3;

	wire horizontal_tile_30_5_to_tile_30_6_0;
	wire horizontal_tile_30_5_to_tile_30_6_1;
	wire horizontal_tile_30_5_to_tile_30_6_2;
	wire horizontal_tile_30_5_to_tile_30_6_3;
	wire horizontal_tile_30_6_to_tile_30_5_0;
	wire horizontal_tile_30_6_to_tile_30_5_1;
	wire horizontal_tile_30_6_to_tile_30_5_2;
	wire horizontal_tile_30_6_to_tile_30_5_3;

	wire horizontal_tile_31_5_to_tile_31_6_0;
	wire horizontal_tile_31_5_to_tile_31_6_1;
	wire horizontal_tile_31_5_to_tile_31_6_2;
	wire horizontal_tile_31_5_to_tile_31_6_3;
	wire horizontal_tile_31_6_to_tile_31_5_0;
	wire horizontal_tile_31_6_to_tile_31_5_1;
	wire horizontal_tile_31_6_to_tile_31_5_2;
	wire horizontal_tile_31_6_to_tile_31_5_3;

	wire horizontal_tile_0_6_to_tile_0_7_0;
	wire horizontal_tile_0_6_to_tile_0_7_1;
	wire horizontal_tile_0_6_to_tile_0_7_2;
	wire horizontal_tile_0_6_to_tile_0_7_3;
	wire horizontal_tile_0_7_to_tile_0_6_0;
	wire horizontal_tile_0_7_to_tile_0_6_1;
	wire horizontal_tile_0_7_to_tile_0_6_2;
	wire horizontal_tile_0_7_to_tile_0_6_3;

	wire horizontal_tile_1_6_to_tile_1_7_0;
	wire horizontal_tile_1_6_to_tile_1_7_1;
	wire horizontal_tile_1_6_to_tile_1_7_2;
	wire horizontal_tile_1_6_to_tile_1_7_3;
	wire horizontal_tile_1_7_to_tile_1_6_0;
	wire horizontal_tile_1_7_to_tile_1_6_1;
	wire horizontal_tile_1_7_to_tile_1_6_2;
	wire horizontal_tile_1_7_to_tile_1_6_3;

	wire horizontal_tile_2_6_to_tile_2_7_0;
	wire horizontal_tile_2_6_to_tile_2_7_1;
	wire horizontal_tile_2_6_to_tile_2_7_2;
	wire horizontal_tile_2_6_to_tile_2_7_3;
	wire horizontal_tile_2_7_to_tile_2_6_0;
	wire horizontal_tile_2_7_to_tile_2_6_1;
	wire horizontal_tile_2_7_to_tile_2_6_2;
	wire horizontal_tile_2_7_to_tile_2_6_3;

	wire horizontal_tile_3_6_to_tile_3_7_0;
	wire horizontal_tile_3_6_to_tile_3_7_1;
	wire horizontal_tile_3_6_to_tile_3_7_2;
	wire horizontal_tile_3_6_to_tile_3_7_3;
	wire horizontal_tile_3_7_to_tile_3_6_0;
	wire horizontal_tile_3_7_to_tile_3_6_1;
	wire horizontal_tile_3_7_to_tile_3_6_2;
	wire horizontal_tile_3_7_to_tile_3_6_3;

	wire horizontal_tile_4_6_to_tile_4_7_0;
	wire horizontal_tile_4_6_to_tile_4_7_1;
	wire horizontal_tile_4_6_to_tile_4_7_2;
	wire horizontal_tile_4_6_to_tile_4_7_3;
	wire horizontal_tile_4_7_to_tile_4_6_0;
	wire horizontal_tile_4_7_to_tile_4_6_1;
	wire horizontal_tile_4_7_to_tile_4_6_2;
	wire horizontal_tile_4_7_to_tile_4_6_3;

	wire horizontal_tile_5_6_to_tile_5_7_0;
	wire horizontal_tile_5_6_to_tile_5_7_1;
	wire horizontal_tile_5_6_to_tile_5_7_2;
	wire horizontal_tile_5_6_to_tile_5_7_3;
	wire horizontal_tile_5_7_to_tile_5_6_0;
	wire horizontal_tile_5_7_to_tile_5_6_1;
	wire horizontal_tile_5_7_to_tile_5_6_2;
	wire horizontal_tile_5_7_to_tile_5_6_3;

	wire horizontal_tile_6_6_to_tile_6_7_0;
	wire horizontal_tile_6_6_to_tile_6_7_1;
	wire horizontal_tile_6_6_to_tile_6_7_2;
	wire horizontal_tile_6_6_to_tile_6_7_3;
	wire horizontal_tile_6_7_to_tile_6_6_0;
	wire horizontal_tile_6_7_to_tile_6_6_1;
	wire horizontal_tile_6_7_to_tile_6_6_2;
	wire horizontal_tile_6_7_to_tile_6_6_3;

	wire horizontal_tile_7_6_to_tile_7_7_0;
	wire horizontal_tile_7_6_to_tile_7_7_1;
	wire horizontal_tile_7_6_to_tile_7_7_2;
	wire horizontal_tile_7_6_to_tile_7_7_3;
	wire horizontal_tile_7_7_to_tile_7_6_0;
	wire horizontal_tile_7_7_to_tile_7_6_1;
	wire horizontal_tile_7_7_to_tile_7_6_2;
	wire horizontal_tile_7_7_to_tile_7_6_3;

	wire horizontal_tile_8_6_to_tile_8_7_0;
	wire horizontal_tile_8_6_to_tile_8_7_1;
	wire horizontal_tile_8_6_to_tile_8_7_2;
	wire horizontal_tile_8_6_to_tile_8_7_3;
	wire horizontal_tile_8_7_to_tile_8_6_0;
	wire horizontal_tile_8_7_to_tile_8_6_1;
	wire horizontal_tile_8_7_to_tile_8_6_2;
	wire horizontal_tile_8_7_to_tile_8_6_3;

	wire horizontal_tile_9_6_to_tile_9_7_0;
	wire horizontal_tile_9_6_to_tile_9_7_1;
	wire horizontal_tile_9_6_to_tile_9_7_2;
	wire horizontal_tile_9_6_to_tile_9_7_3;
	wire horizontal_tile_9_7_to_tile_9_6_0;
	wire horizontal_tile_9_7_to_tile_9_6_1;
	wire horizontal_tile_9_7_to_tile_9_6_2;
	wire horizontal_tile_9_7_to_tile_9_6_3;

	wire horizontal_tile_10_6_to_tile_10_7_0;
	wire horizontal_tile_10_6_to_tile_10_7_1;
	wire horizontal_tile_10_6_to_tile_10_7_2;
	wire horizontal_tile_10_6_to_tile_10_7_3;
	wire horizontal_tile_10_7_to_tile_10_6_0;
	wire horizontal_tile_10_7_to_tile_10_6_1;
	wire horizontal_tile_10_7_to_tile_10_6_2;
	wire horizontal_tile_10_7_to_tile_10_6_3;

	wire horizontal_tile_11_6_to_tile_11_7_0;
	wire horizontal_tile_11_6_to_tile_11_7_1;
	wire horizontal_tile_11_6_to_tile_11_7_2;
	wire horizontal_tile_11_6_to_tile_11_7_3;
	wire horizontal_tile_11_7_to_tile_11_6_0;
	wire horizontal_tile_11_7_to_tile_11_6_1;
	wire horizontal_tile_11_7_to_tile_11_6_2;
	wire horizontal_tile_11_7_to_tile_11_6_3;

	wire horizontal_tile_12_6_to_tile_12_7_0;
	wire horizontal_tile_12_6_to_tile_12_7_1;
	wire horizontal_tile_12_6_to_tile_12_7_2;
	wire horizontal_tile_12_6_to_tile_12_7_3;
	wire horizontal_tile_12_7_to_tile_12_6_0;
	wire horizontal_tile_12_7_to_tile_12_6_1;
	wire horizontal_tile_12_7_to_tile_12_6_2;
	wire horizontal_tile_12_7_to_tile_12_6_3;

	wire horizontal_tile_13_6_to_tile_13_7_0;
	wire horizontal_tile_13_6_to_tile_13_7_1;
	wire horizontal_tile_13_6_to_tile_13_7_2;
	wire horizontal_tile_13_6_to_tile_13_7_3;
	wire horizontal_tile_13_7_to_tile_13_6_0;
	wire horizontal_tile_13_7_to_tile_13_6_1;
	wire horizontal_tile_13_7_to_tile_13_6_2;
	wire horizontal_tile_13_7_to_tile_13_6_3;

	wire horizontal_tile_14_6_to_tile_14_7_0;
	wire horizontal_tile_14_6_to_tile_14_7_1;
	wire horizontal_tile_14_6_to_tile_14_7_2;
	wire horizontal_tile_14_6_to_tile_14_7_3;
	wire horizontal_tile_14_7_to_tile_14_6_0;
	wire horizontal_tile_14_7_to_tile_14_6_1;
	wire horizontal_tile_14_7_to_tile_14_6_2;
	wire horizontal_tile_14_7_to_tile_14_6_3;

	wire horizontal_tile_15_6_to_tile_15_7_0;
	wire horizontal_tile_15_6_to_tile_15_7_1;
	wire horizontal_tile_15_6_to_tile_15_7_2;
	wire horizontal_tile_15_6_to_tile_15_7_3;
	wire horizontal_tile_15_7_to_tile_15_6_0;
	wire horizontal_tile_15_7_to_tile_15_6_1;
	wire horizontal_tile_15_7_to_tile_15_6_2;
	wire horizontal_tile_15_7_to_tile_15_6_3;

	wire horizontal_tile_16_6_to_tile_16_7_0;
	wire horizontal_tile_16_6_to_tile_16_7_1;
	wire horizontal_tile_16_6_to_tile_16_7_2;
	wire horizontal_tile_16_6_to_tile_16_7_3;
	wire horizontal_tile_16_7_to_tile_16_6_0;
	wire horizontal_tile_16_7_to_tile_16_6_1;
	wire horizontal_tile_16_7_to_tile_16_6_2;
	wire horizontal_tile_16_7_to_tile_16_6_3;

	wire horizontal_tile_17_6_to_tile_17_7_0;
	wire horizontal_tile_17_6_to_tile_17_7_1;
	wire horizontal_tile_17_6_to_tile_17_7_2;
	wire horizontal_tile_17_6_to_tile_17_7_3;
	wire horizontal_tile_17_7_to_tile_17_6_0;
	wire horizontal_tile_17_7_to_tile_17_6_1;
	wire horizontal_tile_17_7_to_tile_17_6_2;
	wire horizontal_tile_17_7_to_tile_17_6_3;

	wire horizontal_tile_18_6_to_tile_18_7_0;
	wire horizontal_tile_18_6_to_tile_18_7_1;
	wire horizontal_tile_18_6_to_tile_18_7_2;
	wire horizontal_tile_18_6_to_tile_18_7_3;
	wire horizontal_tile_18_7_to_tile_18_6_0;
	wire horizontal_tile_18_7_to_tile_18_6_1;
	wire horizontal_tile_18_7_to_tile_18_6_2;
	wire horizontal_tile_18_7_to_tile_18_6_3;

	wire horizontal_tile_19_6_to_tile_19_7_0;
	wire horizontal_tile_19_6_to_tile_19_7_1;
	wire horizontal_tile_19_6_to_tile_19_7_2;
	wire horizontal_tile_19_6_to_tile_19_7_3;
	wire horizontal_tile_19_7_to_tile_19_6_0;
	wire horizontal_tile_19_7_to_tile_19_6_1;
	wire horizontal_tile_19_7_to_tile_19_6_2;
	wire horizontal_tile_19_7_to_tile_19_6_3;

	wire horizontal_tile_20_6_to_tile_20_7_0;
	wire horizontal_tile_20_6_to_tile_20_7_1;
	wire horizontal_tile_20_6_to_tile_20_7_2;
	wire horizontal_tile_20_6_to_tile_20_7_3;
	wire horizontal_tile_20_7_to_tile_20_6_0;
	wire horizontal_tile_20_7_to_tile_20_6_1;
	wire horizontal_tile_20_7_to_tile_20_6_2;
	wire horizontal_tile_20_7_to_tile_20_6_3;

	wire horizontal_tile_21_6_to_tile_21_7_0;
	wire horizontal_tile_21_6_to_tile_21_7_1;
	wire horizontal_tile_21_6_to_tile_21_7_2;
	wire horizontal_tile_21_6_to_tile_21_7_3;
	wire horizontal_tile_21_7_to_tile_21_6_0;
	wire horizontal_tile_21_7_to_tile_21_6_1;
	wire horizontal_tile_21_7_to_tile_21_6_2;
	wire horizontal_tile_21_7_to_tile_21_6_3;

	wire horizontal_tile_22_6_to_tile_22_7_0;
	wire horizontal_tile_22_6_to_tile_22_7_1;
	wire horizontal_tile_22_6_to_tile_22_7_2;
	wire horizontal_tile_22_6_to_tile_22_7_3;
	wire horizontal_tile_22_7_to_tile_22_6_0;
	wire horizontal_tile_22_7_to_tile_22_6_1;
	wire horizontal_tile_22_7_to_tile_22_6_2;
	wire horizontal_tile_22_7_to_tile_22_6_3;

	wire horizontal_tile_23_6_to_tile_23_7_0;
	wire horizontal_tile_23_6_to_tile_23_7_1;
	wire horizontal_tile_23_6_to_tile_23_7_2;
	wire horizontal_tile_23_6_to_tile_23_7_3;
	wire horizontal_tile_23_7_to_tile_23_6_0;
	wire horizontal_tile_23_7_to_tile_23_6_1;
	wire horizontal_tile_23_7_to_tile_23_6_2;
	wire horizontal_tile_23_7_to_tile_23_6_3;

	wire horizontal_tile_24_6_to_tile_24_7_0;
	wire horizontal_tile_24_6_to_tile_24_7_1;
	wire horizontal_tile_24_6_to_tile_24_7_2;
	wire horizontal_tile_24_6_to_tile_24_7_3;
	wire horizontal_tile_24_7_to_tile_24_6_0;
	wire horizontal_tile_24_7_to_tile_24_6_1;
	wire horizontal_tile_24_7_to_tile_24_6_2;
	wire horizontal_tile_24_7_to_tile_24_6_3;

	wire horizontal_tile_25_6_to_tile_25_7_0;
	wire horizontal_tile_25_6_to_tile_25_7_1;
	wire horizontal_tile_25_6_to_tile_25_7_2;
	wire horizontal_tile_25_6_to_tile_25_7_3;
	wire horizontal_tile_25_7_to_tile_25_6_0;
	wire horizontal_tile_25_7_to_tile_25_6_1;
	wire horizontal_tile_25_7_to_tile_25_6_2;
	wire horizontal_tile_25_7_to_tile_25_6_3;

	wire horizontal_tile_26_6_to_tile_26_7_0;
	wire horizontal_tile_26_6_to_tile_26_7_1;
	wire horizontal_tile_26_6_to_tile_26_7_2;
	wire horizontal_tile_26_6_to_tile_26_7_3;
	wire horizontal_tile_26_7_to_tile_26_6_0;
	wire horizontal_tile_26_7_to_tile_26_6_1;
	wire horizontal_tile_26_7_to_tile_26_6_2;
	wire horizontal_tile_26_7_to_tile_26_6_3;

	wire horizontal_tile_27_6_to_tile_27_7_0;
	wire horizontal_tile_27_6_to_tile_27_7_1;
	wire horizontal_tile_27_6_to_tile_27_7_2;
	wire horizontal_tile_27_6_to_tile_27_7_3;
	wire horizontal_tile_27_7_to_tile_27_6_0;
	wire horizontal_tile_27_7_to_tile_27_6_1;
	wire horizontal_tile_27_7_to_tile_27_6_2;
	wire horizontal_tile_27_7_to_tile_27_6_3;

	wire horizontal_tile_28_6_to_tile_28_7_0;
	wire horizontal_tile_28_6_to_tile_28_7_1;
	wire horizontal_tile_28_6_to_tile_28_7_2;
	wire horizontal_tile_28_6_to_tile_28_7_3;
	wire horizontal_tile_28_7_to_tile_28_6_0;
	wire horizontal_tile_28_7_to_tile_28_6_1;
	wire horizontal_tile_28_7_to_tile_28_6_2;
	wire horizontal_tile_28_7_to_tile_28_6_3;

	wire horizontal_tile_29_6_to_tile_29_7_0;
	wire horizontal_tile_29_6_to_tile_29_7_1;
	wire horizontal_tile_29_6_to_tile_29_7_2;
	wire horizontal_tile_29_6_to_tile_29_7_3;
	wire horizontal_tile_29_7_to_tile_29_6_0;
	wire horizontal_tile_29_7_to_tile_29_6_1;
	wire horizontal_tile_29_7_to_tile_29_6_2;
	wire horizontal_tile_29_7_to_tile_29_6_3;

	wire horizontal_tile_30_6_to_tile_30_7_0;
	wire horizontal_tile_30_6_to_tile_30_7_1;
	wire horizontal_tile_30_6_to_tile_30_7_2;
	wire horizontal_tile_30_6_to_tile_30_7_3;
	wire horizontal_tile_30_7_to_tile_30_6_0;
	wire horizontal_tile_30_7_to_tile_30_6_1;
	wire horizontal_tile_30_7_to_tile_30_6_2;
	wire horizontal_tile_30_7_to_tile_30_6_3;

	wire horizontal_tile_31_6_to_tile_31_7_0;
	wire horizontal_tile_31_6_to_tile_31_7_1;
	wire horizontal_tile_31_6_to_tile_31_7_2;
	wire horizontal_tile_31_6_to_tile_31_7_3;
	wire horizontal_tile_31_7_to_tile_31_6_0;
	wire horizontal_tile_31_7_to_tile_31_6_1;
	wire horizontal_tile_31_7_to_tile_31_6_2;
	wire horizontal_tile_31_7_to_tile_31_6_3;

	wire horizontal_tile_0_7_to_tile_0_8_0;
	wire horizontal_tile_0_7_to_tile_0_8_1;
	wire horizontal_tile_0_7_to_tile_0_8_2;
	wire horizontal_tile_0_7_to_tile_0_8_3;
	wire horizontal_tile_0_8_to_tile_0_7_0;
	wire horizontal_tile_0_8_to_tile_0_7_1;
	wire horizontal_tile_0_8_to_tile_0_7_2;
	wire horizontal_tile_0_8_to_tile_0_7_3;

	wire horizontal_tile_1_7_to_tile_1_8_0;
	wire horizontal_tile_1_7_to_tile_1_8_1;
	wire horizontal_tile_1_7_to_tile_1_8_2;
	wire horizontal_tile_1_7_to_tile_1_8_3;
	wire horizontal_tile_1_8_to_tile_1_7_0;
	wire horizontal_tile_1_8_to_tile_1_7_1;
	wire horizontal_tile_1_8_to_tile_1_7_2;
	wire horizontal_tile_1_8_to_tile_1_7_3;

	wire horizontal_tile_2_7_to_tile_2_8_0;
	wire horizontal_tile_2_7_to_tile_2_8_1;
	wire horizontal_tile_2_7_to_tile_2_8_2;
	wire horizontal_tile_2_7_to_tile_2_8_3;
	wire horizontal_tile_2_8_to_tile_2_7_0;
	wire horizontal_tile_2_8_to_tile_2_7_1;
	wire horizontal_tile_2_8_to_tile_2_7_2;
	wire horizontal_tile_2_8_to_tile_2_7_3;

	wire horizontal_tile_3_7_to_tile_3_8_0;
	wire horizontal_tile_3_7_to_tile_3_8_1;
	wire horizontal_tile_3_7_to_tile_3_8_2;
	wire horizontal_tile_3_7_to_tile_3_8_3;
	wire horizontal_tile_3_8_to_tile_3_7_0;
	wire horizontal_tile_3_8_to_tile_3_7_1;
	wire horizontal_tile_3_8_to_tile_3_7_2;
	wire horizontal_tile_3_8_to_tile_3_7_3;

	wire horizontal_tile_4_7_to_tile_4_8_0;
	wire horizontal_tile_4_7_to_tile_4_8_1;
	wire horizontal_tile_4_7_to_tile_4_8_2;
	wire horizontal_tile_4_7_to_tile_4_8_3;
	wire horizontal_tile_4_8_to_tile_4_7_0;
	wire horizontal_tile_4_8_to_tile_4_7_1;
	wire horizontal_tile_4_8_to_tile_4_7_2;
	wire horizontal_tile_4_8_to_tile_4_7_3;

	wire horizontal_tile_5_7_to_tile_5_8_0;
	wire horizontal_tile_5_7_to_tile_5_8_1;
	wire horizontal_tile_5_7_to_tile_5_8_2;
	wire horizontal_tile_5_7_to_tile_5_8_3;
	wire horizontal_tile_5_8_to_tile_5_7_0;
	wire horizontal_tile_5_8_to_tile_5_7_1;
	wire horizontal_tile_5_8_to_tile_5_7_2;
	wire horizontal_tile_5_8_to_tile_5_7_3;

	wire horizontal_tile_6_7_to_tile_6_8_0;
	wire horizontal_tile_6_7_to_tile_6_8_1;
	wire horizontal_tile_6_7_to_tile_6_8_2;
	wire horizontal_tile_6_7_to_tile_6_8_3;
	wire horizontal_tile_6_8_to_tile_6_7_0;
	wire horizontal_tile_6_8_to_tile_6_7_1;
	wire horizontal_tile_6_8_to_tile_6_7_2;
	wire horizontal_tile_6_8_to_tile_6_7_3;

	wire horizontal_tile_7_7_to_tile_7_8_0;
	wire horizontal_tile_7_7_to_tile_7_8_1;
	wire horizontal_tile_7_7_to_tile_7_8_2;
	wire horizontal_tile_7_7_to_tile_7_8_3;
	wire horizontal_tile_7_8_to_tile_7_7_0;
	wire horizontal_tile_7_8_to_tile_7_7_1;
	wire horizontal_tile_7_8_to_tile_7_7_2;
	wire horizontal_tile_7_8_to_tile_7_7_3;

	wire horizontal_tile_8_7_to_tile_8_8_0;
	wire horizontal_tile_8_7_to_tile_8_8_1;
	wire horizontal_tile_8_7_to_tile_8_8_2;
	wire horizontal_tile_8_7_to_tile_8_8_3;
	wire horizontal_tile_8_8_to_tile_8_7_0;
	wire horizontal_tile_8_8_to_tile_8_7_1;
	wire horizontal_tile_8_8_to_tile_8_7_2;
	wire horizontal_tile_8_8_to_tile_8_7_3;

	wire horizontal_tile_9_7_to_tile_9_8_0;
	wire horizontal_tile_9_7_to_tile_9_8_1;
	wire horizontal_tile_9_7_to_tile_9_8_2;
	wire horizontal_tile_9_7_to_tile_9_8_3;
	wire horizontal_tile_9_8_to_tile_9_7_0;
	wire horizontal_tile_9_8_to_tile_9_7_1;
	wire horizontal_tile_9_8_to_tile_9_7_2;
	wire horizontal_tile_9_8_to_tile_9_7_3;

	wire horizontal_tile_10_7_to_tile_10_8_0;
	wire horizontal_tile_10_7_to_tile_10_8_1;
	wire horizontal_tile_10_7_to_tile_10_8_2;
	wire horizontal_tile_10_7_to_tile_10_8_3;
	wire horizontal_tile_10_8_to_tile_10_7_0;
	wire horizontal_tile_10_8_to_tile_10_7_1;
	wire horizontal_tile_10_8_to_tile_10_7_2;
	wire horizontal_tile_10_8_to_tile_10_7_3;

	wire horizontal_tile_11_7_to_tile_11_8_0;
	wire horizontal_tile_11_7_to_tile_11_8_1;
	wire horizontal_tile_11_7_to_tile_11_8_2;
	wire horizontal_tile_11_7_to_tile_11_8_3;
	wire horizontal_tile_11_8_to_tile_11_7_0;
	wire horizontal_tile_11_8_to_tile_11_7_1;
	wire horizontal_tile_11_8_to_tile_11_7_2;
	wire horizontal_tile_11_8_to_tile_11_7_3;

	wire horizontal_tile_12_7_to_tile_12_8_0;
	wire horizontal_tile_12_7_to_tile_12_8_1;
	wire horizontal_tile_12_7_to_tile_12_8_2;
	wire horizontal_tile_12_7_to_tile_12_8_3;
	wire horizontal_tile_12_8_to_tile_12_7_0;
	wire horizontal_tile_12_8_to_tile_12_7_1;
	wire horizontal_tile_12_8_to_tile_12_7_2;
	wire horizontal_tile_12_8_to_tile_12_7_3;

	wire horizontal_tile_13_7_to_tile_13_8_0;
	wire horizontal_tile_13_7_to_tile_13_8_1;
	wire horizontal_tile_13_7_to_tile_13_8_2;
	wire horizontal_tile_13_7_to_tile_13_8_3;
	wire horizontal_tile_13_8_to_tile_13_7_0;
	wire horizontal_tile_13_8_to_tile_13_7_1;
	wire horizontal_tile_13_8_to_tile_13_7_2;
	wire horizontal_tile_13_8_to_tile_13_7_3;

	wire horizontal_tile_14_7_to_tile_14_8_0;
	wire horizontal_tile_14_7_to_tile_14_8_1;
	wire horizontal_tile_14_7_to_tile_14_8_2;
	wire horizontal_tile_14_7_to_tile_14_8_3;
	wire horizontal_tile_14_8_to_tile_14_7_0;
	wire horizontal_tile_14_8_to_tile_14_7_1;
	wire horizontal_tile_14_8_to_tile_14_7_2;
	wire horizontal_tile_14_8_to_tile_14_7_3;

	wire horizontal_tile_15_7_to_tile_15_8_0;
	wire horizontal_tile_15_7_to_tile_15_8_1;
	wire horizontal_tile_15_7_to_tile_15_8_2;
	wire horizontal_tile_15_7_to_tile_15_8_3;
	wire horizontal_tile_15_8_to_tile_15_7_0;
	wire horizontal_tile_15_8_to_tile_15_7_1;
	wire horizontal_tile_15_8_to_tile_15_7_2;
	wire horizontal_tile_15_8_to_tile_15_7_3;

	wire horizontal_tile_16_7_to_tile_16_8_0;
	wire horizontal_tile_16_7_to_tile_16_8_1;
	wire horizontal_tile_16_7_to_tile_16_8_2;
	wire horizontal_tile_16_7_to_tile_16_8_3;
	wire horizontal_tile_16_8_to_tile_16_7_0;
	wire horizontal_tile_16_8_to_tile_16_7_1;
	wire horizontal_tile_16_8_to_tile_16_7_2;
	wire horizontal_tile_16_8_to_tile_16_7_3;

	wire horizontal_tile_17_7_to_tile_17_8_0;
	wire horizontal_tile_17_7_to_tile_17_8_1;
	wire horizontal_tile_17_7_to_tile_17_8_2;
	wire horizontal_tile_17_7_to_tile_17_8_3;
	wire horizontal_tile_17_8_to_tile_17_7_0;
	wire horizontal_tile_17_8_to_tile_17_7_1;
	wire horizontal_tile_17_8_to_tile_17_7_2;
	wire horizontal_tile_17_8_to_tile_17_7_3;

	wire horizontal_tile_18_7_to_tile_18_8_0;
	wire horizontal_tile_18_7_to_tile_18_8_1;
	wire horizontal_tile_18_7_to_tile_18_8_2;
	wire horizontal_tile_18_7_to_tile_18_8_3;
	wire horizontal_tile_18_8_to_tile_18_7_0;
	wire horizontal_tile_18_8_to_tile_18_7_1;
	wire horizontal_tile_18_8_to_tile_18_7_2;
	wire horizontal_tile_18_8_to_tile_18_7_3;

	wire horizontal_tile_19_7_to_tile_19_8_0;
	wire horizontal_tile_19_7_to_tile_19_8_1;
	wire horizontal_tile_19_7_to_tile_19_8_2;
	wire horizontal_tile_19_7_to_tile_19_8_3;
	wire horizontal_tile_19_8_to_tile_19_7_0;
	wire horizontal_tile_19_8_to_tile_19_7_1;
	wire horizontal_tile_19_8_to_tile_19_7_2;
	wire horizontal_tile_19_8_to_tile_19_7_3;

	wire horizontal_tile_20_7_to_tile_20_8_0;
	wire horizontal_tile_20_7_to_tile_20_8_1;
	wire horizontal_tile_20_7_to_tile_20_8_2;
	wire horizontal_tile_20_7_to_tile_20_8_3;
	wire horizontal_tile_20_8_to_tile_20_7_0;
	wire horizontal_tile_20_8_to_tile_20_7_1;
	wire horizontal_tile_20_8_to_tile_20_7_2;
	wire horizontal_tile_20_8_to_tile_20_7_3;

	wire horizontal_tile_21_7_to_tile_21_8_0;
	wire horizontal_tile_21_7_to_tile_21_8_1;
	wire horizontal_tile_21_7_to_tile_21_8_2;
	wire horizontal_tile_21_7_to_tile_21_8_3;
	wire horizontal_tile_21_8_to_tile_21_7_0;
	wire horizontal_tile_21_8_to_tile_21_7_1;
	wire horizontal_tile_21_8_to_tile_21_7_2;
	wire horizontal_tile_21_8_to_tile_21_7_3;

	wire horizontal_tile_22_7_to_tile_22_8_0;
	wire horizontal_tile_22_7_to_tile_22_8_1;
	wire horizontal_tile_22_7_to_tile_22_8_2;
	wire horizontal_tile_22_7_to_tile_22_8_3;
	wire horizontal_tile_22_8_to_tile_22_7_0;
	wire horizontal_tile_22_8_to_tile_22_7_1;
	wire horizontal_tile_22_8_to_tile_22_7_2;
	wire horizontal_tile_22_8_to_tile_22_7_3;

	wire horizontal_tile_23_7_to_tile_23_8_0;
	wire horizontal_tile_23_7_to_tile_23_8_1;
	wire horizontal_tile_23_7_to_tile_23_8_2;
	wire horizontal_tile_23_7_to_tile_23_8_3;
	wire horizontal_tile_23_8_to_tile_23_7_0;
	wire horizontal_tile_23_8_to_tile_23_7_1;
	wire horizontal_tile_23_8_to_tile_23_7_2;
	wire horizontal_tile_23_8_to_tile_23_7_3;

	wire horizontal_tile_24_7_to_tile_24_8_0;
	wire horizontal_tile_24_7_to_tile_24_8_1;
	wire horizontal_tile_24_7_to_tile_24_8_2;
	wire horizontal_tile_24_7_to_tile_24_8_3;
	wire horizontal_tile_24_8_to_tile_24_7_0;
	wire horizontal_tile_24_8_to_tile_24_7_1;
	wire horizontal_tile_24_8_to_tile_24_7_2;
	wire horizontal_tile_24_8_to_tile_24_7_3;

	wire horizontal_tile_25_7_to_tile_25_8_0;
	wire horizontal_tile_25_7_to_tile_25_8_1;
	wire horizontal_tile_25_7_to_tile_25_8_2;
	wire horizontal_tile_25_7_to_tile_25_8_3;
	wire horizontal_tile_25_8_to_tile_25_7_0;
	wire horizontal_tile_25_8_to_tile_25_7_1;
	wire horizontal_tile_25_8_to_tile_25_7_2;
	wire horizontal_tile_25_8_to_tile_25_7_3;

	wire horizontal_tile_26_7_to_tile_26_8_0;
	wire horizontal_tile_26_7_to_tile_26_8_1;
	wire horizontal_tile_26_7_to_tile_26_8_2;
	wire horizontal_tile_26_7_to_tile_26_8_3;
	wire horizontal_tile_26_8_to_tile_26_7_0;
	wire horizontal_tile_26_8_to_tile_26_7_1;
	wire horizontal_tile_26_8_to_tile_26_7_2;
	wire horizontal_tile_26_8_to_tile_26_7_3;

	wire horizontal_tile_27_7_to_tile_27_8_0;
	wire horizontal_tile_27_7_to_tile_27_8_1;
	wire horizontal_tile_27_7_to_tile_27_8_2;
	wire horizontal_tile_27_7_to_tile_27_8_3;
	wire horizontal_tile_27_8_to_tile_27_7_0;
	wire horizontal_tile_27_8_to_tile_27_7_1;
	wire horizontal_tile_27_8_to_tile_27_7_2;
	wire horizontal_tile_27_8_to_tile_27_7_3;

	wire horizontal_tile_28_7_to_tile_28_8_0;
	wire horizontal_tile_28_7_to_tile_28_8_1;
	wire horizontal_tile_28_7_to_tile_28_8_2;
	wire horizontal_tile_28_7_to_tile_28_8_3;
	wire horizontal_tile_28_8_to_tile_28_7_0;
	wire horizontal_tile_28_8_to_tile_28_7_1;
	wire horizontal_tile_28_8_to_tile_28_7_2;
	wire horizontal_tile_28_8_to_tile_28_7_3;

	wire horizontal_tile_29_7_to_tile_29_8_0;
	wire horizontal_tile_29_7_to_tile_29_8_1;
	wire horizontal_tile_29_7_to_tile_29_8_2;
	wire horizontal_tile_29_7_to_tile_29_8_3;
	wire horizontal_tile_29_8_to_tile_29_7_0;
	wire horizontal_tile_29_8_to_tile_29_7_1;
	wire horizontal_tile_29_8_to_tile_29_7_2;
	wire horizontal_tile_29_8_to_tile_29_7_3;

	wire horizontal_tile_30_7_to_tile_30_8_0;
	wire horizontal_tile_30_7_to_tile_30_8_1;
	wire horizontal_tile_30_7_to_tile_30_8_2;
	wire horizontal_tile_30_7_to_tile_30_8_3;
	wire horizontal_tile_30_8_to_tile_30_7_0;
	wire horizontal_tile_30_8_to_tile_30_7_1;
	wire horizontal_tile_30_8_to_tile_30_7_2;
	wire horizontal_tile_30_8_to_tile_30_7_3;

	wire horizontal_tile_31_7_to_tile_31_8_0;
	wire horizontal_tile_31_7_to_tile_31_8_1;
	wire horizontal_tile_31_7_to_tile_31_8_2;
	wire horizontal_tile_31_7_to_tile_31_8_3;
	wire horizontal_tile_31_8_to_tile_31_7_0;
	wire horizontal_tile_31_8_to_tile_31_7_1;
	wire horizontal_tile_31_8_to_tile_31_7_2;
	wire horizontal_tile_31_8_to_tile_31_7_3;

	wire horizontal_tile_0_8_to_tile_0_9_0;
	wire horizontal_tile_0_8_to_tile_0_9_1;
	wire horizontal_tile_0_8_to_tile_0_9_2;
	wire horizontal_tile_0_8_to_tile_0_9_3;
	wire horizontal_tile_0_9_to_tile_0_8_0;
	wire horizontal_tile_0_9_to_tile_0_8_1;
	wire horizontal_tile_0_9_to_tile_0_8_2;
	wire horizontal_tile_0_9_to_tile_0_8_3;

	wire horizontal_tile_1_8_to_tile_1_9_0;
	wire horizontal_tile_1_8_to_tile_1_9_1;
	wire horizontal_tile_1_8_to_tile_1_9_2;
	wire horizontal_tile_1_8_to_tile_1_9_3;
	wire horizontal_tile_1_9_to_tile_1_8_0;
	wire horizontal_tile_1_9_to_tile_1_8_1;
	wire horizontal_tile_1_9_to_tile_1_8_2;
	wire horizontal_tile_1_9_to_tile_1_8_3;

	wire horizontal_tile_2_8_to_tile_2_9_0;
	wire horizontal_tile_2_8_to_tile_2_9_1;
	wire horizontal_tile_2_8_to_tile_2_9_2;
	wire horizontal_tile_2_8_to_tile_2_9_3;
	wire horizontal_tile_2_9_to_tile_2_8_0;
	wire horizontal_tile_2_9_to_tile_2_8_1;
	wire horizontal_tile_2_9_to_tile_2_8_2;
	wire horizontal_tile_2_9_to_tile_2_8_3;

	wire horizontal_tile_3_8_to_tile_3_9_0;
	wire horizontal_tile_3_8_to_tile_3_9_1;
	wire horizontal_tile_3_8_to_tile_3_9_2;
	wire horizontal_tile_3_8_to_tile_3_9_3;
	wire horizontal_tile_3_9_to_tile_3_8_0;
	wire horizontal_tile_3_9_to_tile_3_8_1;
	wire horizontal_tile_3_9_to_tile_3_8_2;
	wire horizontal_tile_3_9_to_tile_3_8_3;

	wire horizontal_tile_4_8_to_tile_4_9_0;
	wire horizontal_tile_4_8_to_tile_4_9_1;
	wire horizontal_tile_4_8_to_tile_4_9_2;
	wire horizontal_tile_4_8_to_tile_4_9_3;
	wire horizontal_tile_4_9_to_tile_4_8_0;
	wire horizontal_tile_4_9_to_tile_4_8_1;
	wire horizontal_tile_4_9_to_tile_4_8_2;
	wire horizontal_tile_4_9_to_tile_4_8_3;

	wire horizontal_tile_5_8_to_tile_5_9_0;
	wire horizontal_tile_5_8_to_tile_5_9_1;
	wire horizontal_tile_5_8_to_tile_5_9_2;
	wire horizontal_tile_5_8_to_tile_5_9_3;
	wire horizontal_tile_5_9_to_tile_5_8_0;
	wire horizontal_tile_5_9_to_tile_5_8_1;
	wire horizontal_tile_5_9_to_tile_5_8_2;
	wire horizontal_tile_5_9_to_tile_5_8_3;

	wire horizontal_tile_6_8_to_tile_6_9_0;
	wire horizontal_tile_6_8_to_tile_6_9_1;
	wire horizontal_tile_6_8_to_tile_6_9_2;
	wire horizontal_tile_6_8_to_tile_6_9_3;
	wire horizontal_tile_6_9_to_tile_6_8_0;
	wire horizontal_tile_6_9_to_tile_6_8_1;
	wire horizontal_tile_6_9_to_tile_6_8_2;
	wire horizontal_tile_6_9_to_tile_6_8_3;

	wire horizontal_tile_7_8_to_tile_7_9_0;
	wire horizontal_tile_7_8_to_tile_7_9_1;
	wire horizontal_tile_7_8_to_tile_7_9_2;
	wire horizontal_tile_7_8_to_tile_7_9_3;
	wire horizontal_tile_7_9_to_tile_7_8_0;
	wire horizontal_tile_7_9_to_tile_7_8_1;
	wire horizontal_tile_7_9_to_tile_7_8_2;
	wire horizontal_tile_7_9_to_tile_7_8_3;

	wire horizontal_tile_8_8_to_tile_8_9_0;
	wire horizontal_tile_8_8_to_tile_8_9_1;
	wire horizontal_tile_8_8_to_tile_8_9_2;
	wire horizontal_tile_8_8_to_tile_8_9_3;
	wire horizontal_tile_8_9_to_tile_8_8_0;
	wire horizontal_tile_8_9_to_tile_8_8_1;
	wire horizontal_tile_8_9_to_tile_8_8_2;
	wire horizontal_tile_8_9_to_tile_8_8_3;

	wire horizontal_tile_9_8_to_tile_9_9_0;
	wire horizontal_tile_9_8_to_tile_9_9_1;
	wire horizontal_tile_9_8_to_tile_9_9_2;
	wire horizontal_tile_9_8_to_tile_9_9_3;
	wire horizontal_tile_9_9_to_tile_9_8_0;
	wire horizontal_tile_9_9_to_tile_9_8_1;
	wire horizontal_tile_9_9_to_tile_9_8_2;
	wire horizontal_tile_9_9_to_tile_9_8_3;

	wire horizontal_tile_10_8_to_tile_10_9_0;
	wire horizontal_tile_10_8_to_tile_10_9_1;
	wire horizontal_tile_10_8_to_tile_10_9_2;
	wire horizontal_tile_10_8_to_tile_10_9_3;
	wire horizontal_tile_10_9_to_tile_10_8_0;
	wire horizontal_tile_10_9_to_tile_10_8_1;
	wire horizontal_tile_10_9_to_tile_10_8_2;
	wire horizontal_tile_10_9_to_tile_10_8_3;

	wire horizontal_tile_11_8_to_tile_11_9_0;
	wire horizontal_tile_11_8_to_tile_11_9_1;
	wire horizontal_tile_11_8_to_tile_11_9_2;
	wire horizontal_tile_11_8_to_tile_11_9_3;
	wire horizontal_tile_11_9_to_tile_11_8_0;
	wire horizontal_tile_11_9_to_tile_11_8_1;
	wire horizontal_tile_11_9_to_tile_11_8_2;
	wire horizontal_tile_11_9_to_tile_11_8_3;

	wire horizontal_tile_12_8_to_tile_12_9_0;
	wire horizontal_tile_12_8_to_tile_12_9_1;
	wire horizontal_tile_12_8_to_tile_12_9_2;
	wire horizontal_tile_12_8_to_tile_12_9_3;
	wire horizontal_tile_12_9_to_tile_12_8_0;
	wire horizontal_tile_12_9_to_tile_12_8_1;
	wire horizontal_tile_12_9_to_tile_12_8_2;
	wire horizontal_tile_12_9_to_tile_12_8_3;

	wire horizontal_tile_13_8_to_tile_13_9_0;
	wire horizontal_tile_13_8_to_tile_13_9_1;
	wire horizontal_tile_13_8_to_tile_13_9_2;
	wire horizontal_tile_13_8_to_tile_13_9_3;
	wire horizontal_tile_13_9_to_tile_13_8_0;
	wire horizontal_tile_13_9_to_tile_13_8_1;
	wire horizontal_tile_13_9_to_tile_13_8_2;
	wire horizontal_tile_13_9_to_tile_13_8_3;

	wire horizontal_tile_14_8_to_tile_14_9_0;
	wire horizontal_tile_14_8_to_tile_14_9_1;
	wire horizontal_tile_14_8_to_tile_14_9_2;
	wire horizontal_tile_14_8_to_tile_14_9_3;
	wire horizontal_tile_14_9_to_tile_14_8_0;
	wire horizontal_tile_14_9_to_tile_14_8_1;
	wire horizontal_tile_14_9_to_tile_14_8_2;
	wire horizontal_tile_14_9_to_tile_14_8_3;

	wire horizontal_tile_15_8_to_tile_15_9_0;
	wire horizontal_tile_15_8_to_tile_15_9_1;
	wire horizontal_tile_15_8_to_tile_15_9_2;
	wire horizontal_tile_15_8_to_tile_15_9_3;
	wire horizontal_tile_15_9_to_tile_15_8_0;
	wire horizontal_tile_15_9_to_tile_15_8_1;
	wire horizontal_tile_15_9_to_tile_15_8_2;
	wire horizontal_tile_15_9_to_tile_15_8_3;

	wire horizontal_tile_16_8_to_tile_16_9_0;
	wire horizontal_tile_16_8_to_tile_16_9_1;
	wire horizontal_tile_16_8_to_tile_16_9_2;
	wire horizontal_tile_16_8_to_tile_16_9_3;
	wire horizontal_tile_16_9_to_tile_16_8_0;
	wire horizontal_tile_16_9_to_tile_16_8_1;
	wire horizontal_tile_16_9_to_tile_16_8_2;
	wire horizontal_tile_16_9_to_tile_16_8_3;

	wire horizontal_tile_17_8_to_tile_17_9_0;
	wire horizontal_tile_17_8_to_tile_17_9_1;
	wire horizontal_tile_17_8_to_tile_17_9_2;
	wire horizontal_tile_17_8_to_tile_17_9_3;
	wire horizontal_tile_17_9_to_tile_17_8_0;
	wire horizontal_tile_17_9_to_tile_17_8_1;
	wire horizontal_tile_17_9_to_tile_17_8_2;
	wire horizontal_tile_17_9_to_tile_17_8_3;

	wire horizontal_tile_18_8_to_tile_18_9_0;
	wire horizontal_tile_18_8_to_tile_18_9_1;
	wire horizontal_tile_18_8_to_tile_18_9_2;
	wire horizontal_tile_18_8_to_tile_18_9_3;
	wire horizontal_tile_18_9_to_tile_18_8_0;
	wire horizontal_tile_18_9_to_tile_18_8_1;
	wire horizontal_tile_18_9_to_tile_18_8_2;
	wire horizontal_tile_18_9_to_tile_18_8_3;

	wire horizontal_tile_19_8_to_tile_19_9_0;
	wire horizontal_tile_19_8_to_tile_19_9_1;
	wire horizontal_tile_19_8_to_tile_19_9_2;
	wire horizontal_tile_19_8_to_tile_19_9_3;
	wire horizontal_tile_19_9_to_tile_19_8_0;
	wire horizontal_tile_19_9_to_tile_19_8_1;
	wire horizontal_tile_19_9_to_tile_19_8_2;
	wire horizontal_tile_19_9_to_tile_19_8_3;

	wire horizontal_tile_20_8_to_tile_20_9_0;
	wire horizontal_tile_20_8_to_tile_20_9_1;
	wire horizontal_tile_20_8_to_tile_20_9_2;
	wire horizontal_tile_20_8_to_tile_20_9_3;
	wire horizontal_tile_20_9_to_tile_20_8_0;
	wire horizontal_tile_20_9_to_tile_20_8_1;
	wire horizontal_tile_20_9_to_tile_20_8_2;
	wire horizontal_tile_20_9_to_tile_20_8_3;

	wire horizontal_tile_21_8_to_tile_21_9_0;
	wire horizontal_tile_21_8_to_tile_21_9_1;
	wire horizontal_tile_21_8_to_tile_21_9_2;
	wire horizontal_tile_21_8_to_tile_21_9_3;
	wire horizontal_tile_21_9_to_tile_21_8_0;
	wire horizontal_tile_21_9_to_tile_21_8_1;
	wire horizontal_tile_21_9_to_tile_21_8_2;
	wire horizontal_tile_21_9_to_tile_21_8_3;

	wire horizontal_tile_22_8_to_tile_22_9_0;
	wire horizontal_tile_22_8_to_tile_22_9_1;
	wire horizontal_tile_22_8_to_tile_22_9_2;
	wire horizontal_tile_22_8_to_tile_22_9_3;
	wire horizontal_tile_22_9_to_tile_22_8_0;
	wire horizontal_tile_22_9_to_tile_22_8_1;
	wire horizontal_tile_22_9_to_tile_22_8_2;
	wire horizontal_tile_22_9_to_tile_22_8_3;

	wire horizontal_tile_23_8_to_tile_23_9_0;
	wire horizontal_tile_23_8_to_tile_23_9_1;
	wire horizontal_tile_23_8_to_tile_23_9_2;
	wire horizontal_tile_23_8_to_tile_23_9_3;
	wire horizontal_tile_23_9_to_tile_23_8_0;
	wire horizontal_tile_23_9_to_tile_23_8_1;
	wire horizontal_tile_23_9_to_tile_23_8_2;
	wire horizontal_tile_23_9_to_tile_23_8_3;

	wire horizontal_tile_24_8_to_tile_24_9_0;
	wire horizontal_tile_24_8_to_tile_24_9_1;
	wire horizontal_tile_24_8_to_tile_24_9_2;
	wire horizontal_tile_24_8_to_tile_24_9_3;
	wire horizontal_tile_24_9_to_tile_24_8_0;
	wire horizontal_tile_24_9_to_tile_24_8_1;
	wire horizontal_tile_24_9_to_tile_24_8_2;
	wire horizontal_tile_24_9_to_tile_24_8_3;

	wire horizontal_tile_25_8_to_tile_25_9_0;
	wire horizontal_tile_25_8_to_tile_25_9_1;
	wire horizontal_tile_25_8_to_tile_25_9_2;
	wire horizontal_tile_25_8_to_tile_25_9_3;
	wire horizontal_tile_25_9_to_tile_25_8_0;
	wire horizontal_tile_25_9_to_tile_25_8_1;
	wire horizontal_tile_25_9_to_tile_25_8_2;
	wire horizontal_tile_25_9_to_tile_25_8_3;

	wire horizontal_tile_26_8_to_tile_26_9_0;
	wire horizontal_tile_26_8_to_tile_26_9_1;
	wire horizontal_tile_26_8_to_tile_26_9_2;
	wire horizontal_tile_26_8_to_tile_26_9_3;
	wire horizontal_tile_26_9_to_tile_26_8_0;
	wire horizontal_tile_26_9_to_tile_26_8_1;
	wire horizontal_tile_26_9_to_tile_26_8_2;
	wire horizontal_tile_26_9_to_tile_26_8_3;

	wire horizontal_tile_27_8_to_tile_27_9_0;
	wire horizontal_tile_27_8_to_tile_27_9_1;
	wire horizontal_tile_27_8_to_tile_27_9_2;
	wire horizontal_tile_27_8_to_tile_27_9_3;
	wire horizontal_tile_27_9_to_tile_27_8_0;
	wire horizontal_tile_27_9_to_tile_27_8_1;
	wire horizontal_tile_27_9_to_tile_27_8_2;
	wire horizontal_tile_27_9_to_tile_27_8_3;

	wire horizontal_tile_28_8_to_tile_28_9_0;
	wire horizontal_tile_28_8_to_tile_28_9_1;
	wire horizontal_tile_28_8_to_tile_28_9_2;
	wire horizontal_tile_28_8_to_tile_28_9_3;
	wire horizontal_tile_28_9_to_tile_28_8_0;
	wire horizontal_tile_28_9_to_tile_28_8_1;
	wire horizontal_tile_28_9_to_tile_28_8_2;
	wire horizontal_tile_28_9_to_tile_28_8_3;

	wire horizontal_tile_29_8_to_tile_29_9_0;
	wire horizontal_tile_29_8_to_tile_29_9_1;
	wire horizontal_tile_29_8_to_tile_29_9_2;
	wire horizontal_tile_29_8_to_tile_29_9_3;
	wire horizontal_tile_29_9_to_tile_29_8_0;
	wire horizontal_tile_29_9_to_tile_29_8_1;
	wire horizontal_tile_29_9_to_tile_29_8_2;
	wire horizontal_tile_29_9_to_tile_29_8_3;

	wire horizontal_tile_30_8_to_tile_30_9_0;
	wire horizontal_tile_30_8_to_tile_30_9_1;
	wire horizontal_tile_30_8_to_tile_30_9_2;
	wire horizontal_tile_30_8_to_tile_30_9_3;
	wire horizontal_tile_30_9_to_tile_30_8_0;
	wire horizontal_tile_30_9_to_tile_30_8_1;
	wire horizontal_tile_30_9_to_tile_30_8_2;
	wire horizontal_tile_30_9_to_tile_30_8_3;

	wire horizontal_tile_31_8_to_tile_31_9_0;
	wire horizontal_tile_31_8_to_tile_31_9_1;
	wire horizontal_tile_31_8_to_tile_31_9_2;
	wire horizontal_tile_31_8_to_tile_31_9_3;
	wire horizontal_tile_31_9_to_tile_31_8_0;
	wire horizontal_tile_31_9_to_tile_31_8_1;
	wire horizontal_tile_31_9_to_tile_31_8_2;
	wire horizontal_tile_31_9_to_tile_31_8_3;

	wire horizontal_tile_0_9_to_tile_0_10_0;
	wire horizontal_tile_0_9_to_tile_0_10_1;
	wire horizontal_tile_0_9_to_tile_0_10_2;
	wire horizontal_tile_0_9_to_tile_0_10_3;
	wire horizontal_tile_0_10_to_tile_0_9_0;
	wire horizontal_tile_0_10_to_tile_0_9_1;
	wire horizontal_tile_0_10_to_tile_0_9_2;
	wire horizontal_tile_0_10_to_tile_0_9_3;

	wire horizontal_tile_1_9_to_tile_1_10_0;
	wire horizontal_tile_1_9_to_tile_1_10_1;
	wire horizontal_tile_1_9_to_tile_1_10_2;
	wire horizontal_tile_1_9_to_tile_1_10_3;
	wire horizontal_tile_1_10_to_tile_1_9_0;
	wire horizontal_tile_1_10_to_tile_1_9_1;
	wire horizontal_tile_1_10_to_tile_1_9_2;
	wire horizontal_tile_1_10_to_tile_1_9_3;

	wire horizontal_tile_2_9_to_tile_2_10_0;
	wire horizontal_tile_2_9_to_tile_2_10_1;
	wire horizontal_tile_2_9_to_tile_2_10_2;
	wire horizontal_tile_2_9_to_tile_2_10_3;
	wire horizontal_tile_2_10_to_tile_2_9_0;
	wire horizontal_tile_2_10_to_tile_2_9_1;
	wire horizontal_tile_2_10_to_tile_2_9_2;
	wire horizontal_tile_2_10_to_tile_2_9_3;

	wire horizontal_tile_3_9_to_tile_3_10_0;
	wire horizontal_tile_3_9_to_tile_3_10_1;
	wire horizontal_tile_3_9_to_tile_3_10_2;
	wire horizontal_tile_3_9_to_tile_3_10_3;
	wire horizontal_tile_3_10_to_tile_3_9_0;
	wire horizontal_tile_3_10_to_tile_3_9_1;
	wire horizontal_tile_3_10_to_tile_3_9_2;
	wire horizontal_tile_3_10_to_tile_3_9_3;

	wire horizontal_tile_4_9_to_tile_4_10_0;
	wire horizontal_tile_4_9_to_tile_4_10_1;
	wire horizontal_tile_4_9_to_tile_4_10_2;
	wire horizontal_tile_4_9_to_tile_4_10_3;
	wire horizontal_tile_4_10_to_tile_4_9_0;
	wire horizontal_tile_4_10_to_tile_4_9_1;
	wire horizontal_tile_4_10_to_tile_4_9_2;
	wire horizontal_tile_4_10_to_tile_4_9_3;

	wire horizontal_tile_5_9_to_tile_5_10_0;
	wire horizontal_tile_5_9_to_tile_5_10_1;
	wire horizontal_tile_5_9_to_tile_5_10_2;
	wire horizontal_tile_5_9_to_tile_5_10_3;
	wire horizontal_tile_5_10_to_tile_5_9_0;
	wire horizontal_tile_5_10_to_tile_5_9_1;
	wire horizontal_tile_5_10_to_tile_5_9_2;
	wire horizontal_tile_5_10_to_tile_5_9_3;

	wire horizontal_tile_6_9_to_tile_6_10_0;
	wire horizontal_tile_6_9_to_tile_6_10_1;
	wire horizontal_tile_6_9_to_tile_6_10_2;
	wire horizontal_tile_6_9_to_tile_6_10_3;
	wire horizontal_tile_6_10_to_tile_6_9_0;
	wire horizontal_tile_6_10_to_tile_6_9_1;
	wire horizontal_tile_6_10_to_tile_6_9_2;
	wire horizontal_tile_6_10_to_tile_6_9_3;

	wire horizontal_tile_7_9_to_tile_7_10_0;
	wire horizontal_tile_7_9_to_tile_7_10_1;
	wire horizontal_tile_7_9_to_tile_7_10_2;
	wire horizontal_tile_7_9_to_tile_7_10_3;
	wire horizontal_tile_7_10_to_tile_7_9_0;
	wire horizontal_tile_7_10_to_tile_7_9_1;
	wire horizontal_tile_7_10_to_tile_7_9_2;
	wire horizontal_tile_7_10_to_tile_7_9_3;

	wire horizontal_tile_8_9_to_tile_8_10_0;
	wire horizontal_tile_8_9_to_tile_8_10_1;
	wire horizontal_tile_8_9_to_tile_8_10_2;
	wire horizontal_tile_8_9_to_tile_8_10_3;
	wire horizontal_tile_8_10_to_tile_8_9_0;
	wire horizontal_tile_8_10_to_tile_8_9_1;
	wire horizontal_tile_8_10_to_tile_8_9_2;
	wire horizontal_tile_8_10_to_tile_8_9_3;

	wire horizontal_tile_9_9_to_tile_9_10_0;
	wire horizontal_tile_9_9_to_tile_9_10_1;
	wire horizontal_tile_9_9_to_tile_9_10_2;
	wire horizontal_tile_9_9_to_tile_9_10_3;
	wire horizontal_tile_9_10_to_tile_9_9_0;
	wire horizontal_tile_9_10_to_tile_9_9_1;
	wire horizontal_tile_9_10_to_tile_9_9_2;
	wire horizontal_tile_9_10_to_tile_9_9_3;

	wire horizontal_tile_10_9_to_tile_10_10_0;
	wire horizontal_tile_10_9_to_tile_10_10_1;
	wire horizontal_tile_10_9_to_tile_10_10_2;
	wire horizontal_tile_10_9_to_tile_10_10_3;
	wire horizontal_tile_10_10_to_tile_10_9_0;
	wire horizontal_tile_10_10_to_tile_10_9_1;
	wire horizontal_tile_10_10_to_tile_10_9_2;
	wire horizontal_tile_10_10_to_tile_10_9_3;

	wire horizontal_tile_11_9_to_tile_11_10_0;
	wire horizontal_tile_11_9_to_tile_11_10_1;
	wire horizontal_tile_11_9_to_tile_11_10_2;
	wire horizontal_tile_11_9_to_tile_11_10_3;
	wire horizontal_tile_11_10_to_tile_11_9_0;
	wire horizontal_tile_11_10_to_tile_11_9_1;
	wire horizontal_tile_11_10_to_tile_11_9_2;
	wire horizontal_tile_11_10_to_tile_11_9_3;

	wire horizontal_tile_12_9_to_tile_12_10_0;
	wire horizontal_tile_12_9_to_tile_12_10_1;
	wire horizontal_tile_12_9_to_tile_12_10_2;
	wire horizontal_tile_12_9_to_tile_12_10_3;
	wire horizontal_tile_12_10_to_tile_12_9_0;
	wire horizontal_tile_12_10_to_tile_12_9_1;
	wire horizontal_tile_12_10_to_tile_12_9_2;
	wire horizontal_tile_12_10_to_tile_12_9_3;

	wire horizontal_tile_13_9_to_tile_13_10_0;
	wire horizontal_tile_13_9_to_tile_13_10_1;
	wire horizontal_tile_13_9_to_tile_13_10_2;
	wire horizontal_tile_13_9_to_tile_13_10_3;
	wire horizontal_tile_13_10_to_tile_13_9_0;
	wire horizontal_tile_13_10_to_tile_13_9_1;
	wire horizontal_tile_13_10_to_tile_13_9_2;
	wire horizontal_tile_13_10_to_tile_13_9_3;

	wire horizontal_tile_14_9_to_tile_14_10_0;
	wire horizontal_tile_14_9_to_tile_14_10_1;
	wire horizontal_tile_14_9_to_tile_14_10_2;
	wire horizontal_tile_14_9_to_tile_14_10_3;
	wire horizontal_tile_14_10_to_tile_14_9_0;
	wire horizontal_tile_14_10_to_tile_14_9_1;
	wire horizontal_tile_14_10_to_tile_14_9_2;
	wire horizontal_tile_14_10_to_tile_14_9_3;

	wire horizontal_tile_15_9_to_tile_15_10_0;
	wire horizontal_tile_15_9_to_tile_15_10_1;
	wire horizontal_tile_15_9_to_tile_15_10_2;
	wire horizontal_tile_15_9_to_tile_15_10_3;
	wire horizontal_tile_15_10_to_tile_15_9_0;
	wire horizontal_tile_15_10_to_tile_15_9_1;
	wire horizontal_tile_15_10_to_tile_15_9_2;
	wire horizontal_tile_15_10_to_tile_15_9_3;

	wire horizontal_tile_16_9_to_tile_16_10_0;
	wire horizontal_tile_16_9_to_tile_16_10_1;
	wire horizontal_tile_16_9_to_tile_16_10_2;
	wire horizontal_tile_16_9_to_tile_16_10_3;
	wire horizontal_tile_16_10_to_tile_16_9_0;
	wire horizontal_tile_16_10_to_tile_16_9_1;
	wire horizontal_tile_16_10_to_tile_16_9_2;
	wire horizontal_tile_16_10_to_tile_16_9_3;

	wire horizontal_tile_17_9_to_tile_17_10_0;
	wire horizontal_tile_17_9_to_tile_17_10_1;
	wire horizontal_tile_17_9_to_tile_17_10_2;
	wire horizontal_tile_17_9_to_tile_17_10_3;
	wire horizontal_tile_17_10_to_tile_17_9_0;
	wire horizontal_tile_17_10_to_tile_17_9_1;
	wire horizontal_tile_17_10_to_tile_17_9_2;
	wire horizontal_tile_17_10_to_tile_17_9_3;

	wire horizontal_tile_18_9_to_tile_18_10_0;
	wire horizontal_tile_18_9_to_tile_18_10_1;
	wire horizontal_tile_18_9_to_tile_18_10_2;
	wire horizontal_tile_18_9_to_tile_18_10_3;
	wire horizontal_tile_18_10_to_tile_18_9_0;
	wire horizontal_tile_18_10_to_tile_18_9_1;
	wire horizontal_tile_18_10_to_tile_18_9_2;
	wire horizontal_tile_18_10_to_tile_18_9_3;

	wire horizontal_tile_19_9_to_tile_19_10_0;
	wire horizontal_tile_19_9_to_tile_19_10_1;
	wire horizontal_tile_19_9_to_tile_19_10_2;
	wire horizontal_tile_19_9_to_tile_19_10_3;
	wire horizontal_tile_19_10_to_tile_19_9_0;
	wire horizontal_tile_19_10_to_tile_19_9_1;
	wire horizontal_tile_19_10_to_tile_19_9_2;
	wire horizontal_tile_19_10_to_tile_19_9_3;

	wire horizontal_tile_20_9_to_tile_20_10_0;
	wire horizontal_tile_20_9_to_tile_20_10_1;
	wire horizontal_tile_20_9_to_tile_20_10_2;
	wire horizontal_tile_20_9_to_tile_20_10_3;
	wire horizontal_tile_20_10_to_tile_20_9_0;
	wire horizontal_tile_20_10_to_tile_20_9_1;
	wire horizontal_tile_20_10_to_tile_20_9_2;
	wire horizontal_tile_20_10_to_tile_20_9_3;

	wire horizontal_tile_21_9_to_tile_21_10_0;
	wire horizontal_tile_21_9_to_tile_21_10_1;
	wire horizontal_tile_21_9_to_tile_21_10_2;
	wire horizontal_tile_21_9_to_tile_21_10_3;
	wire horizontal_tile_21_10_to_tile_21_9_0;
	wire horizontal_tile_21_10_to_tile_21_9_1;
	wire horizontal_tile_21_10_to_tile_21_9_2;
	wire horizontal_tile_21_10_to_tile_21_9_3;

	wire horizontal_tile_22_9_to_tile_22_10_0;
	wire horizontal_tile_22_9_to_tile_22_10_1;
	wire horizontal_tile_22_9_to_tile_22_10_2;
	wire horizontal_tile_22_9_to_tile_22_10_3;
	wire horizontal_tile_22_10_to_tile_22_9_0;
	wire horizontal_tile_22_10_to_tile_22_9_1;
	wire horizontal_tile_22_10_to_tile_22_9_2;
	wire horizontal_tile_22_10_to_tile_22_9_3;

	wire horizontal_tile_23_9_to_tile_23_10_0;
	wire horizontal_tile_23_9_to_tile_23_10_1;
	wire horizontal_tile_23_9_to_tile_23_10_2;
	wire horizontal_tile_23_9_to_tile_23_10_3;
	wire horizontal_tile_23_10_to_tile_23_9_0;
	wire horizontal_tile_23_10_to_tile_23_9_1;
	wire horizontal_tile_23_10_to_tile_23_9_2;
	wire horizontal_tile_23_10_to_tile_23_9_3;

	wire horizontal_tile_24_9_to_tile_24_10_0;
	wire horizontal_tile_24_9_to_tile_24_10_1;
	wire horizontal_tile_24_9_to_tile_24_10_2;
	wire horizontal_tile_24_9_to_tile_24_10_3;
	wire horizontal_tile_24_10_to_tile_24_9_0;
	wire horizontal_tile_24_10_to_tile_24_9_1;
	wire horizontal_tile_24_10_to_tile_24_9_2;
	wire horizontal_tile_24_10_to_tile_24_9_3;

	wire horizontal_tile_25_9_to_tile_25_10_0;
	wire horizontal_tile_25_9_to_tile_25_10_1;
	wire horizontal_tile_25_9_to_tile_25_10_2;
	wire horizontal_tile_25_9_to_tile_25_10_3;
	wire horizontal_tile_25_10_to_tile_25_9_0;
	wire horizontal_tile_25_10_to_tile_25_9_1;
	wire horizontal_tile_25_10_to_tile_25_9_2;
	wire horizontal_tile_25_10_to_tile_25_9_3;

	wire horizontal_tile_26_9_to_tile_26_10_0;
	wire horizontal_tile_26_9_to_tile_26_10_1;
	wire horizontal_tile_26_9_to_tile_26_10_2;
	wire horizontal_tile_26_9_to_tile_26_10_3;
	wire horizontal_tile_26_10_to_tile_26_9_0;
	wire horizontal_tile_26_10_to_tile_26_9_1;
	wire horizontal_tile_26_10_to_tile_26_9_2;
	wire horizontal_tile_26_10_to_tile_26_9_3;

	wire horizontal_tile_27_9_to_tile_27_10_0;
	wire horizontal_tile_27_9_to_tile_27_10_1;
	wire horizontal_tile_27_9_to_tile_27_10_2;
	wire horizontal_tile_27_9_to_tile_27_10_3;
	wire horizontal_tile_27_10_to_tile_27_9_0;
	wire horizontal_tile_27_10_to_tile_27_9_1;
	wire horizontal_tile_27_10_to_tile_27_9_2;
	wire horizontal_tile_27_10_to_tile_27_9_3;

	wire horizontal_tile_28_9_to_tile_28_10_0;
	wire horizontal_tile_28_9_to_tile_28_10_1;
	wire horizontal_tile_28_9_to_tile_28_10_2;
	wire horizontal_tile_28_9_to_tile_28_10_3;
	wire horizontal_tile_28_10_to_tile_28_9_0;
	wire horizontal_tile_28_10_to_tile_28_9_1;
	wire horizontal_tile_28_10_to_tile_28_9_2;
	wire horizontal_tile_28_10_to_tile_28_9_3;

	wire horizontal_tile_29_9_to_tile_29_10_0;
	wire horizontal_tile_29_9_to_tile_29_10_1;
	wire horizontal_tile_29_9_to_tile_29_10_2;
	wire horizontal_tile_29_9_to_tile_29_10_3;
	wire horizontal_tile_29_10_to_tile_29_9_0;
	wire horizontal_tile_29_10_to_tile_29_9_1;
	wire horizontal_tile_29_10_to_tile_29_9_2;
	wire horizontal_tile_29_10_to_tile_29_9_3;

	wire horizontal_tile_30_9_to_tile_30_10_0;
	wire horizontal_tile_30_9_to_tile_30_10_1;
	wire horizontal_tile_30_9_to_tile_30_10_2;
	wire horizontal_tile_30_9_to_tile_30_10_3;
	wire horizontal_tile_30_10_to_tile_30_9_0;
	wire horizontal_tile_30_10_to_tile_30_9_1;
	wire horizontal_tile_30_10_to_tile_30_9_2;
	wire horizontal_tile_30_10_to_tile_30_9_3;

	wire horizontal_tile_31_9_to_tile_31_10_0;
	wire horizontal_tile_31_9_to_tile_31_10_1;
	wire horizontal_tile_31_9_to_tile_31_10_2;
	wire horizontal_tile_31_9_to_tile_31_10_3;
	wire horizontal_tile_31_10_to_tile_31_9_0;
	wire horizontal_tile_31_10_to_tile_31_9_1;
	wire horizontal_tile_31_10_to_tile_31_9_2;
	wire horizontal_tile_31_10_to_tile_31_9_3;

	wire horizontal_tile_0_10_to_tile_0_11_0;
	wire horizontal_tile_0_10_to_tile_0_11_1;
	wire horizontal_tile_0_10_to_tile_0_11_2;
	wire horizontal_tile_0_10_to_tile_0_11_3;
	wire horizontal_tile_0_11_to_tile_0_10_0;
	wire horizontal_tile_0_11_to_tile_0_10_1;
	wire horizontal_tile_0_11_to_tile_0_10_2;
	wire horizontal_tile_0_11_to_tile_0_10_3;

	wire horizontal_tile_1_10_to_tile_1_11_0;
	wire horizontal_tile_1_10_to_tile_1_11_1;
	wire horizontal_tile_1_10_to_tile_1_11_2;
	wire horizontal_tile_1_10_to_tile_1_11_3;
	wire horizontal_tile_1_11_to_tile_1_10_0;
	wire horizontal_tile_1_11_to_tile_1_10_1;
	wire horizontal_tile_1_11_to_tile_1_10_2;
	wire horizontal_tile_1_11_to_tile_1_10_3;

	wire horizontal_tile_2_10_to_tile_2_11_0;
	wire horizontal_tile_2_10_to_tile_2_11_1;
	wire horizontal_tile_2_10_to_tile_2_11_2;
	wire horizontal_tile_2_10_to_tile_2_11_3;
	wire horizontal_tile_2_11_to_tile_2_10_0;
	wire horizontal_tile_2_11_to_tile_2_10_1;
	wire horizontal_tile_2_11_to_tile_2_10_2;
	wire horizontal_tile_2_11_to_tile_2_10_3;

	wire horizontal_tile_3_10_to_tile_3_11_0;
	wire horizontal_tile_3_10_to_tile_3_11_1;
	wire horizontal_tile_3_10_to_tile_3_11_2;
	wire horizontal_tile_3_10_to_tile_3_11_3;
	wire horizontal_tile_3_11_to_tile_3_10_0;
	wire horizontal_tile_3_11_to_tile_3_10_1;
	wire horizontal_tile_3_11_to_tile_3_10_2;
	wire horizontal_tile_3_11_to_tile_3_10_3;

	wire horizontal_tile_4_10_to_tile_4_11_0;
	wire horizontal_tile_4_10_to_tile_4_11_1;
	wire horizontal_tile_4_10_to_tile_4_11_2;
	wire horizontal_tile_4_10_to_tile_4_11_3;
	wire horizontal_tile_4_11_to_tile_4_10_0;
	wire horizontal_tile_4_11_to_tile_4_10_1;
	wire horizontal_tile_4_11_to_tile_4_10_2;
	wire horizontal_tile_4_11_to_tile_4_10_3;

	wire horizontal_tile_5_10_to_tile_5_11_0;
	wire horizontal_tile_5_10_to_tile_5_11_1;
	wire horizontal_tile_5_10_to_tile_5_11_2;
	wire horizontal_tile_5_10_to_tile_5_11_3;
	wire horizontal_tile_5_11_to_tile_5_10_0;
	wire horizontal_tile_5_11_to_tile_5_10_1;
	wire horizontal_tile_5_11_to_tile_5_10_2;
	wire horizontal_tile_5_11_to_tile_5_10_3;

	wire horizontal_tile_6_10_to_tile_6_11_0;
	wire horizontal_tile_6_10_to_tile_6_11_1;
	wire horizontal_tile_6_10_to_tile_6_11_2;
	wire horizontal_tile_6_10_to_tile_6_11_3;
	wire horizontal_tile_6_11_to_tile_6_10_0;
	wire horizontal_tile_6_11_to_tile_6_10_1;
	wire horizontal_tile_6_11_to_tile_6_10_2;
	wire horizontal_tile_6_11_to_tile_6_10_3;

	wire horizontal_tile_7_10_to_tile_7_11_0;
	wire horizontal_tile_7_10_to_tile_7_11_1;
	wire horizontal_tile_7_10_to_tile_7_11_2;
	wire horizontal_tile_7_10_to_tile_7_11_3;
	wire horizontal_tile_7_11_to_tile_7_10_0;
	wire horizontal_tile_7_11_to_tile_7_10_1;
	wire horizontal_tile_7_11_to_tile_7_10_2;
	wire horizontal_tile_7_11_to_tile_7_10_3;

	wire horizontal_tile_8_10_to_tile_8_11_0;
	wire horizontal_tile_8_10_to_tile_8_11_1;
	wire horizontal_tile_8_10_to_tile_8_11_2;
	wire horizontal_tile_8_10_to_tile_8_11_3;
	wire horizontal_tile_8_11_to_tile_8_10_0;
	wire horizontal_tile_8_11_to_tile_8_10_1;
	wire horizontal_tile_8_11_to_tile_8_10_2;
	wire horizontal_tile_8_11_to_tile_8_10_3;

	wire horizontal_tile_9_10_to_tile_9_11_0;
	wire horizontal_tile_9_10_to_tile_9_11_1;
	wire horizontal_tile_9_10_to_tile_9_11_2;
	wire horizontal_tile_9_10_to_tile_9_11_3;
	wire horizontal_tile_9_11_to_tile_9_10_0;
	wire horizontal_tile_9_11_to_tile_9_10_1;
	wire horizontal_tile_9_11_to_tile_9_10_2;
	wire horizontal_tile_9_11_to_tile_9_10_3;

	wire horizontal_tile_10_10_to_tile_10_11_0;
	wire horizontal_tile_10_10_to_tile_10_11_1;
	wire horizontal_tile_10_10_to_tile_10_11_2;
	wire horizontal_tile_10_10_to_tile_10_11_3;
	wire horizontal_tile_10_11_to_tile_10_10_0;
	wire horizontal_tile_10_11_to_tile_10_10_1;
	wire horizontal_tile_10_11_to_tile_10_10_2;
	wire horizontal_tile_10_11_to_tile_10_10_3;

	wire horizontal_tile_11_10_to_tile_11_11_0;
	wire horizontal_tile_11_10_to_tile_11_11_1;
	wire horizontal_tile_11_10_to_tile_11_11_2;
	wire horizontal_tile_11_10_to_tile_11_11_3;
	wire horizontal_tile_11_11_to_tile_11_10_0;
	wire horizontal_tile_11_11_to_tile_11_10_1;
	wire horizontal_tile_11_11_to_tile_11_10_2;
	wire horizontal_tile_11_11_to_tile_11_10_3;

	wire horizontal_tile_12_10_to_tile_12_11_0;
	wire horizontal_tile_12_10_to_tile_12_11_1;
	wire horizontal_tile_12_10_to_tile_12_11_2;
	wire horizontal_tile_12_10_to_tile_12_11_3;
	wire horizontal_tile_12_11_to_tile_12_10_0;
	wire horizontal_tile_12_11_to_tile_12_10_1;
	wire horizontal_tile_12_11_to_tile_12_10_2;
	wire horizontal_tile_12_11_to_tile_12_10_3;

	wire horizontal_tile_13_10_to_tile_13_11_0;
	wire horizontal_tile_13_10_to_tile_13_11_1;
	wire horizontal_tile_13_10_to_tile_13_11_2;
	wire horizontal_tile_13_10_to_tile_13_11_3;
	wire horizontal_tile_13_11_to_tile_13_10_0;
	wire horizontal_tile_13_11_to_tile_13_10_1;
	wire horizontal_tile_13_11_to_tile_13_10_2;
	wire horizontal_tile_13_11_to_tile_13_10_3;

	wire horizontal_tile_14_10_to_tile_14_11_0;
	wire horizontal_tile_14_10_to_tile_14_11_1;
	wire horizontal_tile_14_10_to_tile_14_11_2;
	wire horizontal_tile_14_10_to_tile_14_11_3;
	wire horizontal_tile_14_11_to_tile_14_10_0;
	wire horizontal_tile_14_11_to_tile_14_10_1;
	wire horizontal_tile_14_11_to_tile_14_10_2;
	wire horizontal_tile_14_11_to_tile_14_10_3;

	wire horizontal_tile_15_10_to_tile_15_11_0;
	wire horizontal_tile_15_10_to_tile_15_11_1;
	wire horizontal_tile_15_10_to_tile_15_11_2;
	wire horizontal_tile_15_10_to_tile_15_11_3;
	wire horizontal_tile_15_11_to_tile_15_10_0;
	wire horizontal_tile_15_11_to_tile_15_10_1;
	wire horizontal_tile_15_11_to_tile_15_10_2;
	wire horizontal_tile_15_11_to_tile_15_10_3;

	wire horizontal_tile_16_10_to_tile_16_11_0;
	wire horizontal_tile_16_10_to_tile_16_11_1;
	wire horizontal_tile_16_10_to_tile_16_11_2;
	wire horizontal_tile_16_10_to_tile_16_11_3;
	wire horizontal_tile_16_11_to_tile_16_10_0;
	wire horizontal_tile_16_11_to_tile_16_10_1;
	wire horizontal_tile_16_11_to_tile_16_10_2;
	wire horizontal_tile_16_11_to_tile_16_10_3;

	wire horizontal_tile_17_10_to_tile_17_11_0;
	wire horizontal_tile_17_10_to_tile_17_11_1;
	wire horizontal_tile_17_10_to_tile_17_11_2;
	wire horizontal_tile_17_10_to_tile_17_11_3;
	wire horizontal_tile_17_11_to_tile_17_10_0;
	wire horizontal_tile_17_11_to_tile_17_10_1;
	wire horizontal_tile_17_11_to_tile_17_10_2;
	wire horizontal_tile_17_11_to_tile_17_10_3;

	wire horizontal_tile_18_10_to_tile_18_11_0;
	wire horizontal_tile_18_10_to_tile_18_11_1;
	wire horizontal_tile_18_10_to_tile_18_11_2;
	wire horizontal_tile_18_10_to_tile_18_11_3;
	wire horizontal_tile_18_11_to_tile_18_10_0;
	wire horizontal_tile_18_11_to_tile_18_10_1;
	wire horizontal_tile_18_11_to_tile_18_10_2;
	wire horizontal_tile_18_11_to_tile_18_10_3;

	wire horizontal_tile_19_10_to_tile_19_11_0;
	wire horizontal_tile_19_10_to_tile_19_11_1;
	wire horizontal_tile_19_10_to_tile_19_11_2;
	wire horizontal_tile_19_10_to_tile_19_11_3;
	wire horizontal_tile_19_11_to_tile_19_10_0;
	wire horizontal_tile_19_11_to_tile_19_10_1;
	wire horizontal_tile_19_11_to_tile_19_10_2;
	wire horizontal_tile_19_11_to_tile_19_10_3;

	wire horizontal_tile_20_10_to_tile_20_11_0;
	wire horizontal_tile_20_10_to_tile_20_11_1;
	wire horizontal_tile_20_10_to_tile_20_11_2;
	wire horizontal_tile_20_10_to_tile_20_11_3;
	wire horizontal_tile_20_11_to_tile_20_10_0;
	wire horizontal_tile_20_11_to_tile_20_10_1;
	wire horizontal_tile_20_11_to_tile_20_10_2;
	wire horizontal_tile_20_11_to_tile_20_10_3;

	wire horizontal_tile_21_10_to_tile_21_11_0;
	wire horizontal_tile_21_10_to_tile_21_11_1;
	wire horizontal_tile_21_10_to_tile_21_11_2;
	wire horizontal_tile_21_10_to_tile_21_11_3;
	wire horizontal_tile_21_11_to_tile_21_10_0;
	wire horizontal_tile_21_11_to_tile_21_10_1;
	wire horizontal_tile_21_11_to_tile_21_10_2;
	wire horizontal_tile_21_11_to_tile_21_10_3;

	wire horizontal_tile_22_10_to_tile_22_11_0;
	wire horizontal_tile_22_10_to_tile_22_11_1;
	wire horizontal_tile_22_10_to_tile_22_11_2;
	wire horizontal_tile_22_10_to_tile_22_11_3;
	wire horizontal_tile_22_11_to_tile_22_10_0;
	wire horizontal_tile_22_11_to_tile_22_10_1;
	wire horizontal_tile_22_11_to_tile_22_10_2;
	wire horizontal_tile_22_11_to_tile_22_10_3;

	wire horizontal_tile_23_10_to_tile_23_11_0;
	wire horizontal_tile_23_10_to_tile_23_11_1;
	wire horizontal_tile_23_10_to_tile_23_11_2;
	wire horizontal_tile_23_10_to_tile_23_11_3;
	wire horizontal_tile_23_11_to_tile_23_10_0;
	wire horizontal_tile_23_11_to_tile_23_10_1;
	wire horizontal_tile_23_11_to_tile_23_10_2;
	wire horizontal_tile_23_11_to_tile_23_10_3;

	wire horizontal_tile_24_10_to_tile_24_11_0;
	wire horizontal_tile_24_10_to_tile_24_11_1;
	wire horizontal_tile_24_10_to_tile_24_11_2;
	wire horizontal_tile_24_10_to_tile_24_11_3;
	wire horizontal_tile_24_11_to_tile_24_10_0;
	wire horizontal_tile_24_11_to_tile_24_10_1;
	wire horizontal_tile_24_11_to_tile_24_10_2;
	wire horizontal_tile_24_11_to_tile_24_10_3;

	wire horizontal_tile_25_10_to_tile_25_11_0;
	wire horizontal_tile_25_10_to_tile_25_11_1;
	wire horizontal_tile_25_10_to_tile_25_11_2;
	wire horizontal_tile_25_10_to_tile_25_11_3;
	wire horizontal_tile_25_11_to_tile_25_10_0;
	wire horizontal_tile_25_11_to_tile_25_10_1;
	wire horizontal_tile_25_11_to_tile_25_10_2;
	wire horizontal_tile_25_11_to_tile_25_10_3;

	wire horizontal_tile_26_10_to_tile_26_11_0;
	wire horizontal_tile_26_10_to_tile_26_11_1;
	wire horizontal_tile_26_10_to_tile_26_11_2;
	wire horizontal_tile_26_10_to_tile_26_11_3;
	wire horizontal_tile_26_11_to_tile_26_10_0;
	wire horizontal_tile_26_11_to_tile_26_10_1;
	wire horizontal_tile_26_11_to_tile_26_10_2;
	wire horizontal_tile_26_11_to_tile_26_10_3;

	wire horizontal_tile_27_10_to_tile_27_11_0;
	wire horizontal_tile_27_10_to_tile_27_11_1;
	wire horizontal_tile_27_10_to_tile_27_11_2;
	wire horizontal_tile_27_10_to_tile_27_11_3;
	wire horizontal_tile_27_11_to_tile_27_10_0;
	wire horizontal_tile_27_11_to_tile_27_10_1;
	wire horizontal_tile_27_11_to_tile_27_10_2;
	wire horizontal_tile_27_11_to_tile_27_10_3;

	wire horizontal_tile_28_10_to_tile_28_11_0;
	wire horizontal_tile_28_10_to_tile_28_11_1;
	wire horizontal_tile_28_10_to_tile_28_11_2;
	wire horizontal_tile_28_10_to_tile_28_11_3;
	wire horizontal_tile_28_11_to_tile_28_10_0;
	wire horizontal_tile_28_11_to_tile_28_10_1;
	wire horizontal_tile_28_11_to_tile_28_10_2;
	wire horizontal_tile_28_11_to_tile_28_10_3;

	wire horizontal_tile_29_10_to_tile_29_11_0;
	wire horizontal_tile_29_10_to_tile_29_11_1;
	wire horizontal_tile_29_10_to_tile_29_11_2;
	wire horizontal_tile_29_10_to_tile_29_11_3;
	wire horizontal_tile_29_11_to_tile_29_10_0;
	wire horizontal_tile_29_11_to_tile_29_10_1;
	wire horizontal_tile_29_11_to_tile_29_10_2;
	wire horizontal_tile_29_11_to_tile_29_10_3;

	wire horizontal_tile_30_10_to_tile_30_11_0;
	wire horizontal_tile_30_10_to_tile_30_11_1;
	wire horizontal_tile_30_10_to_tile_30_11_2;
	wire horizontal_tile_30_10_to_tile_30_11_3;
	wire horizontal_tile_30_11_to_tile_30_10_0;
	wire horizontal_tile_30_11_to_tile_30_10_1;
	wire horizontal_tile_30_11_to_tile_30_10_2;
	wire horizontal_tile_30_11_to_tile_30_10_3;

	wire horizontal_tile_31_10_to_tile_31_11_0;
	wire horizontal_tile_31_10_to_tile_31_11_1;
	wire horizontal_tile_31_10_to_tile_31_11_2;
	wire horizontal_tile_31_10_to_tile_31_11_3;
	wire horizontal_tile_31_11_to_tile_31_10_0;
	wire horizontal_tile_31_11_to_tile_31_10_1;
	wire horizontal_tile_31_11_to_tile_31_10_2;
	wire horizontal_tile_31_11_to_tile_31_10_3;

	wire horizontal_tile_0_11_to_tile_0_12_0;
	wire horizontal_tile_0_11_to_tile_0_12_1;
	wire horizontal_tile_0_11_to_tile_0_12_2;
	wire horizontal_tile_0_11_to_tile_0_12_3;
	wire horizontal_tile_0_12_to_tile_0_11_0;
	wire horizontal_tile_0_12_to_tile_0_11_1;
	wire horizontal_tile_0_12_to_tile_0_11_2;
	wire horizontal_tile_0_12_to_tile_0_11_3;

	wire horizontal_tile_1_11_to_tile_1_12_0;
	wire horizontal_tile_1_11_to_tile_1_12_1;
	wire horizontal_tile_1_11_to_tile_1_12_2;
	wire horizontal_tile_1_11_to_tile_1_12_3;
	wire horizontal_tile_1_12_to_tile_1_11_0;
	wire horizontal_tile_1_12_to_tile_1_11_1;
	wire horizontal_tile_1_12_to_tile_1_11_2;
	wire horizontal_tile_1_12_to_tile_1_11_3;

	wire horizontal_tile_2_11_to_tile_2_12_0;
	wire horizontal_tile_2_11_to_tile_2_12_1;
	wire horizontal_tile_2_11_to_tile_2_12_2;
	wire horizontal_tile_2_11_to_tile_2_12_3;
	wire horizontal_tile_2_12_to_tile_2_11_0;
	wire horizontal_tile_2_12_to_tile_2_11_1;
	wire horizontal_tile_2_12_to_tile_2_11_2;
	wire horizontal_tile_2_12_to_tile_2_11_3;

	wire horizontal_tile_3_11_to_tile_3_12_0;
	wire horizontal_tile_3_11_to_tile_3_12_1;
	wire horizontal_tile_3_11_to_tile_3_12_2;
	wire horizontal_tile_3_11_to_tile_3_12_3;
	wire horizontal_tile_3_12_to_tile_3_11_0;
	wire horizontal_tile_3_12_to_tile_3_11_1;
	wire horizontal_tile_3_12_to_tile_3_11_2;
	wire horizontal_tile_3_12_to_tile_3_11_3;

	wire horizontal_tile_4_11_to_tile_4_12_0;
	wire horizontal_tile_4_11_to_tile_4_12_1;
	wire horizontal_tile_4_11_to_tile_4_12_2;
	wire horizontal_tile_4_11_to_tile_4_12_3;
	wire horizontal_tile_4_12_to_tile_4_11_0;
	wire horizontal_tile_4_12_to_tile_4_11_1;
	wire horizontal_tile_4_12_to_tile_4_11_2;
	wire horizontal_tile_4_12_to_tile_4_11_3;

	wire horizontal_tile_5_11_to_tile_5_12_0;
	wire horizontal_tile_5_11_to_tile_5_12_1;
	wire horizontal_tile_5_11_to_tile_5_12_2;
	wire horizontal_tile_5_11_to_tile_5_12_3;
	wire horizontal_tile_5_12_to_tile_5_11_0;
	wire horizontal_tile_5_12_to_tile_5_11_1;
	wire horizontal_tile_5_12_to_tile_5_11_2;
	wire horizontal_tile_5_12_to_tile_5_11_3;

	wire horizontal_tile_6_11_to_tile_6_12_0;
	wire horizontal_tile_6_11_to_tile_6_12_1;
	wire horizontal_tile_6_11_to_tile_6_12_2;
	wire horizontal_tile_6_11_to_tile_6_12_3;
	wire horizontal_tile_6_12_to_tile_6_11_0;
	wire horizontal_tile_6_12_to_tile_6_11_1;
	wire horizontal_tile_6_12_to_tile_6_11_2;
	wire horizontal_tile_6_12_to_tile_6_11_3;

	wire horizontal_tile_7_11_to_tile_7_12_0;
	wire horizontal_tile_7_11_to_tile_7_12_1;
	wire horizontal_tile_7_11_to_tile_7_12_2;
	wire horizontal_tile_7_11_to_tile_7_12_3;
	wire horizontal_tile_7_12_to_tile_7_11_0;
	wire horizontal_tile_7_12_to_tile_7_11_1;
	wire horizontal_tile_7_12_to_tile_7_11_2;
	wire horizontal_tile_7_12_to_tile_7_11_3;

	wire horizontal_tile_8_11_to_tile_8_12_0;
	wire horizontal_tile_8_11_to_tile_8_12_1;
	wire horizontal_tile_8_11_to_tile_8_12_2;
	wire horizontal_tile_8_11_to_tile_8_12_3;
	wire horizontal_tile_8_12_to_tile_8_11_0;
	wire horizontal_tile_8_12_to_tile_8_11_1;
	wire horizontal_tile_8_12_to_tile_8_11_2;
	wire horizontal_tile_8_12_to_tile_8_11_3;

	wire horizontal_tile_9_11_to_tile_9_12_0;
	wire horizontal_tile_9_11_to_tile_9_12_1;
	wire horizontal_tile_9_11_to_tile_9_12_2;
	wire horizontal_tile_9_11_to_tile_9_12_3;
	wire horizontal_tile_9_12_to_tile_9_11_0;
	wire horizontal_tile_9_12_to_tile_9_11_1;
	wire horizontal_tile_9_12_to_tile_9_11_2;
	wire horizontal_tile_9_12_to_tile_9_11_3;

	wire horizontal_tile_10_11_to_tile_10_12_0;
	wire horizontal_tile_10_11_to_tile_10_12_1;
	wire horizontal_tile_10_11_to_tile_10_12_2;
	wire horizontal_tile_10_11_to_tile_10_12_3;
	wire horizontal_tile_10_12_to_tile_10_11_0;
	wire horizontal_tile_10_12_to_tile_10_11_1;
	wire horizontal_tile_10_12_to_tile_10_11_2;
	wire horizontal_tile_10_12_to_tile_10_11_3;

	wire horizontal_tile_11_11_to_tile_11_12_0;
	wire horizontal_tile_11_11_to_tile_11_12_1;
	wire horizontal_tile_11_11_to_tile_11_12_2;
	wire horizontal_tile_11_11_to_tile_11_12_3;
	wire horizontal_tile_11_12_to_tile_11_11_0;
	wire horizontal_tile_11_12_to_tile_11_11_1;
	wire horizontal_tile_11_12_to_tile_11_11_2;
	wire horizontal_tile_11_12_to_tile_11_11_3;

	wire horizontal_tile_12_11_to_tile_12_12_0;
	wire horizontal_tile_12_11_to_tile_12_12_1;
	wire horizontal_tile_12_11_to_tile_12_12_2;
	wire horizontal_tile_12_11_to_tile_12_12_3;
	wire horizontal_tile_12_12_to_tile_12_11_0;
	wire horizontal_tile_12_12_to_tile_12_11_1;
	wire horizontal_tile_12_12_to_tile_12_11_2;
	wire horizontal_tile_12_12_to_tile_12_11_3;

	wire horizontal_tile_13_11_to_tile_13_12_0;
	wire horizontal_tile_13_11_to_tile_13_12_1;
	wire horizontal_tile_13_11_to_tile_13_12_2;
	wire horizontal_tile_13_11_to_tile_13_12_3;
	wire horizontal_tile_13_12_to_tile_13_11_0;
	wire horizontal_tile_13_12_to_tile_13_11_1;
	wire horizontal_tile_13_12_to_tile_13_11_2;
	wire horizontal_tile_13_12_to_tile_13_11_3;

	wire horizontal_tile_14_11_to_tile_14_12_0;
	wire horizontal_tile_14_11_to_tile_14_12_1;
	wire horizontal_tile_14_11_to_tile_14_12_2;
	wire horizontal_tile_14_11_to_tile_14_12_3;
	wire horizontal_tile_14_12_to_tile_14_11_0;
	wire horizontal_tile_14_12_to_tile_14_11_1;
	wire horizontal_tile_14_12_to_tile_14_11_2;
	wire horizontal_tile_14_12_to_tile_14_11_3;

	wire horizontal_tile_15_11_to_tile_15_12_0;
	wire horizontal_tile_15_11_to_tile_15_12_1;
	wire horizontal_tile_15_11_to_tile_15_12_2;
	wire horizontal_tile_15_11_to_tile_15_12_3;
	wire horizontal_tile_15_12_to_tile_15_11_0;
	wire horizontal_tile_15_12_to_tile_15_11_1;
	wire horizontal_tile_15_12_to_tile_15_11_2;
	wire horizontal_tile_15_12_to_tile_15_11_3;

	wire horizontal_tile_16_11_to_tile_16_12_0;
	wire horizontal_tile_16_11_to_tile_16_12_1;
	wire horizontal_tile_16_11_to_tile_16_12_2;
	wire horizontal_tile_16_11_to_tile_16_12_3;
	wire horizontal_tile_16_12_to_tile_16_11_0;
	wire horizontal_tile_16_12_to_tile_16_11_1;
	wire horizontal_tile_16_12_to_tile_16_11_2;
	wire horizontal_tile_16_12_to_tile_16_11_3;

	wire horizontal_tile_17_11_to_tile_17_12_0;
	wire horizontal_tile_17_11_to_tile_17_12_1;
	wire horizontal_tile_17_11_to_tile_17_12_2;
	wire horizontal_tile_17_11_to_tile_17_12_3;
	wire horizontal_tile_17_12_to_tile_17_11_0;
	wire horizontal_tile_17_12_to_tile_17_11_1;
	wire horizontal_tile_17_12_to_tile_17_11_2;
	wire horizontal_tile_17_12_to_tile_17_11_3;

	wire horizontal_tile_18_11_to_tile_18_12_0;
	wire horizontal_tile_18_11_to_tile_18_12_1;
	wire horizontal_tile_18_11_to_tile_18_12_2;
	wire horizontal_tile_18_11_to_tile_18_12_3;
	wire horizontal_tile_18_12_to_tile_18_11_0;
	wire horizontal_tile_18_12_to_tile_18_11_1;
	wire horizontal_tile_18_12_to_tile_18_11_2;
	wire horizontal_tile_18_12_to_tile_18_11_3;

	wire horizontal_tile_19_11_to_tile_19_12_0;
	wire horizontal_tile_19_11_to_tile_19_12_1;
	wire horizontal_tile_19_11_to_tile_19_12_2;
	wire horizontal_tile_19_11_to_tile_19_12_3;
	wire horizontal_tile_19_12_to_tile_19_11_0;
	wire horizontal_tile_19_12_to_tile_19_11_1;
	wire horizontal_tile_19_12_to_tile_19_11_2;
	wire horizontal_tile_19_12_to_tile_19_11_3;

	wire horizontal_tile_20_11_to_tile_20_12_0;
	wire horizontal_tile_20_11_to_tile_20_12_1;
	wire horizontal_tile_20_11_to_tile_20_12_2;
	wire horizontal_tile_20_11_to_tile_20_12_3;
	wire horizontal_tile_20_12_to_tile_20_11_0;
	wire horizontal_tile_20_12_to_tile_20_11_1;
	wire horizontal_tile_20_12_to_tile_20_11_2;
	wire horizontal_tile_20_12_to_tile_20_11_3;

	wire horizontal_tile_21_11_to_tile_21_12_0;
	wire horizontal_tile_21_11_to_tile_21_12_1;
	wire horizontal_tile_21_11_to_tile_21_12_2;
	wire horizontal_tile_21_11_to_tile_21_12_3;
	wire horizontal_tile_21_12_to_tile_21_11_0;
	wire horizontal_tile_21_12_to_tile_21_11_1;
	wire horizontal_tile_21_12_to_tile_21_11_2;
	wire horizontal_tile_21_12_to_tile_21_11_3;

	wire horizontal_tile_22_11_to_tile_22_12_0;
	wire horizontal_tile_22_11_to_tile_22_12_1;
	wire horizontal_tile_22_11_to_tile_22_12_2;
	wire horizontal_tile_22_11_to_tile_22_12_3;
	wire horizontal_tile_22_12_to_tile_22_11_0;
	wire horizontal_tile_22_12_to_tile_22_11_1;
	wire horizontal_tile_22_12_to_tile_22_11_2;
	wire horizontal_tile_22_12_to_tile_22_11_3;

	wire horizontal_tile_23_11_to_tile_23_12_0;
	wire horizontal_tile_23_11_to_tile_23_12_1;
	wire horizontal_tile_23_11_to_tile_23_12_2;
	wire horizontal_tile_23_11_to_tile_23_12_3;
	wire horizontal_tile_23_12_to_tile_23_11_0;
	wire horizontal_tile_23_12_to_tile_23_11_1;
	wire horizontal_tile_23_12_to_tile_23_11_2;
	wire horizontal_tile_23_12_to_tile_23_11_3;

	wire horizontal_tile_24_11_to_tile_24_12_0;
	wire horizontal_tile_24_11_to_tile_24_12_1;
	wire horizontal_tile_24_11_to_tile_24_12_2;
	wire horizontal_tile_24_11_to_tile_24_12_3;
	wire horizontal_tile_24_12_to_tile_24_11_0;
	wire horizontal_tile_24_12_to_tile_24_11_1;
	wire horizontal_tile_24_12_to_tile_24_11_2;
	wire horizontal_tile_24_12_to_tile_24_11_3;

	wire horizontal_tile_25_11_to_tile_25_12_0;
	wire horizontal_tile_25_11_to_tile_25_12_1;
	wire horizontal_tile_25_11_to_tile_25_12_2;
	wire horizontal_tile_25_11_to_tile_25_12_3;
	wire horizontal_tile_25_12_to_tile_25_11_0;
	wire horizontal_tile_25_12_to_tile_25_11_1;
	wire horizontal_tile_25_12_to_tile_25_11_2;
	wire horizontal_tile_25_12_to_tile_25_11_3;

	wire horizontal_tile_26_11_to_tile_26_12_0;
	wire horizontal_tile_26_11_to_tile_26_12_1;
	wire horizontal_tile_26_11_to_tile_26_12_2;
	wire horizontal_tile_26_11_to_tile_26_12_3;
	wire horizontal_tile_26_12_to_tile_26_11_0;
	wire horizontal_tile_26_12_to_tile_26_11_1;
	wire horizontal_tile_26_12_to_tile_26_11_2;
	wire horizontal_tile_26_12_to_tile_26_11_3;

	wire horizontal_tile_27_11_to_tile_27_12_0;
	wire horizontal_tile_27_11_to_tile_27_12_1;
	wire horizontal_tile_27_11_to_tile_27_12_2;
	wire horizontal_tile_27_11_to_tile_27_12_3;
	wire horizontal_tile_27_12_to_tile_27_11_0;
	wire horizontal_tile_27_12_to_tile_27_11_1;
	wire horizontal_tile_27_12_to_tile_27_11_2;
	wire horizontal_tile_27_12_to_tile_27_11_3;

	wire horizontal_tile_28_11_to_tile_28_12_0;
	wire horizontal_tile_28_11_to_tile_28_12_1;
	wire horizontal_tile_28_11_to_tile_28_12_2;
	wire horizontal_tile_28_11_to_tile_28_12_3;
	wire horizontal_tile_28_12_to_tile_28_11_0;
	wire horizontal_tile_28_12_to_tile_28_11_1;
	wire horizontal_tile_28_12_to_tile_28_11_2;
	wire horizontal_tile_28_12_to_tile_28_11_3;

	wire horizontal_tile_29_11_to_tile_29_12_0;
	wire horizontal_tile_29_11_to_tile_29_12_1;
	wire horizontal_tile_29_11_to_tile_29_12_2;
	wire horizontal_tile_29_11_to_tile_29_12_3;
	wire horizontal_tile_29_12_to_tile_29_11_0;
	wire horizontal_tile_29_12_to_tile_29_11_1;
	wire horizontal_tile_29_12_to_tile_29_11_2;
	wire horizontal_tile_29_12_to_tile_29_11_3;

	wire horizontal_tile_30_11_to_tile_30_12_0;
	wire horizontal_tile_30_11_to_tile_30_12_1;
	wire horizontal_tile_30_11_to_tile_30_12_2;
	wire horizontal_tile_30_11_to_tile_30_12_3;
	wire horizontal_tile_30_12_to_tile_30_11_0;
	wire horizontal_tile_30_12_to_tile_30_11_1;
	wire horizontal_tile_30_12_to_tile_30_11_2;
	wire horizontal_tile_30_12_to_tile_30_11_3;

	wire horizontal_tile_31_11_to_tile_31_12_0;
	wire horizontal_tile_31_11_to_tile_31_12_1;
	wire horizontal_tile_31_11_to_tile_31_12_2;
	wire horizontal_tile_31_11_to_tile_31_12_3;
	wire horizontal_tile_31_12_to_tile_31_11_0;
	wire horizontal_tile_31_12_to_tile_31_11_1;
	wire horizontal_tile_31_12_to_tile_31_11_2;
	wire horizontal_tile_31_12_to_tile_31_11_3;

	wire horizontal_tile_0_12_to_tile_0_13_0;
	wire horizontal_tile_0_12_to_tile_0_13_1;
	wire horizontal_tile_0_12_to_tile_0_13_2;
	wire horizontal_tile_0_12_to_tile_0_13_3;
	wire horizontal_tile_0_13_to_tile_0_12_0;
	wire horizontal_tile_0_13_to_tile_0_12_1;
	wire horizontal_tile_0_13_to_tile_0_12_2;
	wire horizontal_tile_0_13_to_tile_0_12_3;

	wire horizontal_tile_1_12_to_tile_1_13_0;
	wire horizontal_tile_1_12_to_tile_1_13_1;
	wire horizontal_tile_1_12_to_tile_1_13_2;
	wire horizontal_tile_1_12_to_tile_1_13_3;
	wire horizontal_tile_1_13_to_tile_1_12_0;
	wire horizontal_tile_1_13_to_tile_1_12_1;
	wire horizontal_tile_1_13_to_tile_1_12_2;
	wire horizontal_tile_1_13_to_tile_1_12_3;

	wire horizontal_tile_2_12_to_tile_2_13_0;
	wire horizontal_tile_2_12_to_tile_2_13_1;
	wire horizontal_tile_2_12_to_tile_2_13_2;
	wire horizontal_tile_2_12_to_tile_2_13_3;
	wire horizontal_tile_2_13_to_tile_2_12_0;
	wire horizontal_tile_2_13_to_tile_2_12_1;
	wire horizontal_tile_2_13_to_tile_2_12_2;
	wire horizontal_tile_2_13_to_tile_2_12_3;

	wire horizontal_tile_3_12_to_tile_3_13_0;
	wire horizontal_tile_3_12_to_tile_3_13_1;
	wire horizontal_tile_3_12_to_tile_3_13_2;
	wire horizontal_tile_3_12_to_tile_3_13_3;
	wire horizontal_tile_3_13_to_tile_3_12_0;
	wire horizontal_tile_3_13_to_tile_3_12_1;
	wire horizontal_tile_3_13_to_tile_3_12_2;
	wire horizontal_tile_3_13_to_tile_3_12_3;

	wire horizontal_tile_4_12_to_tile_4_13_0;
	wire horizontal_tile_4_12_to_tile_4_13_1;
	wire horizontal_tile_4_12_to_tile_4_13_2;
	wire horizontal_tile_4_12_to_tile_4_13_3;
	wire horizontal_tile_4_13_to_tile_4_12_0;
	wire horizontal_tile_4_13_to_tile_4_12_1;
	wire horizontal_tile_4_13_to_tile_4_12_2;
	wire horizontal_tile_4_13_to_tile_4_12_3;

	wire horizontal_tile_5_12_to_tile_5_13_0;
	wire horizontal_tile_5_12_to_tile_5_13_1;
	wire horizontal_tile_5_12_to_tile_5_13_2;
	wire horizontal_tile_5_12_to_tile_5_13_3;
	wire horizontal_tile_5_13_to_tile_5_12_0;
	wire horizontal_tile_5_13_to_tile_5_12_1;
	wire horizontal_tile_5_13_to_tile_5_12_2;
	wire horizontal_tile_5_13_to_tile_5_12_3;

	wire horizontal_tile_6_12_to_tile_6_13_0;
	wire horizontal_tile_6_12_to_tile_6_13_1;
	wire horizontal_tile_6_12_to_tile_6_13_2;
	wire horizontal_tile_6_12_to_tile_6_13_3;
	wire horizontal_tile_6_13_to_tile_6_12_0;
	wire horizontal_tile_6_13_to_tile_6_12_1;
	wire horizontal_tile_6_13_to_tile_6_12_2;
	wire horizontal_tile_6_13_to_tile_6_12_3;

	wire horizontal_tile_7_12_to_tile_7_13_0;
	wire horizontal_tile_7_12_to_tile_7_13_1;
	wire horizontal_tile_7_12_to_tile_7_13_2;
	wire horizontal_tile_7_12_to_tile_7_13_3;
	wire horizontal_tile_7_13_to_tile_7_12_0;
	wire horizontal_tile_7_13_to_tile_7_12_1;
	wire horizontal_tile_7_13_to_tile_7_12_2;
	wire horizontal_tile_7_13_to_tile_7_12_3;

	wire horizontal_tile_8_12_to_tile_8_13_0;
	wire horizontal_tile_8_12_to_tile_8_13_1;
	wire horizontal_tile_8_12_to_tile_8_13_2;
	wire horizontal_tile_8_12_to_tile_8_13_3;
	wire horizontal_tile_8_13_to_tile_8_12_0;
	wire horizontal_tile_8_13_to_tile_8_12_1;
	wire horizontal_tile_8_13_to_tile_8_12_2;
	wire horizontal_tile_8_13_to_tile_8_12_3;

	wire horizontal_tile_9_12_to_tile_9_13_0;
	wire horizontal_tile_9_12_to_tile_9_13_1;
	wire horizontal_tile_9_12_to_tile_9_13_2;
	wire horizontal_tile_9_12_to_tile_9_13_3;
	wire horizontal_tile_9_13_to_tile_9_12_0;
	wire horizontal_tile_9_13_to_tile_9_12_1;
	wire horizontal_tile_9_13_to_tile_9_12_2;
	wire horizontal_tile_9_13_to_tile_9_12_3;

	wire horizontal_tile_10_12_to_tile_10_13_0;
	wire horizontal_tile_10_12_to_tile_10_13_1;
	wire horizontal_tile_10_12_to_tile_10_13_2;
	wire horizontal_tile_10_12_to_tile_10_13_3;
	wire horizontal_tile_10_13_to_tile_10_12_0;
	wire horizontal_tile_10_13_to_tile_10_12_1;
	wire horizontal_tile_10_13_to_tile_10_12_2;
	wire horizontal_tile_10_13_to_tile_10_12_3;

	wire horizontal_tile_11_12_to_tile_11_13_0;
	wire horizontal_tile_11_12_to_tile_11_13_1;
	wire horizontal_tile_11_12_to_tile_11_13_2;
	wire horizontal_tile_11_12_to_tile_11_13_3;
	wire horizontal_tile_11_13_to_tile_11_12_0;
	wire horizontal_tile_11_13_to_tile_11_12_1;
	wire horizontal_tile_11_13_to_tile_11_12_2;
	wire horizontal_tile_11_13_to_tile_11_12_3;

	wire horizontal_tile_12_12_to_tile_12_13_0;
	wire horizontal_tile_12_12_to_tile_12_13_1;
	wire horizontal_tile_12_12_to_tile_12_13_2;
	wire horizontal_tile_12_12_to_tile_12_13_3;
	wire horizontal_tile_12_13_to_tile_12_12_0;
	wire horizontal_tile_12_13_to_tile_12_12_1;
	wire horizontal_tile_12_13_to_tile_12_12_2;
	wire horizontal_tile_12_13_to_tile_12_12_3;

	wire horizontal_tile_13_12_to_tile_13_13_0;
	wire horizontal_tile_13_12_to_tile_13_13_1;
	wire horizontal_tile_13_12_to_tile_13_13_2;
	wire horizontal_tile_13_12_to_tile_13_13_3;
	wire horizontal_tile_13_13_to_tile_13_12_0;
	wire horizontal_tile_13_13_to_tile_13_12_1;
	wire horizontal_tile_13_13_to_tile_13_12_2;
	wire horizontal_tile_13_13_to_tile_13_12_3;

	wire horizontal_tile_14_12_to_tile_14_13_0;
	wire horizontal_tile_14_12_to_tile_14_13_1;
	wire horizontal_tile_14_12_to_tile_14_13_2;
	wire horizontal_tile_14_12_to_tile_14_13_3;
	wire horizontal_tile_14_13_to_tile_14_12_0;
	wire horizontal_tile_14_13_to_tile_14_12_1;
	wire horizontal_tile_14_13_to_tile_14_12_2;
	wire horizontal_tile_14_13_to_tile_14_12_3;

	wire horizontal_tile_15_12_to_tile_15_13_0;
	wire horizontal_tile_15_12_to_tile_15_13_1;
	wire horizontal_tile_15_12_to_tile_15_13_2;
	wire horizontal_tile_15_12_to_tile_15_13_3;
	wire horizontal_tile_15_13_to_tile_15_12_0;
	wire horizontal_tile_15_13_to_tile_15_12_1;
	wire horizontal_tile_15_13_to_tile_15_12_2;
	wire horizontal_tile_15_13_to_tile_15_12_3;

	wire horizontal_tile_16_12_to_tile_16_13_0;
	wire horizontal_tile_16_12_to_tile_16_13_1;
	wire horizontal_tile_16_12_to_tile_16_13_2;
	wire horizontal_tile_16_12_to_tile_16_13_3;
	wire horizontal_tile_16_13_to_tile_16_12_0;
	wire horizontal_tile_16_13_to_tile_16_12_1;
	wire horizontal_tile_16_13_to_tile_16_12_2;
	wire horizontal_tile_16_13_to_tile_16_12_3;

	wire horizontal_tile_17_12_to_tile_17_13_0;
	wire horizontal_tile_17_12_to_tile_17_13_1;
	wire horizontal_tile_17_12_to_tile_17_13_2;
	wire horizontal_tile_17_12_to_tile_17_13_3;
	wire horizontal_tile_17_13_to_tile_17_12_0;
	wire horizontal_tile_17_13_to_tile_17_12_1;
	wire horizontal_tile_17_13_to_tile_17_12_2;
	wire horizontal_tile_17_13_to_tile_17_12_3;

	wire horizontal_tile_18_12_to_tile_18_13_0;
	wire horizontal_tile_18_12_to_tile_18_13_1;
	wire horizontal_tile_18_12_to_tile_18_13_2;
	wire horizontal_tile_18_12_to_tile_18_13_3;
	wire horizontal_tile_18_13_to_tile_18_12_0;
	wire horizontal_tile_18_13_to_tile_18_12_1;
	wire horizontal_tile_18_13_to_tile_18_12_2;
	wire horizontal_tile_18_13_to_tile_18_12_3;

	wire horizontal_tile_19_12_to_tile_19_13_0;
	wire horizontal_tile_19_12_to_tile_19_13_1;
	wire horizontal_tile_19_12_to_tile_19_13_2;
	wire horizontal_tile_19_12_to_tile_19_13_3;
	wire horizontal_tile_19_13_to_tile_19_12_0;
	wire horizontal_tile_19_13_to_tile_19_12_1;
	wire horizontal_tile_19_13_to_tile_19_12_2;
	wire horizontal_tile_19_13_to_tile_19_12_3;

	wire horizontal_tile_20_12_to_tile_20_13_0;
	wire horizontal_tile_20_12_to_tile_20_13_1;
	wire horizontal_tile_20_12_to_tile_20_13_2;
	wire horizontal_tile_20_12_to_tile_20_13_3;
	wire horizontal_tile_20_13_to_tile_20_12_0;
	wire horizontal_tile_20_13_to_tile_20_12_1;
	wire horizontal_tile_20_13_to_tile_20_12_2;
	wire horizontal_tile_20_13_to_tile_20_12_3;

	wire horizontal_tile_21_12_to_tile_21_13_0;
	wire horizontal_tile_21_12_to_tile_21_13_1;
	wire horizontal_tile_21_12_to_tile_21_13_2;
	wire horizontal_tile_21_12_to_tile_21_13_3;
	wire horizontal_tile_21_13_to_tile_21_12_0;
	wire horizontal_tile_21_13_to_tile_21_12_1;
	wire horizontal_tile_21_13_to_tile_21_12_2;
	wire horizontal_tile_21_13_to_tile_21_12_3;

	wire horizontal_tile_22_12_to_tile_22_13_0;
	wire horizontal_tile_22_12_to_tile_22_13_1;
	wire horizontal_tile_22_12_to_tile_22_13_2;
	wire horizontal_tile_22_12_to_tile_22_13_3;
	wire horizontal_tile_22_13_to_tile_22_12_0;
	wire horizontal_tile_22_13_to_tile_22_12_1;
	wire horizontal_tile_22_13_to_tile_22_12_2;
	wire horizontal_tile_22_13_to_tile_22_12_3;

	wire horizontal_tile_23_12_to_tile_23_13_0;
	wire horizontal_tile_23_12_to_tile_23_13_1;
	wire horizontal_tile_23_12_to_tile_23_13_2;
	wire horizontal_tile_23_12_to_tile_23_13_3;
	wire horizontal_tile_23_13_to_tile_23_12_0;
	wire horizontal_tile_23_13_to_tile_23_12_1;
	wire horizontal_tile_23_13_to_tile_23_12_2;
	wire horizontal_tile_23_13_to_tile_23_12_3;

	wire horizontal_tile_24_12_to_tile_24_13_0;
	wire horizontal_tile_24_12_to_tile_24_13_1;
	wire horizontal_tile_24_12_to_tile_24_13_2;
	wire horizontal_tile_24_12_to_tile_24_13_3;
	wire horizontal_tile_24_13_to_tile_24_12_0;
	wire horizontal_tile_24_13_to_tile_24_12_1;
	wire horizontal_tile_24_13_to_tile_24_12_2;
	wire horizontal_tile_24_13_to_tile_24_12_3;

	wire horizontal_tile_25_12_to_tile_25_13_0;
	wire horizontal_tile_25_12_to_tile_25_13_1;
	wire horizontal_tile_25_12_to_tile_25_13_2;
	wire horizontal_tile_25_12_to_tile_25_13_3;
	wire horizontal_tile_25_13_to_tile_25_12_0;
	wire horizontal_tile_25_13_to_tile_25_12_1;
	wire horizontal_tile_25_13_to_tile_25_12_2;
	wire horizontal_tile_25_13_to_tile_25_12_3;

	wire horizontal_tile_26_12_to_tile_26_13_0;
	wire horizontal_tile_26_12_to_tile_26_13_1;
	wire horizontal_tile_26_12_to_tile_26_13_2;
	wire horizontal_tile_26_12_to_tile_26_13_3;
	wire horizontal_tile_26_13_to_tile_26_12_0;
	wire horizontal_tile_26_13_to_tile_26_12_1;
	wire horizontal_tile_26_13_to_tile_26_12_2;
	wire horizontal_tile_26_13_to_tile_26_12_3;

	wire horizontal_tile_27_12_to_tile_27_13_0;
	wire horizontal_tile_27_12_to_tile_27_13_1;
	wire horizontal_tile_27_12_to_tile_27_13_2;
	wire horizontal_tile_27_12_to_tile_27_13_3;
	wire horizontal_tile_27_13_to_tile_27_12_0;
	wire horizontal_tile_27_13_to_tile_27_12_1;
	wire horizontal_tile_27_13_to_tile_27_12_2;
	wire horizontal_tile_27_13_to_tile_27_12_3;

	wire horizontal_tile_28_12_to_tile_28_13_0;
	wire horizontal_tile_28_12_to_tile_28_13_1;
	wire horizontal_tile_28_12_to_tile_28_13_2;
	wire horizontal_tile_28_12_to_tile_28_13_3;
	wire horizontal_tile_28_13_to_tile_28_12_0;
	wire horizontal_tile_28_13_to_tile_28_12_1;
	wire horizontal_tile_28_13_to_tile_28_12_2;
	wire horizontal_tile_28_13_to_tile_28_12_3;

	wire horizontal_tile_29_12_to_tile_29_13_0;
	wire horizontal_tile_29_12_to_tile_29_13_1;
	wire horizontal_tile_29_12_to_tile_29_13_2;
	wire horizontal_tile_29_12_to_tile_29_13_3;
	wire horizontal_tile_29_13_to_tile_29_12_0;
	wire horizontal_tile_29_13_to_tile_29_12_1;
	wire horizontal_tile_29_13_to_tile_29_12_2;
	wire horizontal_tile_29_13_to_tile_29_12_3;

	wire horizontal_tile_30_12_to_tile_30_13_0;
	wire horizontal_tile_30_12_to_tile_30_13_1;
	wire horizontal_tile_30_12_to_tile_30_13_2;
	wire horizontal_tile_30_12_to_tile_30_13_3;
	wire horizontal_tile_30_13_to_tile_30_12_0;
	wire horizontal_tile_30_13_to_tile_30_12_1;
	wire horizontal_tile_30_13_to_tile_30_12_2;
	wire horizontal_tile_30_13_to_tile_30_12_3;

	wire horizontal_tile_31_12_to_tile_31_13_0;
	wire horizontal_tile_31_12_to_tile_31_13_1;
	wire horizontal_tile_31_12_to_tile_31_13_2;
	wire horizontal_tile_31_12_to_tile_31_13_3;
	wire horizontal_tile_31_13_to_tile_31_12_0;
	wire horizontal_tile_31_13_to_tile_31_12_1;
	wire horizontal_tile_31_13_to_tile_31_12_2;
	wire horizontal_tile_31_13_to_tile_31_12_3;

	wire horizontal_tile_0_13_to_tile_0_14_0;
	wire horizontal_tile_0_13_to_tile_0_14_1;
	wire horizontal_tile_0_13_to_tile_0_14_2;
	wire horizontal_tile_0_13_to_tile_0_14_3;
	wire horizontal_tile_0_14_to_tile_0_13_0;
	wire horizontal_tile_0_14_to_tile_0_13_1;
	wire horizontal_tile_0_14_to_tile_0_13_2;
	wire horizontal_tile_0_14_to_tile_0_13_3;

	wire horizontal_tile_1_13_to_tile_1_14_0;
	wire horizontal_tile_1_13_to_tile_1_14_1;
	wire horizontal_tile_1_13_to_tile_1_14_2;
	wire horizontal_tile_1_13_to_tile_1_14_3;
	wire horizontal_tile_1_14_to_tile_1_13_0;
	wire horizontal_tile_1_14_to_tile_1_13_1;
	wire horizontal_tile_1_14_to_tile_1_13_2;
	wire horizontal_tile_1_14_to_tile_1_13_3;

	wire horizontal_tile_2_13_to_tile_2_14_0;
	wire horizontal_tile_2_13_to_tile_2_14_1;
	wire horizontal_tile_2_13_to_tile_2_14_2;
	wire horizontal_tile_2_13_to_tile_2_14_3;
	wire horizontal_tile_2_14_to_tile_2_13_0;
	wire horizontal_tile_2_14_to_tile_2_13_1;
	wire horizontal_tile_2_14_to_tile_2_13_2;
	wire horizontal_tile_2_14_to_tile_2_13_3;

	wire horizontal_tile_3_13_to_tile_3_14_0;
	wire horizontal_tile_3_13_to_tile_3_14_1;
	wire horizontal_tile_3_13_to_tile_3_14_2;
	wire horizontal_tile_3_13_to_tile_3_14_3;
	wire horizontal_tile_3_14_to_tile_3_13_0;
	wire horizontal_tile_3_14_to_tile_3_13_1;
	wire horizontal_tile_3_14_to_tile_3_13_2;
	wire horizontal_tile_3_14_to_tile_3_13_3;

	wire horizontal_tile_4_13_to_tile_4_14_0;
	wire horizontal_tile_4_13_to_tile_4_14_1;
	wire horizontal_tile_4_13_to_tile_4_14_2;
	wire horizontal_tile_4_13_to_tile_4_14_3;
	wire horizontal_tile_4_14_to_tile_4_13_0;
	wire horizontal_tile_4_14_to_tile_4_13_1;
	wire horizontal_tile_4_14_to_tile_4_13_2;
	wire horizontal_tile_4_14_to_tile_4_13_3;

	wire horizontal_tile_5_13_to_tile_5_14_0;
	wire horizontal_tile_5_13_to_tile_5_14_1;
	wire horizontal_tile_5_13_to_tile_5_14_2;
	wire horizontal_tile_5_13_to_tile_5_14_3;
	wire horizontal_tile_5_14_to_tile_5_13_0;
	wire horizontal_tile_5_14_to_tile_5_13_1;
	wire horizontal_tile_5_14_to_tile_5_13_2;
	wire horizontal_tile_5_14_to_tile_5_13_3;

	wire horizontal_tile_6_13_to_tile_6_14_0;
	wire horizontal_tile_6_13_to_tile_6_14_1;
	wire horizontal_tile_6_13_to_tile_6_14_2;
	wire horizontal_tile_6_13_to_tile_6_14_3;
	wire horizontal_tile_6_14_to_tile_6_13_0;
	wire horizontal_tile_6_14_to_tile_6_13_1;
	wire horizontal_tile_6_14_to_tile_6_13_2;
	wire horizontal_tile_6_14_to_tile_6_13_3;

	wire horizontal_tile_7_13_to_tile_7_14_0;
	wire horizontal_tile_7_13_to_tile_7_14_1;
	wire horizontal_tile_7_13_to_tile_7_14_2;
	wire horizontal_tile_7_13_to_tile_7_14_3;
	wire horizontal_tile_7_14_to_tile_7_13_0;
	wire horizontal_tile_7_14_to_tile_7_13_1;
	wire horizontal_tile_7_14_to_tile_7_13_2;
	wire horizontal_tile_7_14_to_tile_7_13_3;

	wire horizontal_tile_8_13_to_tile_8_14_0;
	wire horizontal_tile_8_13_to_tile_8_14_1;
	wire horizontal_tile_8_13_to_tile_8_14_2;
	wire horizontal_tile_8_13_to_tile_8_14_3;
	wire horizontal_tile_8_14_to_tile_8_13_0;
	wire horizontal_tile_8_14_to_tile_8_13_1;
	wire horizontal_tile_8_14_to_tile_8_13_2;
	wire horizontal_tile_8_14_to_tile_8_13_3;

	wire horizontal_tile_9_13_to_tile_9_14_0;
	wire horizontal_tile_9_13_to_tile_9_14_1;
	wire horizontal_tile_9_13_to_tile_9_14_2;
	wire horizontal_tile_9_13_to_tile_9_14_3;
	wire horizontal_tile_9_14_to_tile_9_13_0;
	wire horizontal_tile_9_14_to_tile_9_13_1;
	wire horizontal_tile_9_14_to_tile_9_13_2;
	wire horizontal_tile_9_14_to_tile_9_13_3;

	wire horizontal_tile_10_13_to_tile_10_14_0;
	wire horizontal_tile_10_13_to_tile_10_14_1;
	wire horizontal_tile_10_13_to_tile_10_14_2;
	wire horizontal_tile_10_13_to_tile_10_14_3;
	wire horizontal_tile_10_14_to_tile_10_13_0;
	wire horizontal_tile_10_14_to_tile_10_13_1;
	wire horizontal_tile_10_14_to_tile_10_13_2;
	wire horizontal_tile_10_14_to_tile_10_13_3;

	wire horizontal_tile_11_13_to_tile_11_14_0;
	wire horizontal_tile_11_13_to_tile_11_14_1;
	wire horizontal_tile_11_13_to_tile_11_14_2;
	wire horizontal_tile_11_13_to_tile_11_14_3;
	wire horizontal_tile_11_14_to_tile_11_13_0;
	wire horizontal_tile_11_14_to_tile_11_13_1;
	wire horizontal_tile_11_14_to_tile_11_13_2;
	wire horizontal_tile_11_14_to_tile_11_13_3;

	wire horizontal_tile_12_13_to_tile_12_14_0;
	wire horizontal_tile_12_13_to_tile_12_14_1;
	wire horizontal_tile_12_13_to_tile_12_14_2;
	wire horizontal_tile_12_13_to_tile_12_14_3;
	wire horizontal_tile_12_14_to_tile_12_13_0;
	wire horizontal_tile_12_14_to_tile_12_13_1;
	wire horizontal_tile_12_14_to_tile_12_13_2;
	wire horizontal_tile_12_14_to_tile_12_13_3;

	wire horizontal_tile_13_13_to_tile_13_14_0;
	wire horizontal_tile_13_13_to_tile_13_14_1;
	wire horizontal_tile_13_13_to_tile_13_14_2;
	wire horizontal_tile_13_13_to_tile_13_14_3;
	wire horizontal_tile_13_14_to_tile_13_13_0;
	wire horizontal_tile_13_14_to_tile_13_13_1;
	wire horizontal_tile_13_14_to_tile_13_13_2;
	wire horizontal_tile_13_14_to_tile_13_13_3;

	wire horizontal_tile_14_13_to_tile_14_14_0;
	wire horizontal_tile_14_13_to_tile_14_14_1;
	wire horizontal_tile_14_13_to_tile_14_14_2;
	wire horizontal_tile_14_13_to_tile_14_14_3;
	wire horizontal_tile_14_14_to_tile_14_13_0;
	wire horizontal_tile_14_14_to_tile_14_13_1;
	wire horizontal_tile_14_14_to_tile_14_13_2;
	wire horizontal_tile_14_14_to_tile_14_13_3;

	wire horizontal_tile_15_13_to_tile_15_14_0;
	wire horizontal_tile_15_13_to_tile_15_14_1;
	wire horizontal_tile_15_13_to_tile_15_14_2;
	wire horizontal_tile_15_13_to_tile_15_14_3;
	wire horizontal_tile_15_14_to_tile_15_13_0;
	wire horizontal_tile_15_14_to_tile_15_13_1;
	wire horizontal_tile_15_14_to_tile_15_13_2;
	wire horizontal_tile_15_14_to_tile_15_13_3;

	wire horizontal_tile_16_13_to_tile_16_14_0;
	wire horizontal_tile_16_13_to_tile_16_14_1;
	wire horizontal_tile_16_13_to_tile_16_14_2;
	wire horizontal_tile_16_13_to_tile_16_14_3;
	wire horizontal_tile_16_14_to_tile_16_13_0;
	wire horizontal_tile_16_14_to_tile_16_13_1;
	wire horizontal_tile_16_14_to_tile_16_13_2;
	wire horizontal_tile_16_14_to_tile_16_13_3;

	wire horizontal_tile_17_13_to_tile_17_14_0;
	wire horizontal_tile_17_13_to_tile_17_14_1;
	wire horizontal_tile_17_13_to_tile_17_14_2;
	wire horizontal_tile_17_13_to_tile_17_14_3;
	wire horizontal_tile_17_14_to_tile_17_13_0;
	wire horizontal_tile_17_14_to_tile_17_13_1;
	wire horizontal_tile_17_14_to_tile_17_13_2;
	wire horizontal_tile_17_14_to_tile_17_13_3;

	wire horizontal_tile_18_13_to_tile_18_14_0;
	wire horizontal_tile_18_13_to_tile_18_14_1;
	wire horizontal_tile_18_13_to_tile_18_14_2;
	wire horizontal_tile_18_13_to_tile_18_14_3;
	wire horizontal_tile_18_14_to_tile_18_13_0;
	wire horizontal_tile_18_14_to_tile_18_13_1;
	wire horizontal_tile_18_14_to_tile_18_13_2;
	wire horizontal_tile_18_14_to_tile_18_13_3;

	wire horizontal_tile_19_13_to_tile_19_14_0;
	wire horizontal_tile_19_13_to_tile_19_14_1;
	wire horizontal_tile_19_13_to_tile_19_14_2;
	wire horizontal_tile_19_13_to_tile_19_14_3;
	wire horizontal_tile_19_14_to_tile_19_13_0;
	wire horizontal_tile_19_14_to_tile_19_13_1;
	wire horizontal_tile_19_14_to_tile_19_13_2;
	wire horizontal_tile_19_14_to_tile_19_13_3;

	wire horizontal_tile_20_13_to_tile_20_14_0;
	wire horizontal_tile_20_13_to_tile_20_14_1;
	wire horizontal_tile_20_13_to_tile_20_14_2;
	wire horizontal_tile_20_13_to_tile_20_14_3;
	wire horizontal_tile_20_14_to_tile_20_13_0;
	wire horizontal_tile_20_14_to_tile_20_13_1;
	wire horizontal_tile_20_14_to_tile_20_13_2;
	wire horizontal_tile_20_14_to_tile_20_13_3;

	wire horizontal_tile_21_13_to_tile_21_14_0;
	wire horizontal_tile_21_13_to_tile_21_14_1;
	wire horizontal_tile_21_13_to_tile_21_14_2;
	wire horizontal_tile_21_13_to_tile_21_14_3;
	wire horizontal_tile_21_14_to_tile_21_13_0;
	wire horizontal_tile_21_14_to_tile_21_13_1;
	wire horizontal_tile_21_14_to_tile_21_13_2;
	wire horizontal_tile_21_14_to_tile_21_13_3;

	wire horizontal_tile_22_13_to_tile_22_14_0;
	wire horizontal_tile_22_13_to_tile_22_14_1;
	wire horizontal_tile_22_13_to_tile_22_14_2;
	wire horizontal_tile_22_13_to_tile_22_14_3;
	wire horizontal_tile_22_14_to_tile_22_13_0;
	wire horizontal_tile_22_14_to_tile_22_13_1;
	wire horizontal_tile_22_14_to_tile_22_13_2;
	wire horizontal_tile_22_14_to_tile_22_13_3;

	wire horizontal_tile_23_13_to_tile_23_14_0;
	wire horizontal_tile_23_13_to_tile_23_14_1;
	wire horizontal_tile_23_13_to_tile_23_14_2;
	wire horizontal_tile_23_13_to_tile_23_14_3;
	wire horizontal_tile_23_14_to_tile_23_13_0;
	wire horizontal_tile_23_14_to_tile_23_13_1;
	wire horizontal_tile_23_14_to_tile_23_13_2;
	wire horizontal_tile_23_14_to_tile_23_13_3;

	wire horizontal_tile_24_13_to_tile_24_14_0;
	wire horizontal_tile_24_13_to_tile_24_14_1;
	wire horizontal_tile_24_13_to_tile_24_14_2;
	wire horizontal_tile_24_13_to_tile_24_14_3;
	wire horizontal_tile_24_14_to_tile_24_13_0;
	wire horizontal_tile_24_14_to_tile_24_13_1;
	wire horizontal_tile_24_14_to_tile_24_13_2;
	wire horizontal_tile_24_14_to_tile_24_13_3;

	wire horizontal_tile_25_13_to_tile_25_14_0;
	wire horizontal_tile_25_13_to_tile_25_14_1;
	wire horizontal_tile_25_13_to_tile_25_14_2;
	wire horizontal_tile_25_13_to_tile_25_14_3;
	wire horizontal_tile_25_14_to_tile_25_13_0;
	wire horizontal_tile_25_14_to_tile_25_13_1;
	wire horizontal_tile_25_14_to_tile_25_13_2;
	wire horizontal_tile_25_14_to_tile_25_13_3;

	wire horizontal_tile_26_13_to_tile_26_14_0;
	wire horizontal_tile_26_13_to_tile_26_14_1;
	wire horizontal_tile_26_13_to_tile_26_14_2;
	wire horizontal_tile_26_13_to_tile_26_14_3;
	wire horizontal_tile_26_14_to_tile_26_13_0;
	wire horizontal_tile_26_14_to_tile_26_13_1;
	wire horizontal_tile_26_14_to_tile_26_13_2;
	wire horizontal_tile_26_14_to_tile_26_13_3;

	wire horizontal_tile_27_13_to_tile_27_14_0;
	wire horizontal_tile_27_13_to_tile_27_14_1;
	wire horizontal_tile_27_13_to_tile_27_14_2;
	wire horizontal_tile_27_13_to_tile_27_14_3;
	wire horizontal_tile_27_14_to_tile_27_13_0;
	wire horizontal_tile_27_14_to_tile_27_13_1;
	wire horizontal_tile_27_14_to_tile_27_13_2;
	wire horizontal_tile_27_14_to_tile_27_13_3;

	wire horizontal_tile_28_13_to_tile_28_14_0;
	wire horizontal_tile_28_13_to_tile_28_14_1;
	wire horizontal_tile_28_13_to_tile_28_14_2;
	wire horizontal_tile_28_13_to_tile_28_14_3;
	wire horizontal_tile_28_14_to_tile_28_13_0;
	wire horizontal_tile_28_14_to_tile_28_13_1;
	wire horizontal_tile_28_14_to_tile_28_13_2;
	wire horizontal_tile_28_14_to_tile_28_13_3;

	wire horizontal_tile_29_13_to_tile_29_14_0;
	wire horizontal_tile_29_13_to_tile_29_14_1;
	wire horizontal_tile_29_13_to_tile_29_14_2;
	wire horizontal_tile_29_13_to_tile_29_14_3;
	wire horizontal_tile_29_14_to_tile_29_13_0;
	wire horizontal_tile_29_14_to_tile_29_13_1;
	wire horizontal_tile_29_14_to_tile_29_13_2;
	wire horizontal_tile_29_14_to_tile_29_13_3;

	wire horizontal_tile_30_13_to_tile_30_14_0;
	wire horizontal_tile_30_13_to_tile_30_14_1;
	wire horizontal_tile_30_13_to_tile_30_14_2;
	wire horizontal_tile_30_13_to_tile_30_14_3;
	wire horizontal_tile_30_14_to_tile_30_13_0;
	wire horizontal_tile_30_14_to_tile_30_13_1;
	wire horizontal_tile_30_14_to_tile_30_13_2;
	wire horizontal_tile_30_14_to_tile_30_13_3;

	wire horizontal_tile_31_13_to_tile_31_14_0;
	wire horizontal_tile_31_13_to_tile_31_14_1;
	wire horizontal_tile_31_13_to_tile_31_14_2;
	wire horizontal_tile_31_13_to_tile_31_14_3;
	wire horizontal_tile_31_14_to_tile_31_13_0;
	wire horizontal_tile_31_14_to_tile_31_13_1;
	wire horizontal_tile_31_14_to_tile_31_13_2;
	wire horizontal_tile_31_14_to_tile_31_13_3;

	wire horizontal_tile_0_14_to_tile_0_15_0;
	wire horizontal_tile_0_14_to_tile_0_15_1;
	wire horizontal_tile_0_14_to_tile_0_15_2;
	wire horizontal_tile_0_14_to_tile_0_15_3;
	wire horizontal_tile_0_15_to_tile_0_14_0;
	wire horizontal_tile_0_15_to_tile_0_14_1;
	wire horizontal_tile_0_15_to_tile_0_14_2;
	wire horizontal_tile_0_15_to_tile_0_14_3;

	wire horizontal_tile_1_14_to_tile_1_15_0;
	wire horizontal_tile_1_14_to_tile_1_15_1;
	wire horizontal_tile_1_14_to_tile_1_15_2;
	wire horizontal_tile_1_14_to_tile_1_15_3;
	wire horizontal_tile_1_15_to_tile_1_14_0;
	wire horizontal_tile_1_15_to_tile_1_14_1;
	wire horizontal_tile_1_15_to_tile_1_14_2;
	wire horizontal_tile_1_15_to_tile_1_14_3;

	wire horizontal_tile_2_14_to_tile_2_15_0;
	wire horizontal_tile_2_14_to_tile_2_15_1;
	wire horizontal_tile_2_14_to_tile_2_15_2;
	wire horizontal_tile_2_14_to_tile_2_15_3;
	wire horizontal_tile_2_15_to_tile_2_14_0;
	wire horizontal_tile_2_15_to_tile_2_14_1;
	wire horizontal_tile_2_15_to_tile_2_14_2;
	wire horizontal_tile_2_15_to_tile_2_14_3;

	wire horizontal_tile_3_14_to_tile_3_15_0;
	wire horizontal_tile_3_14_to_tile_3_15_1;
	wire horizontal_tile_3_14_to_tile_3_15_2;
	wire horizontal_tile_3_14_to_tile_3_15_3;
	wire horizontal_tile_3_15_to_tile_3_14_0;
	wire horizontal_tile_3_15_to_tile_3_14_1;
	wire horizontal_tile_3_15_to_tile_3_14_2;
	wire horizontal_tile_3_15_to_tile_3_14_3;

	wire horizontal_tile_4_14_to_tile_4_15_0;
	wire horizontal_tile_4_14_to_tile_4_15_1;
	wire horizontal_tile_4_14_to_tile_4_15_2;
	wire horizontal_tile_4_14_to_tile_4_15_3;
	wire horizontal_tile_4_15_to_tile_4_14_0;
	wire horizontal_tile_4_15_to_tile_4_14_1;
	wire horizontal_tile_4_15_to_tile_4_14_2;
	wire horizontal_tile_4_15_to_tile_4_14_3;

	wire horizontal_tile_5_14_to_tile_5_15_0;
	wire horizontal_tile_5_14_to_tile_5_15_1;
	wire horizontal_tile_5_14_to_tile_5_15_2;
	wire horizontal_tile_5_14_to_tile_5_15_3;
	wire horizontal_tile_5_15_to_tile_5_14_0;
	wire horizontal_tile_5_15_to_tile_5_14_1;
	wire horizontal_tile_5_15_to_tile_5_14_2;
	wire horizontal_tile_5_15_to_tile_5_14_3;

	wire horizontal_tile_6_14_to_tile_6_15_0;
	wire horizontal_tile_6_14_to_tile_6_15_1;
	wire horizontal_tile_6_14_to_tile_6_15_2;
	wire horizontal_tile_6_14_to_tile_6_15_3;
	wire horizontal_tile_6_15_to_tile_6_14_0;
	wire horizontal_tile_6_15_to_tile_6_14_1;
	wire horizontal_tile_6_15_to_tile_6_14_2;
	wire horizontal_tile_6_15_to_tile_6_14_3;

	wire horizontal_tile_7_14_to_tile_7_15_0;
	wire horizontal_tile_7_14_to_tile_7_15_1;
	wire horizontal_tile_7_14_to_tile_7_15_2;
	wire horizontal_tile_7_14_to_tile_7_15_3;
	wire horizontal_tile_7_15_to_tile_7_14_0;
	wire horizontal_tile_7_15_to_tile_7_14_1;
	wire horizontal_tile_7_15_to_tile_7_14_2;
	wire horizontal_tile_7_15_to_tile_7_14_3;

	wire horizontal_tile_8_14_to_tile_8_15_0;
	wire horizontal_tile_8_14_to_tile_8_15_1;
	wire horizontal_tile_8_14_to_tile_8_15_2;
	wire horizontal_tile_8_14_to_tile_8_15_3;
	wire horizontal_tile_8_15_to_tile_8_14_0;
	wire horizontal_tile_8_15_to_tile_8_14_1;
	wire horizontal_tile_8_15_to_tile_8_14_2;
	wire horizontal_tile_8_15_to_tile_8_14_3;

	wire horizontal_tile_9_14_to_tile_9_15_0;
	wire horizontal_tile_9_14_to_tile_9_15_1;
	wire horizontal_tile_9_14_to_tile_9_15_2;
	wire horizontal_tile_9_14_to_tile_9_15_3;
	wire horizontal_tile_9_15_to_tile_9_14_0;
	wire horizontal_tile_9_15_to_tile_9_14_1;
	wire horizontal_tile_9_15_to_tile_9_14_2;
	wire horizontal_tile_9_15_to_tile_9_14_3;

	wire horizontal_tile_10_14_to_tile_10_15_0;
	wire horizontal_tile_10_14_to_tile_10_15_1;
	wire horizontal_tile_10_14_to_tile_10_15_2;
	wire horizontal_tile_10_14_to_tile_10_15_3;
	wire horizontal_tile_10_15_to_tile_10_14_0;
	wire horizontal_tile_10_15_to_tile_10_14_1;
	wire horizontal_tile_10_15_to_tile_10_14_2;
	wire horizontal_tile_10_15_to_tile_10_14_3;

	wire horizontal_tile_11_14_to_tile_11_15_0;
	wire horizontal_tile_11_14_to_tile_11_15_1;
	wire horizontal_tile_11_14_to_tile_11_15_2;
	wire horizontal_tile_11_14_to_tile_11_15_3;
	wire horizontal_tile_11_15_to_tile_11_14_0;
	wire horizontal_tile_11_15_to_tile_11_14_1;
	wire horizontal_tile_11_15_to_tile_11_14_2;
	wire horizontal_tile_11_15_to_tile_11_14_3;

	wire horizontal_tile_12_14_to_tile_12_15_0;
	wire horizontal_tile_12_14_to_tile_12_15_1;
	wire horizontal_tile_12_14_to_tile_12_15_2;
	wire horizontal_tile_12_14_to_tile_12_15_3;
	wire horizontal_tile_12_15_to_tile_12_14_0;
	wire horizontal_tile_12_15_to_tile_12_14_1;
	wire horizontal_tile_12_15_to_tile_12_14_2;
	wire horizontal_tile_12_15_to_tile_12_14_3;

	wire horizontal_tile_13_14_to_tile_13_15_0;
	wire horizontal_tile_13_14_to_tile_13_15_1;
	wire horizontal_tile_13_14_to_tile_13_15_2;
	wire horizontal_tile_13_14_to_tile_13_15_3;
	wire horizontal_tile_13_15_to_tile_13_14_0;
	wire horizontal_tile_13_15_to_tile_13_14_1;
	wire horizontal_tile_13_15_to_tile_13_14_2;
	wire horizontal_tile_13_15_to_tile_13_14_3;

	wire horizontal_tile_14_14_to_tile_14_15_0;
	wire horizontal_tile_14_14_to_tile_14_15_1;
	wire horizontal_tile_14_14_to_tile_14_15_2;
	wire horizontal_tile_14_14_to_tile_14_15_3;
	wire horizontal_tile_14_15_to_tile_14_14_0;
	wire horizontal_tile_14_15_to_tile_14_14_1;
	wire horizontal_tile_14_15_to_tile_14_14_2;
	wire horizontal_tile_14_15_to_tile_14_14_3;

	wire horizontal_tile_15_14_to_tile_15_15_0;
	wire horizontal_tile_15_14_to_tile_15_15_1;
	wire horizontal_tile_15_14_to_tile_15_15_2;
	wire horizontal_tile_15_14_to_tile_15_15_3;
	wire horizontal_tile_15_15_to_tile_15_14_0;
	wire horizontal_tile_15_15_to_tile_15_14_1;
	wire horizontal_tile_15_15_to_tile_15_14_2;
	wire horizontal_tile_15_15_to_tile_15_14_3;

	wire horizontal_tile_16_14_to_tile_16_15_0;
	wire horizontal_tile_16_14_to_tile_16_15_1;
	wire horizontal_tile_16_14_to_tile_16_15_2;
	wire horizontal_tile_16_14_to_tile_16_15_3;
	wire horizontal_tile_16_15_to_tile_16_14_0;
	wire horizontal_tile_16_15_to_tile_16_14_1;
	wire horizontal_tile_16_15_to_tile_16_14_2;
	wire horizontal_tile_16_15_to_tile_16_14_3;

	wire horizontal_tile_17_14_to_tile_17_15_0;
	wire horizontal_tile_17_14_to_tile_17_15_1;
	wire horizontal_tile_17_14_to_tile_17_15_2;
	wire horizontal_tile_17_14_to_tile_17_15_3;
	wire horizontal_tile_17_15_to_tile_17_14_0;
	wire horizontal_tile_17_15_to_tile_17_14_1;
	wire horizontal_tile_17_15_to_tile_17_14_2;
	wire horizontal_tile_17_15_to_tile_17_14_3;

	wire horizontal_tile_18_14_to_tile_18_15_0;
	wire horizontal_tile_18_14_to_tile_18_15_1;
	wire horizontal_tile_18_14_to_tile_18_15_2;
	wire horizontal_tile_18_14_to_tile_18_15_3;
	wire horizontal_tile_18_15_to_tile_18_14_0;
	wire horizontal_tile_18_15_to_tile_18_14_1;
	wire horizontal_tile_18_15_to_tile_18_14_2;
	wire horizontal_tile_18_15_to_tile_18_14_3;

	wire horizontal_tile_19_14_to_tile_19_15_0;
	wire horizontal_tile_19_14_to_tile_19_15_1;
	wire horizontal_tile_19_14_to_tile_19_15_2;
	wire horizontal_tile_19_14_to_tile_19_15_3;
	wire horizontal_tile_19_15_to_tile_19_14_0;
	wire horizontal_tile_19_15_to_tile_19_14_1;
	wire horizontal_tile_19_15_to_tile_19_14_2;
	wire horizontal_tile_19_15_to_tile_19_14_3;

	wire horizontal_tile_20_14_to_tile_20_15_0;
	wire horizontal_tile_20_14_to_tile_20_15_1;
	wire horizontal_tile_20_14_to_tile_20_15_2;
	wire horizontal_tile_20_14_to_tile_20_15_3;
	wire horizontal_tile_20_15_to_tile_20_14_0;
	wire horizontal_tile_20_15_to_tile_20_14_1;
	wire horizontal_tile_20_15_to_tile_20_14_2;
	wire horizontal_tile_20_15_to_tile_20_14_3;

	wire horizontal_tile_21_14_to_tile_21_15_0;
	wire horizontal_tile_21_14_to_tile_21_15_1;
	wire horizontal_tile_21_14_to_tile_21_15_2;
	wire horizontal_tile_21_14_to_tile_21_15_3;
	wire horizontal_tile_21_15_to_tile_21_14_0;
	wire horizontal_tile_21_15_to_tile_21_14_1;
	wire horizontal_tile_21_15_to_tile_21_14_2;
	wire horizontal_tile_21_15_to_tile_21_14_3;

	wire horizontal_tile_22_14_to_tile_22_15_0;
	wire horizontal_tile_22_14_to_tile_22_15_1;
	wire horizontal_tile_22_14_to_tile_22_15_2;
	wire horizontal_tile_22_14_to_tile_22_15_3;
	wire horizontal_tile_22_15_to_tile_22_14_0;
	wire horizontal_tile_22_15_to_tile_22_14_1;
	wire horizontal_tile_22_15_to_tile_22_14_2;
	wire horizontal_tile_22_15_to_tile_22_14_3;

	wire horizontal_tile_23_14_to_tile_23_15_0;
	wire horizontal_tile_23_14_to_tile_23_15_1;
	wire horizontal_tile_23_14_to_tile_23_15_2;
	wire horizontal_tile_23_14_to_tile_23_15_3;
	wire horizontal_tile_23_15_to_tile_23_14_0;
	wire horizontal_tile_23_15_to_tile_23_14_1;
	wire horizontal_tile_23_15_to_tile_23_14_2;
	wire horizontal_tile_23_15_to_tile_23_14_3;

	wire horizontal_tile_24_14_to_tile_24_15_0;
	wire horizontal_tile_24_14_to_tile_24_15_1;
	wire horizontal_tile_24_14_to_tile_24_15_2;
	wire horizontal_tile_24_14_to_tile_24_15_3;
	wire horizontal_tile_24_15_to_tile_24_14_0;
	wire horizontal_tile_24_15_to_tile_24_14_1;
	wire horizontal_tile_24_15_to_tile_24_14_2;
	wire horizontal_tile_24_15_to_tile_24_14_3;

	wire horizontal_tile_25_14_to_tile_25_15_0;
	wire horizontal_tile_25_14_to_tile_25_15_1;
	wire horizontal_tile_25_14_to_tile_25_15_2;
	wire horizontal_tile_25_14_to_tile_25_15_3;
	wire horizontal_tile_25_15_to_tile_25_14_0;
	wire horizontal_tile_25_15_to_tile_25_14_1;
	wire horizontal_tile_25_15_to_tile_25_14_2;
	wire horizontal_tile_25_15_to_tile_25_14_3;

	wire horizontal_tile_26_14_to_tile_26_15_0;
	wire horizontal_tile_26_14_to_tile_26_15_1;
	wire horizontal_tile_26_14_to_tile_26_15_2;
	wire horizontal_tile_26_14_to_tile_26_15_3;
	wire horizontal_tile_26_15_to_tile_26_14_0;
	wire horizontal_tile_26_15_to_tile_26_14_1;
	wire horizontal_tile_26_15_to_tile_26_14_2;
	wire horizontal_tile_26_15_to_tile_26_14_3;

	wire horizontal_tile_27_14_to_tile_27_15_0;
	wire horizontal_tile_27_14_to_tile_27_15_1;
	wire horizontal_tile_27_14_to_tile_27_15_2;
	wire horizontal_tile_27_14_to_tile_27_15_3;
	wire horizontal_tile_27_15_to_tile_27_14_0;
	wire horizontal_tile_27_15_to_tile_27_14_1;
	wire horizontal_tile_27_15_to_tile_27_14_2;
	wire horizontal_tile_27_15_to_tile_27_14_3;

	wire horizontal_tile_28_14_to_tile_28_15_0;
	wire horizontal_tile_28_14_to_tile_28_15_1;
	wire horizontal_tile_28_14_to_tile_28_15_2;
	wire horizontal_tile_28_14_to_tile_28_15_3;
	wire horizontal_tile_28_15_to_tile_28_14_0;
	wire horizontal_tile_28_15_to_tile_28_14_1;
	wire horizontal_tile_28_15_to_tile_28_14_2;
	wire horizontal_tile_28_15_to_tile_28_14_3;

	wire horizontal_tile_29_14_to_tile_29_15_0;
	wire horizontal_tile_29_14_to_tile_29_15_1;
	wire horizontal_tile_29_14_to_tile_29_15_2;
	wire horizontal_tile_29_14_to_tile_29_15_3;
	wire horizontal_tile_29_15_to_tile_29_14_0;
	wire horizontal_tile_29_15_to_tile_29_14_1;
	wire horizontal_tile_29_15_to_tile_29_14_2;
	wire horizontal_tile_29_15_to_tile_29_14_3;

	wire horizontal_tile_30_14_to_tile_30_15_0;
	wire horizontal_tile_30_14_to_tile_30_15_1;
	wire horizontal_tile_30_14_to_tile_30_15_2;
	wire horizontal_tile_30_14_to_tile_30_15_3;
	wire horizontal_tile_30_15_to_tile_30_14_0;
	wire horizontal_tile_30_15_to_tile_30_14_1;
	wire horizontal_tile_30_15_to_tile_30_14_2;
	wire horizontal_tile_30_15_to_tile_30_14_3;

	wire horizontal_tile_31_14_to_tile_31_15_0;
	wire horizontal_tile_31_14_to_tile_31_15_1;
	wire horizontal_tile_31_14_to_tile_31_15_2;
	wire horizontal_tile_31_14_to_tile_31_15_3;
	wire horizontal_tile_31_15_to_tile_31_14_0;
	wire horizontal_tile_31_15_to_tile_31_14_1;
	wire horizontal_tile_31_15_to_tile_31_14_2;
	wire horizontal_tile_31_15_to_tile_31_14_3;

	wire horizontal_tile_0_15_to_tile_0_16_0;
	wire horizontal_tile_0_15_to_tile_0_16_1;
	wire horizontal_tile_0_15_to_tile_0_16_2;
	wire horizontal_tile_0_15_to_tile_0_16_3;
	wire horizontal_tile_0_16_to_tile_0_15_0;
	wire horizontal_tile_0_16_to_tile_0_15_1;
	wire horizontal_tile_0_16_to_tile_0_15_2;
	wire horizontal_tile_0_16_to_tile_0_15_3;

	wire horizontal_tile_1_15_to_tile_1_16_0;
	wire horizontal_tile_1_15_to_tile_1_16_1;
	wire horizontal_tile_1_15_to_tile_1_16_2;
	wire horizontal_tile_1_15_to_tile_1_16_3;
	wire horizontal_tile_1_16_to_tile_1_15_0;
	wire horizontal_tile_1_16_to_tile_1_15_1;
	wire horizontal_tile_1_16_to_tile_1_15_2;
	wire horizontal_tile_1_16_to_tile_1_15_3;

	wire horizontal_tile_2_15_to_tile_2_16_0;
	wire horizontal_tile_2_15_to_tile_2_16_1;
	wire horizontal_tile_2_15_to_tile_2_16_2;
	wire horizontal_tile_2_15_to_tile_2_16_3;
	wire horizontal_tile_2_16_to_tile_2_15_0;
	wire horizontal_tile_2_16_to_tile_2_15_1;
	wire horizontal_tile_2_16_to_tile_2_15_2;
	wire horizontal_tile_2_16_to_tile_2_15_3;

	wire horizontal_tile_3_15_to_tile_3_16_0;
	wire horizontal_tile_3_15_to_tile_3_16_1;
	wire horizontal_tile_3_15_to_tile_3_16_2;
	wire horizontal_tile_3_15_to_tile_3_16_3;
	wire horizontal_tile_3_16_to_tile_3_15_0;
	wire horizontal_tile_3_16_to_tile_3_15_1;
	wire horizontal_tile_3_16_to_tile_3_15_2;
	wire horizontal_tile_3_16_to_tile_3_15_3;

	wire horizontal_tile_4_15_to_tile_4_16_0;
	wire horizontal_tile_4_15_to_tile_4_16_1;
	wire horizontal_tile_4_15_to_tile_4_16_2;
	wire horizontal_tile_4_15_to_tile_4_16_3;
	wire horizontal_tile_4_16_to_tile_4_15_0;
	wire horizontal_tile_4_16_to_tile_4_15_1;
	wire horizontal_tile_4_16_to_tile_4_15_2;
	wire horizontal_tile_4_16_to_tile_4_15_3;

	wire horizontal_tile_5_15_to_tile_5_16_0;
	wire horizontal_tile_5_15_to_tile_5_16_1;
	wire horizontal_tile_5_15_to_tile_5_16_2;
	wire horizontal_tile_5_15_to_tile_5_16_3;
	wire horizontal_tile_5_16_to_tile_5_15_0;
	wire horizontal_tile_5_16_to_tile_5_15_1;
	wire horizontal_tile_5_16_to_tile_5_15_2;
	wire horizontal_tile_5_16_to_tile_5_15_3;

	wire horizontal_tile_6_15_to_tile_6_16_0;
	wire horizontal_tile_6_15_to_tile_6_16_1;
	wire horizontal_tile_6_15_to_tile_6_16_2;
	wire horizontal_tile_6_15_to_tile_6_16_3;
	wire horizontal_tile_6_16_to_tile_6_15_0;
	wire horizontal_tile_6_16_to_tile_6_15_1;
	wire horizontal_tile_6_16_to_tile_6_15_2;
	wire horizontal_tile_6_16_to_tile_6_15_3;

	wire horizontal_tile_7_15_to_tile_7_16_0;
	wire horizontal_tile_7_15_to_tile_7_16_1;
	wire horizontal_tile_7_15_to_tile_7_16_2;
	wire horizontal_tile_7_15_to_tile_7_16_3;
	wire horizontal_tile_7_16_to_tile_7_15_0;
	wire horizontal_tile_7_16_to_tile_7_15_1;
	wire horizontal_tile_7_16_to_tile_7_15_2;
	wire horizontal_tile_7_16_to_tile_7_15_3;

	wire horizontal_tile_8_15_to_tile_8_16_0;
	wire horizontal_tile_8_15_to_tile_8_16_1;
	wire horizontal_tile_8_15_to_tile_8_16_2;
	wire horizontal_tile_8_15_to_tile_8_16_3;
	wire horizontal_tile_8_16_to_tile_8_15_0;
	wire horizontal_tile_8_16_to_tile_8_15_1;
	wire horizontal_tile_8_16_to_tile_8_15_2;
	wire horizontal_tile_8_16_to_tile_8_15_3;

	wire horizontal_tile_9_15_to_tile_9_16_0;
	wire horizontal_tile_9_15_to_tile_9_16_1;
	wire horizontal_tile_9_15_to_tile_9_16_2;
	wire horizontal_tile_9_15_to_tile_9_16_3;
	wire horizontal_tile_9_16_to_tile_9_15_0;
	wire horizontal_tile_9_16_to_tile_9_15_1;
	wire horizontal_tile_9_16_to_tile_9_15_2;
	wire horizontal_tile_9_16_to_tile_9_15_3;

	wire horizontal_tile_10_15_to_tile_10_16_0;
	wire horizontal_tile_10_15_to_tile_10_16_1;
	wire horizontal_tile_10_15_to_tile_10_16_2;
	wire horizontal_tile_10_15_to_tile_10_16_3;
	wire horizontal_tile_10_16_to_tile_10_15_0;
	wire horizontal_tile_10_16_to_tile_10_15_1;
	wire horizontal_tile_10_16_to_tile_10_15_2;
	wire horizontal_tile_10_16_to_tile_10_15_3;

	wire horizontal_tile_11_15_to_tile_11_16_0;
	wire horizontal_tile_11_15_to_tile_11_16_1;
	wire horizontal_tile_11_15_to_tile_11_16_2;
	wire horizontal_tile_11_15_to_tile_11_16_3;
	wire horizontal_tile_11_16_to_tile_11_15_0;
	wire horizontal_tile_11_16_to_tile_11_15_1;
	wire horizontal_tile_11_16_to_tile_11_15_2;
	wire horizontal_tile_11_16_to_tile_11_15_3;

	wire horizontal_tile_12_15_to_tile_12_16_0;
	wire horizontal_tile_12_15_to_tile_12_16_1;
	wire horizontal_tile_12_15_to_tile_12_16_2;
	wire horizontal_tile_12_15_to_tile_12_16_3;
	wire horizontal_tile_12_16_to_tile_12_15_0;
	wire horizontal_tile_12_16_to_tile_12_15_1;
	wire horizontal_tile_12_16_to_tile_12_15_2;
	wire horizontal_tile_12_16_to_tile_12_15_3;

	wire horizontal_tile_13_15_to_tile_13_16_0;
	wire horizontal_tile_13_15_to_tile_13_16_1;
	wire horizontal_tile_13_15_to_tile_13_16_2;
	wire horizontal_tile_13_15_to_tile_13_16_3;
	wire horizontal_tile_13_16_to_tile_13_15_0;
	wire horizontal_tile_13_16_to_tile_13_15_1;
	wire horizontal_tile_13_16_to_tile_13_15_2;
	wire horizontal_tile_13_16_to_tile_13_15_3;

	wire horizontal_tile_14_15_to_tile_14_16_0;
	wire horizontal_tile_14_15_to_tile_14_16_1;
	wire horizontal_tile_14_15_to_tile_14_16_2;
	wire horizontal_tile_14_15_to_tile_14_16_3;
	wire horizontal_tile_14_16_to_tile_14_15_0;
	wire horizontal_tile_14_16_to_tile_14_15_1;
	wire horizontal_tile_14_16_to_tile_14_15_2;
	wire horizontal_tile_14_16_to_tile_14_15_3;

	wire horizontal_tile_15_15_to_tile_15_16_0;
	wire horizontal_tile_15_15_to_tile_15_16_1;
	wire horizontal_tile_15_15_to_tile_15_16_2;
	wire horizontal_tile_15_15_to_tile_15_16_3;
	wire horizontal_tile_15_16_to_tile_15_15_0;
	wire horizontal_tile_15_16_to_tile_15_15_1;
	wire horizontal_tile_15_16_to_tile_15_15_2;
	wire horizontal_tile_15_16_to_tile_15_15_3;

	wire horizontal_tile_16_15_to_tile_16_16_0;
	wire horizontal_tile_16_15_to_tile_16_16_1;
	wire horizontal_tile_16_15_to_tile_16_16_2;
	wire horizontal_tile_16_15_to_tile_16_16_3;
	wire horizontal_tile_16_16_to_tile_16_15_0;
	wire horizontal_tile_16_16_to_tile_16_15_1;
	wire horizontal_tile_16_16_to_tile_16_15_2;
	wire horizontal_tile_16_16_to_tile_16_15_3;

	wire horizontal_tile_17_15_to_tile_17_16_0;
	wire horizontal_tile_17_15_to_tile_17_16_1;
	wire horizontal_tile_17_15_to_tile_17_16_2;
	wire horizontal_tile_17_15_to_tile_17_16_3;
	wire horizontal_tile_17_16_to_tile_17_15_0;
	wire horizontal_tile_17_16_to_tile_17_15_1;
	wire horizontal_tile_17_16_to_tile_17_15_2;
	wire horizontal_tile_17_16_to_tile_17_15_3;

	wire horizontal_tile_18_15_to_tile_18_16_0;
	wire horizontal_tile_18_15_to_tile_18_16_1;
	wire horizontal_tile_18_15_to_tile_18_16_2;
	wire horizontal_tile_18_15_to_tile_18_16_3;
	wire horizontal_tile_18_16_to_tile_18_15_0;
	wire horizontal_tile_18_16_to_tile_18_15_1;
	wire horizontal_tile_18_16_to_tile_18_15_2;
	wire horizontal_tile_18_16_to_tile_18_15_3;

	wire horizontal_tile_19_15_to_tile_19_16_0;
	wire horizontal_tile_19_15_to_tile_19_16_1;
	wire horizontal_tile_19_15_to_tile_19_16_2;
	wire horizontal_tile_19_15_to_tile_19_16_3;
	wire horizontal_tile_19_16_to_tile_19_15_0;
	wire horizontal_tile_19_16_to_tile_19_15_1;
	wire horizontal_tile_19_16_to_tile_19_15_2;
	wire horizontal_tile_19_16_to_tile_19_15_3;

	wire horizontal_tile_20_15_to_tile_20_16_0;
	wire horizontal_tile_20_15_to_tile_20_16_1;
	wire horizontal_tile_20_15_to_tile_20_16_2;
	wire horizontal_tile_20_15_to_tile_20_16_3;
	wire horizontal_tile_20_16_to_tile_20_15_0;
	wire horizontal_tile_20_16_to_tile_20_15_1;
	wire horizontal_tile_20_16_to_tile_20_15_2;
	wire horizontal_tile_20_16_to_tile_20_15_3;

	wire horizontal_tile_21_15_to_tile_21_16_0;
	wire horizontal_tile_21_15_to_tile_21_16_1;
	wire horizontal_tile_21_15_to_tile_21_16_2;
	wire horizontal_tile_21_15_to_tile_21_16_3;
	wire horizontal_tile_21_16_to_tile_21_15_0;
	wire horizontal_tile_21_16_to_tile_21_15_1;
	wire horizontal_tile_21_16_to_tile_21_15_2;
	wire horizontal_tile_21_16_to_tile_21_15_3;

	wire horizontal_tile_22_15_to_tile_22_16_0;
	wire horizontal_tile_22_15_to_tile_22_16_1;
	wire horizontal_tile_22_15_to_tile_22_16_2;
	wire horizontal_tile_22_15_to_tile_22_16_3;
	wire horizontal_tile_22_16_to_tile_22_15_0;
	wire horizontal_tile_22_16_to_tile_22_15_1;
	wire horizontal_tile_22_16_to_tile_22_15_2;
	wire horizontal_tile_22_16_to_tile_22_15_3;

	wire horizontal_tile_23_15_to_tile_23_16_0;
	wire horizontal_tile_23_15_to_tile_23_16_1;
	wire horizontal_tile_23_15_to_tile_23_16_2;
	wire horizontal_tile_23_15_to_tile_23_16_3;
	wire horizontal_tile_23_16_to_tile_23_15_0;
	wire horizontal_tile_23_16_to_tile_23_15_1;
	wire horizontal_tile_23_16_to_tile_23_15_2;
	wire horizontal_tile_23_16_to_tile_23_15_3;

	wire horizontal_tile_24_15_to_tile_24_16_0;
	wire horizontal_tile_24_15_to_tile_24_16_1;
	wire horizontal_tile_24_15_to_tile_24_16_2;
	wire horizontal_tile_24_15_to_tile_24_16_3;
	wire horizontal_tile_24_16_to_tile_24_15_0;
	wire horizontal_tile_24_16_to_tile_24_15_1;
	wire horizontal_tile_24_16_to_tile_24_15_2;
	wire horizontal_tile_24_16_to_tile_24_15_3;

	wire horizontal_tile_25_15_to_tile_25_16_0;
	wire horizontal_tile_25_15_to_tile_25_16_1;
	wire horizontal_tile_25_15_to_tile_25_16_2;
	wire horizontal_tile_25_15_to_tile_25_16_3;
	wire horizontal_tile_25_16_to_tile_25_15_0;
	wire horizontal_tile_25_16_to_tile_25_15_1;
	wire horizontal_tile_25_16_to_tile_25_15_2;
	wire horizontal_tile_25_16_to_tile_25_15_3;

	wire horizontal_tile_26_15_to_tile_26_16_0;
	wire horizontal_tile_26_15_to_tile_26_16_1;
	wire horizontal_tile_26_15_to_tile_26_16_2;
	wire horizontal_tile_26_15_to_tile_26_16_3;
	wire horizontal_tile_26_16_to_tile_26_15_0;
	wire horizontal_tile_26_16_to_tile_26_15_1;
	wire horizontal_tile_26_16_to_tile_26_15_2;
	wire horizontal_tile_26_16_to_tile_26_15_3;

	wire horizontal_tile_27_15_to_tile_27_16_0;
	wire horizontal_tile_27_15_to_tile_27_16_1;
	wire horizontal_tile_27_15_to_tile_27_16_2;
	wire horizontal_tile_27_15_to_tile_27_16_3;
	wire horizontal_tile_27_16_to_tile_27_15_0;
	wire horizontal_tile_27_16_to_tile_27_15_1;
	wire horizontal_tile_27_16_to_tile_27_15_2;
	wire horizontal_tile_27_16_to_tile_27_15_3;

	wire horizontal_tile_28_15_to_tile_28_16_0;
	wire horizontal_tile_28_15_to_tile_28_16_1;
	wire horizontal_tile_28_15_to_tile_28_16_2;
	wire horizontal_tile_28_15_to_tile_28_16_3;
	wire horizontal_tile_28_16_to_tile_28_15_0;
	wire horizontal_tile_28_16_to_tile_28_15_1;
	wire horizontal_tile_28_16_to_tile_28_15_2;
	wire horizontal_tile_28_16_to_tile_28_15_3;

	wire horizontal_tile_29_15_to_tile_29_16_0;
	wire horizontal_tile_29_15_to_tile_29_16_1;
	wire horizontal_tile_29_15_to_tile_29_16_2;
	wire horizontal_tile_29_15_to_tile_29_16_3;
	wire horizontal_tile_29_16_to_tile_29_15_0;
	wire horizontal_tile_29_16_to_tile_29_15_1;
	wire horizontal_tile_29_16_to_tile_29_15_2;
	wire horizontal_tile_29_16_to_tile_29_15_3;

	wire horizontal_tile_30_15_to_tile_30_16_0;
	wire horizontal_tile_30_15_to_tile_30_16_1;
	wire horizontal_tile_30_15_to_tile_30_16_2;
	wire horizontal_tile_30_15_to_tile_30_16_3;
	wire horizontal_tile_30_16_to_tile_30_15_0;
	wire horizontal_tile_30_16_to_tile_30_15_1;
	wire horizontal_tile_30_16_to_tile_30_15_2;
	wire horizontal_tile_30_16_to_tile_30_15_3;

	wire horizontal_tile_31_15_to_tile_31_16_0;
	wire horizontal_tile_31_15_to_tile_31_16_1;
	wire horizontal_tile_31_15_to_tile_31_16_2;
	wire horizontal_tile_31_15_to_tile_31_16_3;
	wire horizontal_tile_31_16_to_tile_31_15_0;
	wire horizontal_tile_31_16_to_tile_31_15_1;
	wire horizontal_tile_31_16_to_tile_31_15_2;
	wire horizontal_tile_31_16_to_tile_31_15_3;

	wire horizontal_tile_0_16_to_tile_0_17_0;
	wire horizontal_tile_0_16_to_tile_0_17_1;
	wire horizontal_tile_0_16_to_tile_0_17_2;
	wire horizontal_tile_0_16_to_tile_0_17_3;
	wire horizontal_tile_0_17_to_tile_0_16_0;
	wire horizontal_tile_0_17_to_tile_0_16_1;
	wire horizontal_tile_0_17_to_tile_0_16_2;
	wire horizontal_tile_0_17_to_tile_0_16_3;

	wire horizontal_tile_1_16_to_tile_1_17_0;
	wire horizontal_tile_1_16_to_tile_1_17_1;
	wire horizontal_tile_1_16_to_tile_1_17_2;
	wire horizontal_tile_1_16_to_tile_1_17_3;
	wire horizontal_tile_1_17_to_tile_1_16_0;
	wire horizontal_tile_1_17_to_tile_1_16_1;
	wire horizontal_tile_1_17_to_tile_1_16_2;
	wire horizontal_tile_1_17_to_tile_1_16_3;

	wire horizontal_tile_2_16_to_tile_2_17_0;
	wire horizontal_tile_2_16_to_tile_2_17_1;
	wire horizontal_tile_2_16_to_tile_2_17_2;
	wire horizontal_tile_2_16_to_tile_2_17_3;
	wire horizontal_tile_2_17_to_tile_2_16_0;
	wire horizontal_tile_2_17_to_tile_2_16_1;
	wire horizontal_tile_2_17_to_tile_2_16_2;
	wire horizontal_tile_2_17_to_tile_2_16_3;

	wire horizontal_tile_3_16_to_tile_3_17_0;
	wire horizontal_tile_3_16_to_tile_3_17_1;
	wire horizontal_tile_3_16_to_tile_3_17_2;
	wire horizontal_tile_3_16_to_tile_3_17_3;
	wire horizontal_tile_3_17_to_tile_3_16_0;
	wire horizontal_tile_3_17_to_tile_3_16_1;
	wire horizontal_tile_3_17_to_tile_3_16_2;
	wire horizontal_tile_3_17_to_tile_3_16_3;

	wire horizontal_tile_4_16_to_tile_4_17_0;
	wire horizontal_tile_4_16_to_tile_4_17_1;
	wire horizontal_tile_4_16_to_tile_4_17_2;
	wire horizontal_tile_4_16_to_tile_4_17_3;
	wire horizontal_tile_4_17_to_tile_4_16_0;
	wire horizontal_tile_4_17_to_tile_4_16_1;
	wire horizontal_tile_4_17_to_tile_4_16_2;
	wire horizontal_tile_4_17_to_tile_4_16_3;

	wire horizontal_tile_5_16_to_tile_5_17_0;
	wire horizontal_tile_5_16_to_tile_5_17_1;
	wire horizontal_tile_5_16_to_tile_5_17_2;
	wire horizontal_tile_5_16_to_tile_5_17_3;
	wire horizontal_tile_5_17_to_tile_5_16_0;
	wire horizontal_tile_5_17_to_tile_5_16_1;
	wire horizontal_tile_5_17_to_tile_5_16_2;
	wire horizontal_tile_5_17_to_tile_5_16_3;

	wire horizontal_tile_6_16_to_tile_6_17_0;
	wire horizontal_tile_6_16_to_tile_6_17_1;
	wire horizontal_tile_6_16_to_tile_6_17_2;
	wire horizontal_tile_6_16_to_tile_6_17_3;
	wire horizontal_tile_6_17_to_tile_6_16_0;
	wire horizontal_tile_6_17_to_tile_6_16_1;
	wire horizontal_tile_6_17_to_tile_6_16_2;
	wire horizontal_tile_6_17_to_tile_6_16_3;

	wire horizontal_tile_7_16_to_tile_7_17_0;
	wire horizontal_tile_7_16_to_tile_7_17_1;
	wire horizontal_tile_7_16_to_tile_7_17_2;
	wire horizontal_tile_7_16_to_tile_7_17_3;
	wire horizontal_tile_7_17_to_tile_7_16_0;
	wire horizontal_tile_7_17_to_tile_7_16_1;
	wire horizontal_tile_7_17_to_tile_7_16_2;
	wire horizontal_tile_7_17_to_tile_7_16_3;

	wire horizontal_tile_8_16_to_tile_8_17_0;
	wire horizontal_tile_8_16_to_tile_8_17_1;
	wire horizontal_tile_8_16_to_tile_8_17_2;
	wire horizontal_tile_8_16_to_tile_8_17_3;
	wire horizontal_tile_8_17_to_tile_8_16_0;
	wire horizontal_tile_8_17_to_tile_8_16_1;
	wire horizontal_tile_8_17_to_tile_8_16_2;
	wire horizontal_tile_8_17_to_tile_8_16_3;

	wire horizontal_tile_9_16_to_tile_9_17_0;
	wire horizontal_tile_9_16_to_tile_9_17_1;
	wire horizontal_tile_9_16_to_tile_9_17_2;
	wire horizontal_tile_9_16_to_tile_9_17_3;
	wire horizontal_tile_9_17_to_tile_9_16_0;
	wire horizontal_tile_9_17_to_tile_9_16_1;
	wire horizontal_tile_9_17_to_tile_9_16_2;
	wire horizontal_tile_9_17_to_tile_9_16_3;

	wire horizontal_tile_10_16_to_tile_10_17_0;
	wire horizontal_tile_10_16_to_tile_10_17_1;
	wire horizontal_tile_10_16_to_tile_10_17_2;
	wire horizontal_tile_10_16_to_tile_10_17_3;
	wire horizontal_tile_10_17_to_tile_10_16_0;
	wire horizontal_tile_10_17_to_tile_10_16_1;
	wire horizontal_tile_10_17_to_tile_10_16_2;
	wire horizontal_tile_10_17_to_tile_10_16_3;

	wire horizontal_tile_11_16_to_tile_11_17_0;
	wire horizontal_tile_11_16_to_tile_11_17_1;
	wire horizontal_tile_11_16_to_tile_11_17_2;
	wire horizontal_tile_11_16_to_tile_11_17_3;
	wire horizontal_tile_11_17_to_tile_11_16_0;
	wire horizontal_tile_11_17_to_tile_11_16_1;
	wire horizontal_tile_11_17_to_tile_11_16_2;
	wire horizontal_tile_11_17_to_tile_11_16_3;

	wire horizontal_tile_12_16_to_tile_12_17_0;
	wire horizontal_tile_12_16_to_tile_12_17_1;
	wire horizontal_tile_12_16_to_tile_12_17_2;
	wire horizontal_tile_12_16_to_tile_12_17_3;
	wire horizontal_tile_12_17_to_tile_12_16_0;
	wire horizontal_tile_12_17_to_tile_12_16_1;
	wire horizontal_tile_12_17_to_tile_12_16_2;
	wire horizontal_tile_12_17_to_tile_12_16_3;

	wire horizontal_tile_13_16_to_tile_13_17_0;
	wire horizontal_tile_13_16_to_tile_13_17_1;
	wire horizontal_tile_13_16_to_tile_13_17_2;
	wire horizontal_tile_13_16_to_tile_13_17_3;
	wire horizontal_tile_13_17_to_tile_13_16_0;
	wire horizontal_tile_13_17_to_tile_13_16_1;
	wire horizontal_tile_13_17_to_tile_13_16_2;
	wire horizontal_tile_13_17_to_tile_13_16_3;

	wire horizontal_tile_14_16_to_tile_14_17_0;
	wire horizontal_tile_14_16_to_tile_14_17_1;
	wire horizontal_tile_14_16_to_tile_14_17_2;
	wire horizontal_tile_14_16_to_tile_14_17_3;
	wire horizontal_tile_14_17_to_tile_14_16_0;
	wire horizontal_tile_14_17_to_tile_14_16_1;
	wire horizontal_tile_14_17_to_tile_14_16_2;
	wire horizontal_tile_14_17_to_tile_14_16_3;

	wire horizontal_tile_15_16_to_tile_15_17_0;
	wire horizontal_tile_15_16_to_tile_15_17_1;
	wire horizontal_tile_15_16_to_tile_15_17_2;
	wire horizontal_tile_15_16_to_tile_15_17_3;
	wire horizontal_tile_15_17_to_tile_15_16_0;
	wire horizontal_tile_15_17_to_tile_15_16_1;
	wire horizontal_tile_15_17_to_tile_15_16_2;
	wire horizontal_tile_15_17_to_tile_15_16_3;

	wire horizontal_tile_16_16_to_tile_16_17_0;
	wire horizontal_tile_16_16_to_tile_16_17_1;
	wire horizontal_tile_16_16_to_tile_16_17_2;
	wire horizontal_tile_16_16_to_tile_16_17_3;
	wire horizontal_tile_16_17_to_tile_16_16_0;
	wire horizontal_tile_16_17_to_tile_16_16_1;
	wire horizontal_tile_16_17_to_tile_16_16_2;
	wire horizontal_tile_16_17_to_tile_16_16_3;

	wire horizontal_tile_17_16_to_tile_17_17_0;
	wire horizontal_tile_17_16_to_tile_17_17_1;
	wire horizontal_tile_17_16_to_tile_17_17_2;
	wire horizontal_tile_17_16_to_tile_17_17_3;
	wire horizontal_tile_17_17_to_tile_17_16_0;
	wire horizontal_tile_17_17_to_tile_17_16_1;
	wire horizontal_tile_17_17_to_tile_17_16_2;
	wire horizontal_tile_17_17_to_tile_17_16_3;

	wire horizontal_tile_18_16_to_tile_18_17_0;
	wire horizontal_tile_18_16_to_tile_18_17_1;
	wire horizontal_tile_18_16_to_tile_18_17_2;
	wire horizontal_tile_18_16_to_tile_18_17_3;
	wire horizontal_tile_18_17_to_tile_18_16_0;
	wire horizontal_tile_18_17_to_tile_18_16_1;
	wire horizontal_tile_18_17_to_tile_18_16_2;
	wire horizontal_tile_18_17_to_tile_18_16_3;

	wire horizontal_tile_19_16_to_tile_19_17_0;
	wire horizontal_tile_19_16_to_tile_19_17_1;
	wire horizontal_tile_19_16_to_tile_19_17_2;
	wire horizontal_tile_19_16_to_tile_19_17_3;
	wire horizontal_tile_19_17_to_tile_19_16_0;
	wire horizontal_tile_19_17_to_tile_19_16_1;
	wire horizontal_tile_19_17_to_tile_19_16_2;
	wire horizontal_tile_19_17_to_tile_19_16_3;

	wire horizontal_tile_20_16_to_tile_20_17_0;
	wire horizontal_tile_20_16_to_tile_20_17_1;
	wire horizontal_tile_20_16_to_tile_20_17_2;
	wire horizontal_tile_20_16_to_tile_20_17_3;
	wire horizontal_tile_20_17_to_tile_20_16_0;
	wire horizontal_tile_20_17_to_tile_20_16_1;
	wire horizontal_tile_20_17_to_tile_20_16_2;
	wire horizontal_tile_20_17_to_tile_20_16_3;

	wire horizontal_tile_21_16_to_tile_21_17_0;
	wire horizontal_tile_21_16_to_tile_21_17_1;
	wire horizontal_tile_21_16_to_tile_21_17_2;
	wire horizontal_tile_21_16_to_tile_21_17_3;
	wire horizontal_tile_21_17_to_tile_21_16_0;
	wire horizontal_tile_21_17_to_tile_21_16_1;
	wire horizontal_tile_21_17_to_tile_21_16_2;
	wire horizontal_tile_21_17_to_tile_21_16_3;

	wire horizontal_tile_22_16_to_tile_22_17_0;
	wire horizontal_tile_22_16_to_tile_22_17_1;
	wire horizontal_tile_22_16_to_tile_22_17_2;
	wire horizontal_tile_22_16_to_tile_22_17_3;
	wire horizontal_tile_22_17_to_tile_22_16_0;
	wire horizontal_tile_22_17_to_tile_22_16_1;
	wire horizontal_tile_22_17_to_tile_22_16_2;
	wire horizontal_tile_22_17_to_tile_22_16_3;

	wire horizontal_tile_23_16_to_tile_23_17_0;
	wire horizontal_tile_23_16_to_tile_23_17_1;
	wire horizontal_tile_23_16_to_tile_23_17_2;
	wire horizontal_tile_23_16_to_tile_23_17_3;
	wire horizontal_tile_23_17_to_tile_23_16_0;
	wire horizontal_tile_23_17_to_tile_23_16_1;
	wire horizontal_tile_23_17_to_tile_23_16_2;
	wire horizontal_tile_23_17_to_tile_23_16_3;

	wire horizontal_tile_24_16_to_tile_24_17_0;
	wire horizontal_tile_24_16_to_tile_24_17_1;
	wire horizontal_tile_24_16_to_tile_24_17_2;
	wire horizontal_tile_24_16_to_tile_24_17_3;
	wire horizontal_tile_24_17_to_tile_24_16_0;
	wire horizontal_tile_24_17_to_tile_24_16_1;
	wire horizontal_tile_24_17_to_tile_24_16_2;
	wire horizontal_tile_24_17_to_tile_24_16_3;

	wire horizontal_tile_25_16_to_tile_25_17_0;
	wire horizontal_tile_25_16_to_tile_25_17_1;
	wire horizontal_tile_25_16_to_tile_25_17_2;
	wire horizontal_tile_25_16_to_tile_25_17_3;
	wire horizontal_tile_25_17_to_tile_25_16_0;
	wire horizontal_tile_25_17_to_tile_25_16_1;
	wire horizontal_tile_25_17_to_tile_25_16_2;
	wire horizontal_tile_25_17_to_tile_25_16_3;

	wire horizontal_tile_26_16_to_tile_26_17_0;
	wire horizontal_tile_26_16_to_tile_26_17_1;
	wire horizontal_tile_26_16_to_tile_26_17_2;
	wire horizontal_tile_26_16_to_tile_26_17_3;
	wire horizontal_tile_26_17_to_tile_26_16_0;
	wire horizontal_tile_26_17_to_tile_26_16_1;
	wire horizontal_tile_26_17_to_tile_26_16_2;
	wire horizontal_tile_26_17_to_tile_26_16_3;

	wire horizontal_tile_27_16_to_tile_27_17_0;
	wire horizontal_tile_27_16_to_tile_27_17_1;
	wire horizontal_tile_27_16_to_tile_27_17_2;
	wire horizontal_tile_27_16_to_tile_27_17_3;
	wire horizontal_tile_27_17_to_tile_27_16_0;
	wire horizontal_tile_27_17_to_tile_27_16_1;
	wire horizontal_tile_27_17_to_tile_27_16_2;
	wire horizontal_tile_27_17_to_tile_27_16_3;

	wire horizontal_tile_28_16_to_tile_28_17_0;
	wire horizontal_tile_28_16_to_tile_28_17_1;
	wire horizontal_tile_28_16_to_tile_28_17_2;
	wire horizontal_tile_28_16_to_tile_28_17_3;
	wire horizontal_tile_28_17_to_tile_28_16_0;
	wire horizontal_tile_28_17_to_tile_28_16_1;
	wire horizontal_tile_28_17_to_tile_28_16_2;
	wire horizontal_tile_28_17_to_tile_28_16_3;

	wire horizontal_tile_29_16_to_tile_29_17_0;
	wire horizontal_tile_29_16_to_tile_29_17_1;
	wire horizontal_tile_29_16_to_tile_29_17_2;
	wire horizontal_tile_29_16_to_tile_29_17_3;
	wire horizontal_tile_29_17_to_tile_29_16_0;
	wire horizontal_tile_29_17_to_tile_29_16_1;
	wire horizontal_tile_29_17_to_tile_29_16_2;
	wire horizontal_tile_29_17_to_tile_29_16_3;

	wire horizontal_tile_30_16_to_tile_30_17_0;
	wire horizontal_tile_30_16_to_tile_30_17_1;
	wire horizontal_tile_30_16_to_tile_30_17_2;
	wire horizontal_tile_30_16_to_tile_30_17_3;
	wire horizontal_tile_30_17_to_tile_30_16_0;
	wire horizontal_tile_30_17_to_tile_30_16_1;
	wire horizontal_tile_30_17_to_tile_30_16_2;
	wire horizontal_tile_30_17_to_tile_30_16_3;

	wire horizontal_tile_31_16_to_tile_31_17_0;
	wire horizontal_tile_31_16_to_tile_31_17_1;
	wire horizontal_tile_31_16_to_tile_31_17_2;
	wire horizontal_tile_31_16_to_tile_31_17_3;
	wire horizontal_tile_31_17_to_tile_31_16_0;
	wire horizontal_tile_31_17_to_tile_31_16_1;
	wire horizontal_tile_31_17_to_tile_31_16_2;
	wire horizontal_tile_31_17_to_tile_31_16_3;

	wire horizontal_tile_0_17_to_tile_0_18_0;
	wire horizontal_tile_0_17_to_tile_0_18_1;
	wire horizontal_tile_0_17_to_tile_0_18_2;
	wire horizontal_tile_0_17_to_tile_0_18_3;
	wire horizontal_tile_0_18_to_tile_0_17_0;
	wire horizontal_tile_0_18_to_tile_0_17_1;
	wire horizontal_tile_0_18_to_tile_0_17_2;
	wire horizontal_tile_0_18_to_tile_0_17_3;

	wire horizontal_tile_1_17_to_tile_1_18_0;
	wire horizontal_tile_1_17_to_tile_1_18_1;
	wire horizontal_tile_1_17_to_tile_1_18_2;
	wire horizontal_tile_1_17_to_tile_1_18_3;
	wire horizontal_tile_1_18_to_tile_1_17_0;
	wire horizontal_tile_1_18_to_tile_1_17_1;
	wire horizontal_tile_1_18_to_tile_1_17_2;
	wire horizontal_tile_1_18_to_tile_1_17_3;

	wire horizontal_tile_2_17_to_tile_2_18_0;
	wire horizontal_tile_2_17_to_tile_2_18_1;
	wire horizontal_tile_2_17_to_tile_2_18_2;
	wire horizontal_tile_2_17_to_tile_2_18_3;
	wire horizontal_tile_2_18_to_tile_2_17_0;
	wire horizontal_tile_2_18_to_tile_2_17_1;
	wire horizontal_tile_2_18_to_tile_2_17_2;
	wire horizontal_tile_2_18_to_tile_2_17_3;

	wire horizontal_tile_3_17_to_tile_3_18_0;
	wire horizontal_tile_3_17_to_tile_3_18_1;
	wire horizontal_tile_3_17_to_tile_3_18_2;
	wire horizontal_tile_3_17_to_tile_3_18_3;
	wire horizontal_tile_3_18_to_tile_3_17_0;
	wire horizontal_tile_3_18_to_tile_3_17_1;
	wire horizontal_tile_3_18_to_tile_3_17_2;
	wire horizontal_tile_3_18_to_tile_3_17_3;

	wire horizontal_tile_4_17_to_tile_4_18_0;
	wire horizontal_tile_4_17_to_tile_4_18_1;
	wire horizontal_tile_4_17_to_tile_4_18_2;
	wire horizontal_tile_4_17_to_tile_4_18_3;
	wire horizontal_tile_4_18_to_tile_4_17_0;
	wire horizontal_tile_4_18_to_tile_4_17_1;
	wire horizontal_tile_4_18_to_tile_4_17_2;
	wire horizontal_tile_4_18_to_tile_4_17_3;

	wire horizontal_tile_5_17_to_tile_5_18_0;
	wire horizontal_tile_5_17_to_tile_5_18_1;
	wire horizontal_tile_5_17_to_tile_5_18_2;
	wire horizontal_tile_5_17_to_tile_5_18_3;
	wire horizontal_tile_5_18_to_tile_5_17_0;
	wire horizontal_tile_5_18_to_tile_5_17_1;
	wire horizontal_tile_5_18_to_tile_5_17_2;
	wire horizontal_tile_5_18_to_tile_5_17_3;

	wire horizontal_tile_6_17_to_tile_6_18_0;
	wire horizontal_tile_6_17_to_tile_6_18_1;
	wire horizontal_tile_6_17_to_tile_6_18_2;
	wire horizontal_tile_6_17_to_tile_6_18_3;
	wire horizontal_tile_6_18_to_tile_6_17_0;
	wire horizontal_tile_6_18_to_tile_6_17_1;
	wire horizontal_tile_6_18_to_tile_6_17_2;
	wire horizontal_tile_6_18_to_tile_6_17_3;

	wire horizontal_tile_7_17_to_tile_7_18_0;
	wire horizontal_tile_7_17_to_tile_7_18_1;
	wire horizontal_tile_7_17_to_tile_7_18_2;
	wire horizontal_tile_7_17_to_tile_7_18_3;
	wire horizontal_tile_7_18_to_tile_7_17_0;
	wire horizontal_tile_7_18_to_tile_7_17_1;
	wire horizontal_tile_7_18_to_tile_7_17_2;
	wire horizontal_tile_7_18_to_tile_7_17_3;

	wire horizontal_tile_8_17_to_tile_8_18_0;
	wire horizontal_tile_8_17_to_tile_8_18_1;
	wire horizontal_tile_8_17_to_tile_8_18_2;
	wire horizontal_tile_8_17_to_tile_8_18_3;
	wire horizontal_tile_8_18_to_tile_8_17_0;
	wire horizontal_tile_8_18_to_tile_8_17_1;
	wire horizontal_tile_8_18_to_tile_8_17_2;
	wire horizontal_tile_8_18_to_tile_8_17_3;

	wire horizontal_tile_9_17_to_tile_9_18_0;
	wire horizontal_tile_9_17_to_tile_9_18_1;
	wire horizontal_tile_9_17_to_tile_9_18_2;
	wire horizontal_tile_9_17_to_tile_9_18_3;
	wire horizontal_tile_9_18_to_tile_9_17_0;
	wire horizontal_tile_9_18_to_tile_9_17_1;
	wire horizontal_tile_9_18_to_tile_9_17_2;
	wire horizontal_tile_9_18_to_tile_9_17_3;

	wire horizontal_tile_10_17_to_tile_10_18_0;
	wire horizontal_tile_10_17_to_tile_10_18_1;
	wire horizontal_tile_10_17_to_tile_10_18_2;
	wire horizontal_tile_10_17_to_tile_10_18_3;
	wire horizontal_tile_10_18_to_tile_10_17_0;
	wire horizontal_tile_10_18_to_tile_10_17_1;
	wire horizontal_tile_10_18_to_tile_10_17_2;
	wire horizontal_tile_10_18_to_tile_10_17_3;

	wire horizontal_tile_11_17_to_tile_11_18_0;
	wire horizontal_tile_11_17_to_tile_11_18_1;
	wire horizontal_tile_11_17_to_tile_11_18_2;
	wire horizontal_tile_11_17_to_tile_11_18_3;
	wire horizontal_tile_11_18_to_tile_11_17_0;
	wire horizontal_tile_11_18_to_tile_11_17_1;
	wire horizontal_tile_11_18_to_tile_11_17_2;
	wire horizontal_tile_11_18_to_tile_11_17_3;

	wire horizontal_tile_12_17_to_tile_12_18_0;
	wire horizontal_tile_12_17_to_tile_12_18_1;
	wire horizontal_tile_12_17_to_tile_12_18_2;
	wire horizontal_tile_12_17_to_tile_12_18_3;
	wire horizontal_tile_12_18_to_tile_12_17_0;
	wire horizontal_tile_12_18_to_tile_12_17_1;
	wire horizontal_tile_12_18_to_tile_12_17_2;
	wire horizontal_tile_12_18_to_tile_12_17_3;

	wire horizontal_tile_13_17_to_tile_13_18_0;
	wire horizontal_tile_13_17_to_tile_13_18_1;
	wire horizontal_tile_13_17_to_tile_13_18_2;
	wire horizontal_tile_13_17_to_tile_13_18_3;
	wire horizontal_tile_13_18_to_tile_13_17_0;
	wire horizontal_tile_13_18_to_tile_13_17_1;
	wire horizontal_tile_13_18_to_tile_13_17_2;
	wire horizontal_tile_13_18_to_tile_13_17_3;

	wire horizontal_tile_14_17_to_tile_14_18_0;
	wire horizontal_tile_14_17_to_tile_14_18_1;
	wire horizontal_tile_14_17_to_tile_14_18_2;
	wire horizontal_tile_14_17_to_tile_14_18_3;
	wire horizontal_tile_14_18_to_tile_14_17_0;
	wire horizontal_tile_14_18_to_tile_14_17_1;
	wire horizontal_tile_14_18_to_tile_14_17_2;
	wire horizontal_tile_14_18_to_tile_14_17_3;

	wire horizontal_tile_15_17_to_tile_15_18_0;
	wire horizontal_tile_15_17_to_tile_15_18_1;
	wire horizontal_tile_15_17_to_tile_15_18_2;
	wire horizontal_tile_15_17_to_tile_15_18_3;
	wire horizontal_tile_15_18_to_tile_15_17_0;
	wire horizontal_tile_15_18_to_tile_15_17_1;
	wire horizontal_tile_15_18_to_tile_15_17_2;
	wire horizontal_tile_15_18_to_tile_15_17_3;

	wire horizontal_tile_16_17_to_tile_16_18_0;
	wire horizontal_tile_16_17_to_tile_16_18_1;
	wire horizontal_tile_16_17_to_tile_16_18_2;
	wire horizontal_tile_16_17_to_tile_16_18_3;
	wire horizontal_tile_16_18_to_tile_16_17_0;
	wire horizontal_tile_16_18_to_tile_16_17_1;
	wire horizontal_tile_16_18_to_tile_16_17_2;
	wire horizontal_tile_16_18_to_tile_16_17_3;

	wire horizontal_tile_17_17_to_tile_17_18_0;
	wire horizontal_tile_17_17_to_tile_17_18_1;
	wire horizontal_tile_17_17_to_tile_17_18_2;
	wire horizontal_tile_17_17_to_tile_17_18_3;
	wire horizontal_tile_17_18_to_tile_17_17_0;
	wire horizontal_tile_17_18_to_tile_17_17_1;
	wire horizontal_tile_17_18_to_tile_17_17_2;
	wire horizontal_tile_17_18_to_tile_17_17_3;

	wire horizontal_tile_18_17_to_tile_18_18_0;
	wire horizontal_tile_18_17_to_tile_18_18_1;
	wire horizontal_tile_18_17_to_tile_18_18_2;
	wire horizontal_tile_18_17_to_tile_18_18_3;
	wire horizontal_tile_18_18_to_tile_18_17_0;
	wire horizontal_tile_18_18_to_tile_18_17_1;
	wire horizontal_tile_18_18_to_tile_18_17_2;
	wire horizontal_tile_18_18_to_tile_18_17_3;

	wire horizontal_tile_19_17_to_tile_19_18_0;
	wire horizontal_tile_19_17_to_tile_19_18_1;
	wire horizontal_tile_19_17_to_tile_19_18_2;
	wire horizontal_tile_19_17_to_tile_19_18_3;
	wire horizontal_tile_19_18_to_tile_19_17_0;
	wire horizontal_tile_19_18_to_tile_19_17_1;
	wire horizontal_tile_19_18_to_tile_19_17_2;
	wire horizontal_tile_19_18_to_tile_19_17_3;

	wire horizontal_tile_20_17_to_tile_20_18_0;
	wire horizontal_tile_20_17_to_tile_20_18_1;
	wire horizontal_tile_20_17_to_tile_20_18_2;
	wire horizontal_tile_20_17_to_tile_20_18_3;
	wire horizontal_tile_20_18_to_tile_20_17_0;
	wire horizontal_tile_20_18_to_tile_20_17_1;
	wire horizontal_tile_20_18_to_tile_20_17_2;
	wire horizontal_tile_20_18_to_tile_20_17_3;

	wire horizontal_tile_21_17_to_tile_21_18_0;
	wire horizontal_tile_21_17_to_tile_21_18_1;
	wire horizontal_tile_21_17_to_tile_21_18_2;
	wire horizontal_tile_21_17_to_tile_21_18_3;
	wire horizontal_tile_21_18_to_tile_21_17_0;
	wire horizontal_tile_21_18_to_tile_21_17_1;
	wire horizontal_tile_21_18_to_tile_21_17_2;
	wire horizontal_tile_21_18_to_tile_21_17_3;

	wire horizontal_tile_22_17_to_tile_22_18_0;
	wire horizontal_tile_22_17_to_tile_22_18_1;
	wire horizontal_tile_22_17_to_tile_22_18_2;
	wire horizontal_tile_22_17_to_tile_22_18_3;
	wire horizontal_tile_22_18_to_tile_22_17_0;
	wire horizontal_tile_22_18_to_tile_22_17_1;
	wire horizontal_tile_22_18_to_tile_22_17_2;
	wire horizontal_tile_22_18_to_tile_22_17_3;

	wire horizontal_tile_23_17_to_tile_23_18_0;
	wire horizontal_tile_23_17_to_tile_23_18_1;
	wire horizontal_tile_23_17_to_tile_23_18_2;
	wire horizontal_tile_23_17_to_tile_23_18_3;
	wire horizontal_tile_23_18_to_tile_23_17_0;
	wire horizontal_tile_23_18_to_tile_23_17_1;
	wire horizontal_tile_23_18_to_tile_23_17_2;
	wire horizontal_tile_23_18_to_tile_23_17_3;

	wire horizontal_tile_24_17_to_tile_24_18_0;
	wire horizontal_tile_24_17_to_tile_24_18_1;
	wire horizontal_tile_24_17_to_tile_24_18_2;
	wire horizontal_tile_24_17_to_tile_24_18_3;
	wire horizontal_tile_24_18_to_tile_24_17_0;
	wire horizontal_tile_24_18_to_tile_24_17_1;
	wire horizontal_tile_24_18_to_tile_24_17_2;
	wire horizontal_tile_24_18_to_tile_24_17_3;

	wire horizontal_tile_25_17_to_tile_25_18_0;
	wire horizontal_tile_25_17_to_tile_25_18_1;
	wire horizontal_tile_25_17_to_tile_25_18_2;
	wire horizontal_tile_25_17_to_tile_25_18_3;
	wire horizontal_tile_25_18_to_tile_25_17_0;
	wire horizontal_tile_25_18_to_tile_25_17_1;
	wire horizontal_tile_25_18_to_tile_25_17_2;
	wire horizontal_tile_25_18_to_tile_25_17_3;

	wire horizontal_tile_26_17_to_tile_26_18_0;
	wire horizontal_tile_26_17_to_tile_26_18_1;
	wire horizontal_tile_26_17_to_tile_26_18_2;
	wire horizontal_tile_26_17_to_tile_26_18_3;
	wire horizontal_tile_26_18_to_tile_26_17_0;
	wire horizontal_tile_26_18_to_tile_26_17_1;
	wire horizontal_tile_26_18_to_tile_26_17_2;
	wire horizontal_tile_26_18_to_tile_26_17_3;

	wire horizontal_tile_27_17_to_tile_27_18_0;
	wire horizontal_tile_27_17_to_tile_27_18_1;
	wire horizontal_tile_27_17_to_tile_27_18_2;
	wire horizontal_tile_27_17_to_tile_27_18_3;
	wire horizontal_tile_27_18_to_tile_27_17_0;
	wire horizontal_tile_27_18_to_tile_27_17_1;
	wire horizontal_tile_27_18_to_tile_27_17_2;
	wire horizontal_tile_27_18_to_tile_27_17_3;

	wire horizontal_tile_28_17_to_tile_28_18_0;
	wire horizontal_tile_28_17_to_tile_28_18_1;
	wire horizontal_tile_28_17_to_tile_28_18_2;
	wire horizontal_tile_28_17_to_tile_28_18_3;
	wire horizontal_tile_28_18_to_tile_28_17_0;
	wire horizontal_tile_28_18_to_tile_28_17_1;
	wire horizontal_tile_28_18_to_tile_28_17_2;
	wire horizontal_tile_28_18_to_tile_28_17_3;

	wire horizontal_tile_29_17_to_tile_29_18_0;
	wire horizontal_tile_29_17_to_tile_29_18_1;
	wire horizontal_tile_29_17_to_tile_29_18_2;
	wire horizontal_tile_29_17_to_tile_29_18_3;
	wire horizontal_tile_29_18_to_tile_29_17_0;
	wire horizontal_tile_29_18_to_tile_29_17_1;
	wire horizontal_tile_29_18_to_tile_29_17_2;
	wire horizontal_tile_29_18_to_tile_29_17_3;

	wire horizontal_tile_30_17_to_tile_30_18_0;
	wire horizontal_tile_30_17_to_tile_30_18_1;
	wire horizontal_tile_30_17_to_tile_30_18_2;
	wire horizontal_tile_30_17_to_tile_30_18_3;
	wire horizontal_tile_30_18_to_tile_30_17_0;
	wire horizontal_tile_30_18_to_tile_30_17_1;
	wire horizontal_tile_30_18_to_tile_30_17_2;
	wire horizontal_tile_30_18_to_tile_30_17_3;

	wire horizontal_tile_31_17_to_tile_31_18_0;
	wire horizontal_tile_31_17_to_tile_31_18_1;
	wire horizontal_tile_31_17_to_tile_31_18_2;
	wire horizontal_tile_31_17_to_tile_31_18_3;
	wire horizontal_tile_31_18_to_tile_31_17_0;
	wire horizontal_tile_31_18_to_tile_31_17_1;
	wire horizontal_tile_31_18_to_tile_31_17_2;
	wire horizontal_tile_31_18_to_tile_31_17_3;

	wire horizontal_tile_0_18_to_tile_0_19_0;
	wire horizontal_tile_0_18_to_tile_0_19_1;
	wire horizontal_tile_0_18_to_tile_0_19_2;
	wire horizontal_tile_0_18_to_tile_0_19_3;
	wire horizontal_tile_0_19_to_tile_0_18_0;
	wire horizontal_tile_0_19_to_tile_0_18_1;
	wire horizontal_tile_0_19_to_tile_0_18_2;
	wire horizontal_tile_0_19_to_tile_0_18_3;

	wire horizontal_tile_1_18_to_tile_1_19_0;
	wire horizontal_tile_1_18_to_tile_1_19_1;
	wire horizontal_tile_1_18_to_tile_1_19_2;
	wire horizontal_tile_1_18_to_tile_1_19_3;
	wire horizontal_tile_1_19_to_tile_1_18_0;
	wire horizontal_tile_1_19_to_tile_1_18_1;
	wire horizontal_tile_1_19_to_tile_1_18_2;
	wire horizontal_tile_1_19_to_tile_1_18_3;

	wire horizontal_tile_2_18_to_tile_2_19_0;
	wire horizontal_tile_2_18_to_tile_2_19_1;
	wire horizontal_tile_2_18_to_tile_2_19_2;
	wire horizontal_tile_2_18_to_tile_2_19_3;
	wire horizontal_tile_2_19_to_tile_2_18_0;
	wire horizontal_tile_2_19_to_tile_2_18_1;
	wire horizontal_tile_2_19_to_tile_2_18_2;
	wire horizontal_tile_2_19_to_tile_2_18_3;

	wire horizontal_tile_3_18_to_tile_3_19_0;
	wire horizontal_tile_3_18_to_tile_3_19_1;
	wire horizontal_tile_3_18_to_tile_3_19_2;
	wire horizontal_tile_3_18_to_tile_3_19_3;
	wire horizontal_tile_3_19_to_tile_3_18_0;
	wire horizontal_tile_3_19_to_tile_3_18_1;
	wire horizontal_tile_3_19_to_tile_3_18_2;
	wire horizontal_tile_3_19_to_tile_3_18_3;

	wire horizontal_tile_4_18_to_tile_4_19_0;
	wire horizontal_tile_4_18_to_tile_4_19_1;
	wire horizontal_tile_4_18_to_tile_4_19_2;
	wire horizontal_tile_4_18_to_tile_4_19_3;
	wire horizontal_tile_4_19_to_tile_4_18_0;
	wire horizontal_tile_4_19_to_tile_4_18_1;
	wire horizontal_tile_4_19_to_tile_4_18_2;
	wire horizontal_tile_4_19_to_tile_4_18_3;

	wire horizontal_tile_5_18_to_tile_5_19_0;
	wire horizontal_tile_5_18_to_tile_5_19_1;
	wire horizontal_tile_5_18_to_tile_5_19_2;
	wire horizontal_tile_5_18_to_tile_5_19_3;
	wire horizontal_tile_5_19_to_tile_5_18_0;
	wire horizontal_tile_5_19_to_tile_5_18_1;
	wire horizontal_tile_5_19_to_tile_5_18_2;
	wire horizontal_tile_5_19_to_tile_5_18_3;

	wire horizontal_tile_6_18_to_tile_6_19_0;
	wire horizontal_tile_6_18_to_tile_6_19_1;
	wire horizontal_tile_6_18_to_tile_6_19_2;
	wire horizontal_tile_6_18_to_tile_6_19_3;
	wire horizontal_tile_6_19_to_tile_6_18_0;
	wire horizontal_tile_6_19_to_tile_6_18_1;
	wire horizontal_tile_6_19_to_tile_6_18_2;
	wire horizontal_tile_6_19_to_tile_6_18_3;

	wire horizontal_tile_7_18_to_tile_7_19_0;
	wire horizontal_tile_7_18_to_tile_7_19_1;
	wire horizontal_tile_7_18_to_tile_7_19_2;
	wire horizontal_tile_7_18_to_tile_7_19_3;
	wire horizontal_tile_7_19_to_tile_7_18_0;
	wire horizontal_tile_7_19_to_tile_7_18_1;
	wire horizontal_tile_7_19_to_tile_7_18_2;
	wire horizontal_tile_7_19_to_tile_7_18_3;

	wire horizontal_tile_8_18_to_tile_8_19_0;
	wire horizontal_tile_8_18_to_tile_8_19_1;
	wire horizontal_tile_8_18_to_tile_8_19_2;
	wire horizontal_tile_8_18_to_tile_8_19_3;
	wire horizontal_tile_8_19_to_tile_8_18_0;
	wire horizontal_tile_8_19_to_tile_8_18_1;
	wire horizontal_tile_8_19_to_tile_8_18_2;
	wire horizontal_tile_8_19_to_tile_8_18_3;

	wire horizontal_tile_9_18_to_tile_9_19_0;
	wire horizontal_tile_9_18_to_tile_9_19_1;
	wire horizontal_tile_9_18_to_tile_9_19_2;
	wire horizontal_tile_9_18_to_tile_9_19_3;
	wire horizontal_tile_9_19_to_tile_9_18_0;
	wire horizontal_tile_9_19_to_tile_9_18_1;
	wire horizontal_tile_9_19_to_tile_9_18_2;
	wire horizontal_tile_9_19_to_tile_9_18_3;

	wire horizontal_tile_10_18_to_tile_10_19_0;
	wire horizontal_tile_10_18_to_tile_10_19_1;
	wire horizontal_tile_10_18_to_tile_10_19_2;
	wire horizontal_tile_10_18_to_tile_10_19_3;
	wire horizontal_tile_10_19_to_tile_10_18_0;
	wire horizontal_tile_10_19_to_tile_10_18_1;
	wire horizontal_tile_10_19_to_tile_10_18_2;
	wire horizontal_tile_10_19_to_tile_10_18_3;

	wire horizontal_tile_11_18_to_tile_11_19_0;
	wire horizontal_tile_11_18_to_tile_11_19_1;
	wire horizontal_tile_11_18_to_tile_11_19_2;
	wire horizontal_tile_11_18_to_tile_11_19_3;
	wire horizontal_tile_11_19_to_tile_11_18_0;
	wire horizontal_tile_11_19_to_tile_11_18_1;
	wire horizontal_tile_11_19_to_tile_11_18_2;
	wire horizontal_tile_11_19_to_tile_11_18_3;

	wire horizontal_tile_12_18_to_tile_12_19_0;
	wire horizontal_tile_12_18_to_tile_12_19_1;
	wire horizontal_tile_12_18_to_tile_12_19_2;
	wire horizontal_tile_12_18_to_tile_12_19_3;
	wire horizontal_tile_12_19_to_tile_12_18_0;
	wire horizontal_tile_12_19_to_tile_12_18_1;
	wire horizontal_tile_12_19_to_tile_12_18_2;
	wire horizontal_tile_12_19_to_tile_12_18_3;

	wire horizontal_tile_13_18_to_tile_13_19_0;
	wire horizontal_tile_13_18_to_tile_13_19_1;
	wire horizontal_tile_13_18_to_tile_13_19_2;
	wire horizontal_tile_13_18_to_tile_13_19_3;
	wire horizontal_tile_13_19_to_tile_13_18_0;
	wire horizontal_tile_13_19_to_tile_13_18_1;
	wire horizontal_tile_13_19_to_tile_13_18_2;
	wire horizontal_tile_13_19_to_tile_13_18_3;

	wire horizontal_tile_14_18_to_tile_14_19_0;
	wire horizontal_tile_14_18_to_tile_14_19_1;
	wire horizontal_tile_14_18_to_tile_14_19_2;
	wire horizontal_tile_14_18_to_tile_14_19_3;
	wire horizontal_tile_14_19_to_tile_14_18_0;
	wire horizontal_tile_14_19_to_tile_14_18_1;
	wire horizontal_tile_14_19_to_tile_14_18_2;
	wire horizontal_tile_14_19_to_tile_14_18_3;

	wire horizontal_tile_15_18_to_tile_15_19_0;
	wire horizontal_tile_15_18_to_tile_15_19_1;
	wire horizontal_tile_15_18_to_tile_15_19_2;
	wire horizontal_tile_15_18_to_tile_15_19_3;
	wire horizontal_tile_15_19_to_tile_15_18_0;
	wire horizontal_tile_15_19_to_tile_15_18_1;
	wire horizontal_tile_15_19_to_tile_15_18_2;
	wire horizontal_tile_15_19_to_tile_15_18_3;

	wire horizontal_tile_16_18_to_tile_16_19_0;
	wire horizontal_tile_16_18_to_tile_16_19_1;
	wire horizontal_tile_16_18_to_tile_16_19_2;
	wire horizontal_tile_16_18_to_tile_16_19_3;
	wire horizontal_tile_16_19_to_tile_16_18_0;
	wire horizontal_tile_16_19_to_tile_16_18_1;
	wire horizontal_tile_16_19_to_tile_16_18_2;
	wire horizontal_tile_16_19_to_tile_16_18_3;

	wire horizontal_tile_17_18_to_tile_17_19_0;
	wire horizontal_tile_17_18_to_tile_17_19_1;
	wire horizontal_tile_17_18_to_tile_17_19_2;
	wire horizontal_tile_17_18_to_tile_17_19_3;
	wire horizontal_tile_17_19_to_tile_17_18_0;
	wire horizontal_tile_17_19_to_tile_17_18_1;
	wire horizontal_tile_17_19_to_tile_17_18_2;
	wire horizontal_tile_17_19_to_tile_17_18_3;

	wire horizontal_tile_18_18_to_tile_18_19_0;
	wire horizontal_tile_18_18_to_tile_18_19_1;
	wire horizontal_tile_18_18_to_tile_18_19_2;
	wire horizontal_tile_18_18_to_tile_18_19_3;
	wire horizontal_tile_18_19_to_tile_18_18_0;
	wire horizontal_tile_18_19_to_tile_18_18_1;
	wire horizontal_tile_18_19_to_tile_18_18_2;
	wire horizontal_tile_18_19_to_tile_18_18_3;

	wire horizontal_tile_19_18_to_tile_19_19_0;
	wire horizontal_tile_19_18_to_tile_19_19_1;
	wire horizontal_tile_19_18_to_tile_19_19_2;
	wire horizontal_tile_19_18_to_tile_19_19_3;
	wire horizontal_tile_19_19_to_tile_19_18_0;
	wire horizontal_tile_19_19_to_tile_19_18_1;
	wire horizontal_tile_19_19_to_tile_19_18_2;
	wire horizontal_tile_19_19_to_tile_19_18_3;

	wire horizontal_tile_20_18_to_tile_20_19_0;
	wire horizontal_tile_20_18_to_tile_20_19_1;
	wire horizontal_tile_20_18_to_tile_20_19_2;
	wire horizontal_tile_20_18_to_tile_20_19_3;
	wire horizontal_tile_20_19_to_tile_20_18_0;
	wire horizontal_tile_20_19_to_tile_20_18_1;
	wire horizontal_tile_20_19_to_tile_20_18_2;
	wire horizontal_tile_20_19_to_tile_20_18_3;

	wire horizontal_tile_21_18_to_tile_21_19_0;
	wire horizontal_tile_21_18_to_tile_21_19_1;
	wire horizontal_tile_21_18_to_tile_21_19_2;
	wire horizontal_tile_21_18_to_tile_21_19_3;
	wire horizontal_tile_21_19_to_tile_21_18_0;
	wire horizontal_tile_21_19_to_tile_21_18_1;
	wire horizontal_tile_21_19_to_tile_21_18_2;
	wire horizontal_tile_21_19_to_tile_21_18_3;

	wire horizontal_tile_22_18_to_tile_22_19_0;
	wire horizontal_tile_22_18_to_tile_22_19_1;
	wire horizontal_tile_22_18_to_tile_22_19_2;
	wire horizontal_tile_22_18_to_tile_22_19_3;
	wire horizontal_tile_22_19_to_tile_22_18_0;
	wire horizontal_tile_22_19_to_tile_22_18_1;
	wire horizontal_tile_22_19_to_tile_22_18_2;
	wire horizontal_tile_22_19_to_tile_22_18_3;

	wire horizontal_tile_23_18_to_tile_23_19_0;
	wire horizontal_tile_23_18_to_tile_23_19_1;
	wire horizontal_tile_23_18_to_tile_23_19_2;
	wire horizontal_tile_23_18_to_tile_23_19_3;
	wire horizontal_tile_23_19_to_tile_23_18_0;
	wire horizontal_tile_23_19_to_tile_23_18_1;
	wire horizontal_tile_23_19_to_tile_23_18_2;
	wire horizontal_tile_23_19_to_tile_23_18_3;

	wire horizontal_tile_24_18_to_tile_24_19_0;
	wire horizontal_tile_24_18_to_tile_24_19_1;
	wire horizontal_tile_24_18_to_tile_24_19_2;
	wire horizontal_tile_24_18_to_tile_24_19_3;
	wire horizontal_tile_24_19_to_tile_24_18_0;
	wire horizontal_tile_24_19_to_tile_24_18_1;
	wire horizontal_tile_24_19_to_tile_24_18_2;
	wire horizontal_tile_24_19_to_tile_24_18_3;

	wire horizontal_tile_25_18_to_tile_25_19_0;
	wire horizontal_tile_25_18_to_tile_25_19_1;
	wire horizontal_tile_25_18_to_tile_25_19_2;
	wire horizontal_tile_25_18_to_tile_25_19_3;
	wire horizontal_tile_25_19_to_tile_25_18_0;
	wire horizontal_tile_25_19_to_tile_25_18_1;
	wire horizontal_tile_25_19_to_tile_25_18_2;
	wire horizontal_tile_25_19_to_tile_25_18_3;

	wire horizontal_tile_26_18_to_tile_26_19_0;
	wire horizontal_tile_26_18_to_tile_26_19_1;
	wire horizontal_tile_26_18_to_tile_26_19_2;
	wire horizontal_tile_26_18_to_tile_26_19_3;
	wire horizontal_tile_26_19_to_tile_26_18_0;
	wire horizontal_tile_26_19_to_tile_26_18_1;
	wire horizontal_tile_26_19_to_tile_26_18_2;
	wire horizontal_tile_26_19_to_tile_26_18_3;

	wire horizontal_tile_27_18_to_tile_27_19_0;
	wire horizontal_tile_27_18_to_tile_27_19_1;
	wire horizontal_tile_27_18_to_tile_27_19_2;
	wire horizontal_tile_27_18_to_tile_27_19_3;
	wire horizontal_tile_27_19_to_tile_27_18_0;
	wire horizontal_tile_27_19_to_tile_27_18_1;
	wire horizontal_tile_27_19_to_tile_27_18_2;
	wire horizontal_tile_27_19_to_tile_27_18_3;

	wire horizontal_tile_28_18_to_tile_28_19_0;
	wire horizontal_tile_28_18_to_tile_28_19_1;
	wire horizontal_tile_28_18_to_tile_28_19_2;
	wire horizontal_tile_28_18_to_tile_28_19_3;
	wire horizontal_tile_28_19_to_tile_28_18_0;
	wire horizontal_tile_28_19_to_tile_28_18_1;
	wire horizontal_tile_28_19_to_tile_28_18_2;
	wire horizontal_tile_28_19_to_tile_28_18_3;

	wire horizontal_tile_29_18_to_tile_29_19_0;
	wire horizontal_tile_29_18_to_tile_29_19_1;
	wire horizontal_tile_29_18_to_tile_29_19_2;
	wire horizontal_tile_29_18_to_tile_29_19_3;
	wire horizontal_tile_29_19_to_tile_29_18_0;
	wire horizontal_tile_29_19_to_tile_29_18_1;
	wire horizontal_tile_29_19_to_tile_29_18_2;
	wire horizontal_tile_29_19_to_tile_29_18_3;

	wire horizontal_tile_30_18_to_tile_30_19_0;
	wire horizontal_tile_30_18_to_tile_30_19_1;
	wire horizontal_tile_30_18_to_tile_30_19_2;
	wire horizontal_tile_30_18_to_tile_30_19_3;
	wire horizontal_tile_30_19_to_tile_30_18_0;
	wire horizontal_tile_30_19_to_tile_30_18_1;
	wire horizontal_tile_30_19_to_tile_30_18_2;
	wire horizontal_tile_30_19_to_tile_30_18_3;

	wire horizontal_tile_31_18_to_tile_31_19_0;
	wire horizontal_tile_31_18_to_tile_31_19_1;
	wire horizontal_tile_31_18_to_tile_31_19_2;
	wire horizontal_tile_31_18_to_tile_31_19_3;
	wire horizontal_tile_31_19_to_tile_31_18_0;
	wire horizontal_tile_31_19_to_tile_31_18_1;
	wire horizontal_tile_31_19_to_tile_31_18_2;
	wire horizontal_tile_31_19_to_tile_31_18_3;

	wire horizontal_tile_0_19_to_tile_0_20_0;
	wire horizontal_tile_0_19_to_tile_0_20_1;
	wire horizontal_tile_0_19_to_tile_0_20_2;
	wire horizontal_tile_0_19_to_tile_0_20_3;
	wire horizontal_tile_0_20_to_tile_0_19_0;
	wire horizontal_tile_0_20_to_tile_0_19_1;
	wire horizontal_tile_0_20_to_tile_0_19_2;
	wire horizontal_tile_0_20_to_tile_0_19_3;

	wire horizontal_tile_1_19_to_tile_1_20_0;
	wire horizontal_tile_1_19_to_tile_1_20_1;
	wire horizontal_tile_1_19_to_tile_1_20_2;
	wire horizontal_tile_1_19_to_tile_1_20_3;
	wire horizontal_tile_1_20_to_tile_1_19_0;
	wire horizontal_tile_1_20_to_tile_1_19_1;
	wire horizontal_tile_1_20_to_tile_1_19_2;
	wire horizontal_tile_1_20_to_tile_1_19_3;

	wire horizontal_tile_2_19_to_tile_2_20_0;
	wire horizontal_tile_2_19_to_tile_2_20_1;
	wire horizontal_tile_2_19_to_tile_2_20_2;
	wire horizontal_tile_2_19_to_tile_2_20_3;
	wire horizontal_tile_2_20_to_tile_2_19_0;
	wire horizontal_tile_2_20_to_tile_2_19_1;
	wire horizontal_tile_2_20_to_tile_2_19_2;
	wire horizontal_tile_2_20_to_tile_2_19_3;

	wire horizontal_tile_3_19_to_tile_3_20_0;
	wire horizontal_tile_3_19_to_tile_3_20_1;
	wire horizontal_tile_3_19_to_tile_3_20_2;
	wire horizontal_tile_3_19_to_tile_3_20_3;
	wire horizontal_tile_3_20_to_tile_3_19_0;
	wire horizontal_tile_3_20_to_tile_3_19_1;
	wire horizontal_tile_3_20_to_tile_3_19_2;
	wire horizontal_tile_3_20_to_tile_3_19_3;

	wire horizontal_tile_4_19_to_tile_4_20_0;
	wire horizontal_tile_4_19_to_tile_4_20_1;
	wire horizontal_tile_4_19_to_tile_4_20_2;
	wire horizontal_tile_4_19_to_tile_4_20_3;
	wire horizontal_tile_4_20_to_tile_4_19_0;
	wire horizontal_tile_4_20_to_tile_4_19_1;
	wire horizontal_tile_4_20_to_tile_4_19_2;
	wire horizontal_tile_4_20_to_tile_4_19_3;

	wire horizontal_tile_5_19_to_tile_5_20_0;
	wire horizontal_tile_5_19_to_tile_5_20_1;
	wire horizontal_tile_5_19_to_tile_5_20_2;
	wire horizontal_tile_5_19_to_tile_5_20_3;
	wire horizontal_tile_5_20_to_tile_5_19_0;
	wire horizontal_tile_5_20_to_tile_5_19_1;
	wire horizontal_tile_5_20_to_tile_5_19_2;
	wire horizontal_tile_5_20_to_tile_5_19_3;

	wire horizontal_tile_6_19_to_tile_6_20_0;
	wire horizontal_tile_6_19_to_tile_6_20_1;
	wire horizontal_tile_6_19_to_tile_6_20_2;
	wire horizontal_tile_6_19_to_tile_6_20_3;
	wire horizontal_tile_6_20_to_tile_6_19_0;
	wire horizontal_tile_6_20_to_tile_6_19_1;
	wire horizontal_tile_6_20_to_tile_6_19_2;
	wire horizontal_tile_6_20_to_tile_6_19_3;

	wire horizontal_tile_7_19_to_tile_7_20_0;
	wire horizontal_tile_7_19_to_tile_7_20_1;
	wire horizontal_tile_7_19_to_tile_7_20_2;
	wire horizontal_tile_7_19_to_tile_7_20_3;
	wire horizontal_tile_7_20_to_tile_7_19_0;
	wire horizontal_tile_7_20_to_tile_7_19_1;
	wire horizontal_tile_7_20_to_tile_7_19_2;
	wire horizontal_tile_7_20_to_tile_7_19_3;

	wire horizontal_tile_8_19_to_tile_8_20_0;
	wire horizontal_tile_8_19_to_tile_8_20_1;
	wire horizontal_tile_8_19_to_tile_8_20_2;
	wire horizontal_tile_8_19_to_tile_8_20_3;
	wire horizontal_tile_8_20_to_tile_8_19_0;
	wire horizontal_tile_8_20_to_tile_8_19_1;
	wire horizontal_tile_8_20_to_tile_8_19_2;
	wire horizontal_tile_8_20_to_tile_8_19_3;

	wire horizontal_tile_9_19_to_tile_9_20_0;
	wire horizontal_tile_9_19_to_tile_9_20_1;
	wire horizontal_tile_9_19_to_tile_9_20_2;
	wire horizontal_tile_9_19_to_tile_9_20_3;
	wire horizontal_tile_9_20_to_tile_9_19_0;
	wire horizontal_tile_9_20_to_tile_9_19_1;
	wire horizontal_tile_9_20_to_tile_9_19_2;
	wire horizontal_tile_9_20_to_tile_9_19_3;

	wire horizontal_tile_10_19_to_tile_10_20_0;
	wire horizontal_tile_10_19_to_tile_10_20_1;
	wire horizontal_tile_10_19_to_tile_10_20_2;
	wire horizontal_tile_10_19_to_tile_10_20_3;
	wire horizontal_tile_10_20_to_tile_10_19_0;
	wire horizontal_tile_10_20_to_tile_10_19_1;
	wire horizontal_tile_10_20_to_tile_10_19_2;
	wire horizontal_tile_10_20_to_tile_10_19_3;

	wire horizontal_tile_11_19_to_tile_11_20_0;
	wire horizontal_tile_11_19_to_tile_11_20_1;
	wire horizontal_tile_11_19_to_tile_11_20_2;
	wire horizontal_tile_11_19_to_tile_11_20_3;
	wire horizontal_tile_11_20_to_tile_11_19_0;
	wire horizontal_tile_11_20_to_tile_11_19_1;
	wire horizontal_tile_11_20_to_tile_11_19_2;
	wire horizontal_tile_11_20_to_tile_11_19_3;

	wire horizontal_tile_12_19_to_tile_12_20_0;
	wire horizontal_tile_12_19_to_tile_12_20_1;
	wire horizontal_tile_12_19_to_tile_12_20_2;
	wire horizontal_tile_12_19_to_tile_12_20_3;
	wire horizontal_tile_12_20_to_tile_12_19_0;
	wire horizontal_tile_12_20_to_tile_12_19_1;
	wire horizontal_tile_12_20_to_tile_12_19_2;
	wire horizontal_tile_12_20_to_tile_12_19_3;

	wire horizontal_tile_13_19_to_tile_13_20_0;
	wire horizontal_tile_13_19_to_tile_13_20_1;
	wire horizontal_tile_13_19_to_tile_13_20_2;
	wire horizontal_tile_13_19_to_tile_13_20_3;
	wire horizontal_tile_13_20_to_tile_13_19_0;
	wire horizontal_tile_13_20_to_tile_13_19_1;
	wire horizontal_tile_13_20_to_tile_13_19_2;
	wire horizontal_tile_13_20_to_tile_13_19_3;

	wire horizontal_tile_14_19_to_tile_14_20_0;
	wire horizontal_tile_14_19_to_tile_14_20_1;
	wire horizontal_tile_14_19_to_tile_14_20_2;
	wire horizontal_tile_14_19_to_tile_14_20_3;
	wire horizontal_tile_14_20_to_tile_14_19_0;
	wire horizontal_tile_14_20_to_tile_14_19_1;
	wire horizontal_tile_14_20_to_tile_14_19_2;
	wire horizontal_tile_14_20_to_tile_14_19_3;

	wire horizontal_tile_15_19_to_tile_15_20_0;
	wire horizontal_tile_15_19_to_tile_15_20_1;
	wire horizontal_tile_15_19_to_tile_15_20_2;
	wire horizontal_tile_15_19_to_tile_15_20_3;
	wire horizontal_tile_15_20_to_tile_15_19_0;
	wire horizontal_tile_15_20_to_tile_15_19_1;
	wire horizontal_tile_15_20_to_tile_15_19_2;
	wire horizontal_tile_15_20_to_tile_15_19_3;

	wire horizontal_tile_16_19_to_tile_16_20_0;
	wire horizontal_tile_16_19_to_tile_16_20_1;
	wire horizontal_tile_16_19_to_tile_16_20_2;
	wire horizontal_tile_16_19_to_tile_16_20_3;
	wire horizontal_tile_16_20_to_tile_16_19_0;
	wire horizontal_tile_16_20_to_tile_16_19_1;
	wire horizontal_tile_16_20_to_tile_16_19_2;
	wire horizontal_tile_16_20_to_tile_16_19_3;

	wire horizontal_tile_17_19_to_tile_17_20_0;
	wire horizontal_tile_17_19_to_tile_17_20_1;
	wire horizontal_tile_17_19_to_tile_17_20_2;
	wire horizontal_tile_17_19_to_tile_17_20_3;
	wire horizontal_tile_17_20_to_tile_17_19_0;
	wire horizontal_tile_17_20_to_tile_17_19_1;
	wire horizontal_tile_17_20_to_tile_17_19_2;
	wire horizontal_tile_17_20_to_tile_17_19_3;

	wire horizontal_tile_18_19_to_tile_18_20_0;
	wire horizontal_tile_18_19_to_tile_18_20_1;
	wire horizontal_tile_18_19_to_tile_18_20_2;
	wire horizontal_tile_18_19_to_tile_18_20_3;
	wire horizontal_tile_18_20_to_tile_18_19_0;
	wire horizontal_tile_18_20_to_tile_18_19_1;
	wire horizontal_tile_18_20_to_tile_18_19_2;
	wire horizontal_tile_18_20_to_tile_18_19_3;

	wire horizontal_tile_19_19_to_tile_19_20_0;
	wire horizontal_tile_19_19_to_tile_19_20_1;
	wire horizontal_tile_19_19_to_tile_19_20_2;
	wire horizontal_tile_19_19_to_tile_19_20_3;
	wire horizontal_tile_19_20_to_tile_19_19_0;
	wire horizontal_tile_19_20_to_tile_19_19_1;
	wire horizontal_tile_19_20_to_tile_19_19_2;
	wire horizontal_tile_19_20_to_tile_19_19_3;

	wire horizontal_tile_20_19_to_tile_20_20_0;
	wire horizontal_tile_20_19_to_tile_20_20_1;
	wire horizontal_tile_20_19_to_tile_20_20_2;
	wire horizontal_tile_20_19_to_tile_20_20_3;
	wire horizontal_tile_20_20_to_tile_20_19_0;
	wire horizontal_tile_20_20_to_tile_20_19_1;
	wire horizontal_tile_20_20_to_tile_20_19_2;
	wire horizontal_tile_20_20_to_tile_20_19_3;

	wire horizontal_tile_21_19_to_tile_21_20_0;
	wire horizontal_tile_21_19_to_tile_21_20_1;
	wire horizontal_tile_21_19_to_tile_21_20_2;
	wire horizontal_tile_21_19_to_tile_21_20_3;
	wire horizontal_tile_21_20_to_tile_21_19_0;
	wire horizontal_tile_21_20_to_tile_21_19_1;
	wire horizontal_tile_21_20_to_tile_21_19_2;
	wire horizontal_tile_21_20_to_tile_21_19_3;

	wire horizontal_tile_22_19_to_tile_22_20_0;
	wire horizontal_tile_22_19_to_tile_22_20_1;
	wire horizontal_tile_22_19_to_tile_22_20_2;
	wire horizontal_tile_22_19_to_tile_22_20_3;
	wire horizontal_tile_22_20_to_tile_22_19_0;
	wire horizontal_tile_22_20_to_tile_22_19_1;
	wire horizontal_tile_22_20_to_tile_22_19_2;
	wire horizontal_tile_22_20_to_tile_22_19_3;

	wire horizontal_tile_23_19_to_tile_23_20_0;
	wire horizontal_tile_23_19_to_tile_23_20_1;
	wire horizontal_tile_23_19_to_tile_23_20_2;
	wire horizontal_tile_23_19_to_tile_23_20_3;
	wire horizontal_tile_23_20_to_tile_23_19_0;
	wire horizontal_tile_23_20_to_tile_23_19_1;
	wire horizontal_tile_23_20_to_tile_23_19_2;
	wire horizontal_tile_23_20_to_tile_23_19_3;

	wire horizontal_tile_24_19_to_tile_24_20_0;
	wire horizontal_tile_24_19_to_tile_24_20_1;
	wire horizontal_tile_24_19_to_tile_24_20_2;
	wire horizontal_tile_24_19_to_tile_24_20_3;
	wire horizontal_tile_24_20_to_tile_24_19_0;
	wire horizontal_tile_24_20_to_tile_24_19_1;
	wire horizontal_tile_24_20_to_tile_24_19_2;
	wire horizontal_tile_24_20_to_tile_24_19_3;

	wire horizontal_tile_25_19_to_tile_25_20_0;
	wire horizontal_tile_25_19_to_tile_25_20_1;
	wire horizontal_tile_25_19_to_tile_25_20_2;
	wire horizontal_tile_25_19_to_tile_25_20_3;
	wire horizontal_tile_25_20_to_tile_25_19_0;
	wire horizontal_tile_25_20_to_tile_25_19_1;
	wire horizontal_tile_25_20_to_tile_25_19_2;
	wire horizontal_tile_25_20_to_tile_25_19_3;

	wire horizontal_tile_26_19_to_tile_26_20_0;
	wire horizontal_tile_26_19_to_tile_26_20_1;
	wire horizontal_tile_26_19_to_tile_26_20_2;
	wire horizontal_tile_26_19_to_tile_26_20_3;
	wire horizontal_tile_26_20_to_tile_26_19_0;
	wire horizontal_tile_26_20_to_tile_26_19_1;
	wire horizontal_tile_26_20_to_tile_26_19_2;
	wire horizontal_tile_26_20_to_tile_26_19_3;

	wire horizontal_tile_27_19_to_tile_27_20_0;
	wire horizontal_tile_27_19_to_tile_27_20_1;
	wire horizontal_tile_27_19_to_tile_27_20_2;
	wire horizontal_tile_27_19_to_tile_27_20_3;
	wire horizontal_tile_27_20_to_tile_27_19_0;
	wire horizontal_tile_27_20_to_tile_27_19_1;
	wire horizontal_tile_27_20_to_tile_27_19_2;
	wire horizontal_tile_27_20_to_tile_27_19_3;

	wire horizontal_tile_28_19_to_tile_28_20_0;
	wire horizontal_tile_28_19_to_tile_28_20_1;
	wire horizontal_tile_28_19_to_tile_28_20_2;
	wire horizontal_tile_28_19_to_tile_28_20_3;
	wire horizontal_tile_28_20_to_tile_28_19_0;
	wire horizontal_tile_28_20_to_tile_28_19_1;
	wire horizontal_tile_28_20_to_tile_28_19_2;
	wire horizontal_tile_28_20_to_tile_28_19_3;

	wire horizontal_tile_29_19_to_tile_29_20_0;
	wire horizontal_tile_29_19_to_tile_29_20_1;
	wire horizontal_tile_29_19_to_tile_29_20_2;
	wire horizontal_tile_29_19_to_tile_29_20_3;
	wire horizontal_tile_29_20_to_tile_29_19_0;
	wire horizontal_tile_29_20_to_tile_29_19_1;
	wire horizontal_tile_29_20_to_tile_29_19_2;
	wire horizontal_tile_29_20_to_tile_29_19_3;

	wire horizontal_tile_30_19_to_tile_30_20_0;
	wire horizontal_tile_30_19_to_tile_30_20_1;
	wire horizontal_tile_30_19_to_tile_30_20_2;
	wire horizontal_tile_30_19_to_tile_30_20_3;
	wire horizontal_tile_30_20_to_tile_30_19_0;
	wire horizontal_tile_30_20_to_tile_30_19_1;
	wire horizontal_tile_30_20_to_tile_30_19_2;
	wire horizontal_tile_30_20_to_tile_30_19_3;

	wire horizontal_tile_31_19_to_tile_31_20_0;
	wire horizontal_tile_31_19_to_tile_31_20_1;
	wire horizontal_tile_31_19_to_tile_31_20_2;
	wire horizontal_tile_31_19_to_tile_31_20_3;
	wire horizontal_tile_31_20_to_tile_31_19_0;
	wire horizontal_tile_31_20_to_tile_31_19_1;
	wire horizontal_tile_31_20_to_tile_31_19_2;
	wire horizontal_tile_31_20_to_tile_31_19_3;

	wire horizontal_tile_0_20_to_tile_0_21_0;
	wire horizontal_tile_0_20_to_tile_0_21_1;
	wire horizontal_tile_0_20_to_tile_0_21_2;
	wire horizontal_tile_0_20_to_tile_0_21_3;
	wire horizontal_tile_0_21_to_tile_0_20_0;
	wire horizontal_tile_0_21_to_tile_0_20_1;
	wire horizontal_tile_0_21_to_tile_0_20_2;
	wire horizontal_tile_0_21_to_tile_0_20_3;

	wire horizontal_tile_1_20_to_tile_1_21_0;
	wire horizontal_tile_1_20_to_tile_1_21_1;
	wire horizontal_tile_1_20_to_tile_1_21_2;
	wire horizontal_tile_1_20_to_tile_1_21_3;
	wire horizontal_tile_1_21_to_tile_1_20_0;
	wire horizontal_tile_1_21_to_tile_1_20_1;
	wire horizontal_tile_1_21_to_tile_1_20_2;
	wire horizontal_tile_1_21_to_tile_1_20_3;

	wire horizontal_tile_2_20_to_tile_2_21_0;
	wire horizontal_tile_2_20_to_tile_2_21_1;
	wire horizontal_tile_2_20_to_tile_2_21_2;
	wire horizontal_tile_2_20_to_tile_2_21_3;
	wire horizontal_tile_2_21_to_tile_2_20_0;
	wire horizontal_tile_2_21_to_tile_2_20_1;
	wire horizontal_tile_2_21_to_tile_2_20_2;
	wire horizontal_tile_2_21_to_tile_2_20_3;

	wire horizontal_tile_3_20_to_tile_3_21_0;
	wire horizontal_tile_3_20_to_tile_3_21_1;
	wire horizontal_tile_3_20_to_tile_3_21_2;
	wire horizontal_tile_3_20_to_tile_3_21_3;
	wire horizontal_tile_3_21_to_tile_3_20_0;
	wire horizontal_tile_3_21_to_tile_3_20_1;
	wire horizontal_tile_3_21_to_tile_3_20_2;
	wire horizontal_tile_3_21_to_tile_3_20_3;

	wire horizontal_tile_4_20_to_tile_4_21_0;
	wire horizontal_tile_4_20_to_tile_4_21_1;
	wire horizontal_tile_4_20_to_tile_4_21_2;
	wire horizontal_tile_4_20_to_tile_4_21_3;
	wire horizontal_tile_4_21_to_tile_4_20_0;
	wire horizontal_tile_4_21_to_tile_4_20_1;
	wire horizontal_tile_4_21_to_tile_4_20_2;
	wire horizontal_tile_4_21_to_tile_4_20_3;

	wire horizontal_tile_5_20_to_tile_5_21_0;
	wire horizontal_tile_5_20_to_tile_5_21_1;
	wire horizontal_tile_5_20_to_tile_5_21_2;
	wire horizontal_tile_5_20_to_tile_5_21_3;
	wire horizontal_tile_5_21_to_tile_5_20_0;
	wire horizontal_tile_5_21_to_tile_5_20_1;
	wire horizontal_tile_5_21_to_tile_5_20_2;
	wire horizontal_tile_5_21_to_tile_5_20_3;

	wire horizontal_tile_6_20_to_tile_6_21_0;
	wire horizontal_tile_6_20_to_tile_6_21_1;
	wire horizontal_tile_6_20_to_tile_6_21_2;
	wire horizontal_tile_6_20_to_tile_6_21_3;
	wire horizontal_tile_6_21_to_tile_6_20_0;
	wire horizontal_tile_6_21_to_tile_6_20_1;
	wire horizontal_tile_6_21_to_tile_6_20_2;
	wire horizontal_tile_6_21_to_tile_6_20_3;

	wire horizontal_tile_7_20_to_tile_7_21_0;
	wire horizontal_tile_7_20_to_tile_7_21_1;
	wire horizontal_tile_7_20_to_tile_7_21_2;
	wire horizontal_tile_7_20_to_tile_7_21_3;
	wire horizontal_tile_7_21_to_tile_7_20_0;
	wire horizontal_tile_7_21_to_tile_7_20_1;
	wire horizontal_tile_7_21_to_tile_7_20_2;
	wire horizontal_tile_7_21_to_tile_7_20_3;

	wire horizontal_tile_8_20_to_tile_8_21_0;
	wire horizontal_tile_8_20_to_tile_8_21_1;
	wire horizontal_tile_8_20_to_tile_8_21_2;
	wire horizontal_tile_8_20_to_tile_8_21_3;
	wire horizontal_tile_8_21_to_tile_8_20_0;
	wire horizontal_tile_8_21_to_tile_8_20_1;
	wire horizontal_tile_8_21_to_tile_8_20_2;
	wire horizontal_tile_8_21_to_tile_8_20_3;

	wire horizontal_tile_9_20_to_tile_9_21_0;
	wire horizontal_tile_9_20_to_tile_9_21_1;
	wire horizontal_tile_9_20_to_tile_9_21_2;
	wire horizontal_tile_9_20_to_tile_9_21_3;
	wire horizontal_tile_9_21_to_tile_9_20_0;
	wire horizontal_tile_9_21_to_tile_9_20_1;
	wire horizontal_tile_9_21_to_tile_9_20_2;
	wire horizontal_tile_9_21_to_tile_9_20_3;

	wire horizontal_tile_10_20_to_tile_10_21_0;
	wire horizontal_tile_10_20_to_tile_10_21_1;
	wire horizontal_tile_10_20_to_tile_10_21_2;
	wire horizontal_tile_10_20_to_tile_10_21_3;
	wire horizontal_tile_10_21_to_tile_10_20_0;
	wire horizontal_tile_10_21_to_tile_10_20_1;
	wire horizontal_tile_10_21_to_tile_10_20_2;
	wire horizontal_tile_10_21_to_tile_10_20_3;

	wire horizontal_tile_11_20_to_tile_11_21_0;
	wire horizontal_tile_11_20_to_tile_11_21_1;
	wire horizontal_tile_11_20_to_tile_11_21_2;
	wire horizontal_tile_11_20_to_tile_11_21_3;
	wire horizontal_tile_11_21_to_tile_11_20_0;
	wire horizontal_tile_11_21_to_tile_11_20_1;
	wire horizontal_tile_11_21_to_tile_11_20_2;
	wire horizontal_tile_11_21_to_tile_11_20_3;

	wire horizontal_tile_12_20_to_tile_12_21_0;
	wire horizontal_tile_12_20_to_tile_12_21_1;
	wire horizontal_tile_12_20_to_tile_12_21_2;
	wire horizontal_tile_12_20_to_tile_12_21_3;
	wire horizontal_tile_12_21_to_tile_12_20_0;
	wire horizontal_tile_12_21_to_tile_12_20_1;
	wire horizontal_tile_12_21_to_tile_12_20_2;
	wire horizontal_tile_12_21_to_tile_12_20_3;

	wire horizontal_tile_13_20_to_tile_13_21_0;
	wire horizontal_tile_13_20_to_tile_13_21_1;
	wire horizontal_tile_13_20_to_tile_13_21_2;
	wire horizontal_tile_13_20_to_tile_13_21_3;
	wire horizontal_tile_13_21_to_tile_13_20_0;
	wire horizontal_tile_13_21_to_tile_13_20_1;
	wire horizontal_tile_13_21_to_tile_13_20_2;
	wire horizontal_tile_13_21_to_tile_13_20_3;

	wire horizontal_tile_14_20_to_tile_14_21_0;
	wire horizontal_tile_14_20_to_tile_14_21_1;
	wire horizontal_tile_14_20_to_tile_14_21_2;
	wire horizontal_tile_14_20_to_tile_14_21_3;
	wire horizontal_tile_14_21_to_tile_14_20_0;
	wire horizontal_tile_14_21_to_tile_14_20_1;
	wire horizontal_tile_14_21_to_tile_14_20_2;
	wire horizontal_tile_14_21_to_tile_14_20_3;

	wire horizontal_tile_15_20_to_tile_15_21_0;
	wire horizontal_tile_15_20_to_tile_15_21_1;
	wire horizontal_tile_15_20_to_tile_15_21_2;
	wire horizontal_tile_15_20_to_tile_15_21_3;
	wire horizontal_tile_15_21_to_tile_15_20_0;
	wire horizontal_tile_15_21_to_tile_15_20_1;
	wire horizontal_tile_15_21_to_tile_15_20_2;
	wire horizontal_tile_15_21_to_tile_15_20_3;

	wire horizontal_tile_16_20_to_tile_16_21_0;
	wire horizontal_tile_16_20_to_tile_16_21_1;
	wire horizontal_tile_16_20_to_tile_16_21_2;
	wire horizontal_tile_16_20_to_tile_16_21_3;
	wire horizontal_tile_16_21_to_tile_16_20_0;
	wire horizontal_tile_16_21_to_tile_16_20_1;
	wire horizontal_tile_16_21_to_tile_16_20_2;
	wire horizontal_tile_16_21_to_tile_16_20_3;

	wire horizontal_tile_17_20_to_tile_17_21_0;
	wire horizontal_tile_17_20_to_tile_17_21_1;
	wire horizontal_tile_17_20_to_tile_17_21_2;
	wire horizontal_tile_17_20_to_tile_17_21_3;
	wire horizontal_tile_17_21_to_tile_17_20_0;
	wire horizontal_tile_17_21_to_tile_17_20_1;
	wire horizontal_tile_17_21_to_tile_17_20_2;
	wire horizontal_tile_17_21_to_tile_17_20_3;

	wire horizontal_tile_18_20_to_tile_18_21_0;
	wire horizontal_tile_18_20_to_tile_18_21_1;
	wire horizontal_tile_18_20_to_tile_18_21_2;
	wire horizontal_tile_18_20_to_tile_18_21_3;
	wire horizontal_tile_18_21_to_tile_18_20_0;
	wire horizontal_tile_18_21_to_tile_18_20_1;
	wire horizontal_tile_18_21_to_tile_18_20_2;
	wire horizontal_tile_18_21_to_tile_18_20_3;

	wire horizontal_tile_19_20_to_tile_19_21_0;
	wire horizontal_tile_19_20_to_tile_19_21_1;
	wire horizontal_tile_19_20_to_tile_19_21_2;
	wire horizontal_tile_19_20_to_tile_19_21_3;
	wire horizontal_tile_19_21_to_tile_19_20_0;
	wire horizontal_tile_19_21_to_tile_19_20_1;
	wire horizontal_tile_19_21_to_tile_19_20_2;
	wire horizontal_tile_19_21_to_tile_19_20_3;

	wire horizontal_tile_20_20_to_tile_20_21_0;
	wire horizontal_tile_20_20_to_tile_20_21_1;
	wire horizontal_tile_20_20_to_tile_20_21_2;
	wire horizontal_tile_20_20_to_tile_20_21_3;
	wire horizontal_tile_20_21_to_tile_20_20_0;
	wire horizontal_tile_20_21_to_tile_20_20_1;
	wire horizontal_tile_20_21_to_tile_20_20_2;
	wire horizontal_tile_20_21_to_tile_20_20_3;

	wire horizontal_tile_21_20_to_tile_21_21_0;
	wire horizontal_tile_21_20_to_tile_21_21_1;
	wire horizontal_tile_21_20_to_tile_21_21_2;
	wire horizontal_tile_21_20_to_tile_21_21_3;
	wire horizontal_tile_21_21_to_tile_21_20_0;
	wire horizontal_tile_21_21_to_tile_21_20_1;
	wire horizontal_tile_21_21_to_tile_21_20_2;
	wire horizontal_tile_21_21_to_tile_21_20_3;

	wire horizontal_tile_22_20_to_tile_22_21_0;
	wire horizontal_tile_22_20_to_tile_22_21_1;
	wire horizontal_tile_22_20_to_tile_22_21_2;
	wire horizontal_tile_22_20_to_tile_22_21_3;
	wire horizontal_tile_22_21_to_tile_22_20_0;
	wire horizontal_tile_22_21_to_tile_22_20_1;
	wire horizontal_tile_22_21_to_tile_22_20_2;
	wire horizontal_tile_22_21_to_tile_22_20_3;

	wire horizontal_tile_23_20_to_tile_23_21_0;
	wire horizontal_tile_23_20_to_tile_23_21_1;
	wire horizontal_tile_23_20_to_tile_23_21_2;
	wire horizontal_tile_23_20_to_tile_23_21_3;
	wire horizontal_tile_23_21_to_tile_23_20_0;
	wire horizontal_tile_23_21_to_tile_23_20_1;
	wire horizontal_tile_23_21_to_tile_23_20_2;
	wire horizontal_tile_23_21_to_tile_23_20_3;

	wire horizontal_tile_24_20_to_tile_24_21_0;
	wire horizontal_tile_24_20_to_tile_24_21_1;
	wire horizontal_tile_24_20_to_tile_24_21_2;
	wire horizontal_tile_24_20_to_tile_24_21_3;
	wire horizontal_tile_24_21_to_tile_24_20_0;
	wire horizontal_tile_24_21_to_tile_24_20_1;
	wire horizontal_tile_24_21_to_tile_24_20_2;
	wire horizontal_tile_24_21_to_tile_24_20_3;

	wire horizontal_tile_25_20_to_tile_25_21_0;
	wire horizontal_tile_25_20_to_tile_25_21_1;
	wire horizontal_tile_25_20_to_tile_25_21_2;
	wire horizontal_tile_25_20_to_tile_25_21_3;
	wire horizontal_tile_25_21_to_tile_25_20_0;
	wire horizontal_tile_25_21_to_tile_25_20_1;
	wire horizontal_tile_25_21_to_tile_25_20_2;
	wire horizontal_tile_25_21_to_tile_25_20_3;

	wire horizontal_tile_26_20_to_tile_26_21_0;
	wire horizontal_tile_26_20_to_tile_26_21_1;
	wire horizontal_tile_26_20_to_tile_26_21_2;
	wire horizontal_tile_26_20_to_tile_26_21_3;
	wire horizontal_tile_26_21_to_tile_26_20_0;
	wire horizontal_tile_26_21_to_tile_26_20_1;
	wire horizontal_tile_26_21_to_tile_26_20_2;
	wire horizontal_tile_26_21_to_tile_26_20_3;

	wire horizontal_tile_27_20_to_tile_27_21_0;
	wire horizontal_tile_27_20_to_tile_27_21_1;
	wire horizontal_tile_27_20_to_tile_27_21_2;
	wire horizontal_tile_27_20_to_tile_27_21_3;
	wire horizontal_tile_27_21_to_tile_27_20_0;
	wire horizontal_tile_27_21_to_tile_27_20_1;
	wire horizontal_tile_27_21_to_tile_27_20_2;
	wire horizontal_tile_27_21_to_tile_27_20_3;

	wire horizontal_tile_28_20_to_tile_28_21_0;
	wire horizontal_tile_28_20_to_tile_28_21_1;
	wire horizontal_tile_28_20_to_tile_28_21_2;
	wire horizontal_tile_28_20_to_tile_28_21_3;
	wire horizontal_tile_28_21_to_tile_28_20_0;
	wire horizontal_tile_28_21_to_tile_28_20_1;
	wire horizontal_tile_28_21_to_tile_28_20_2;
	wire horizontal_tile_28_21_to_tile_28_20_3;

	wire horizontal_tile_29_20_to_tile_29_21_0;
	wire horizontal_tile_29_20_to_tile_29_21_1;
	wire horizontal_tile_29_20_to_tile_29_21_2;
	wire horizontal_tile_29_20_to_tile_29_21_3;
	wire horizontal_tile_29_21_to_tile_29_20_0;
	wire horizontal_tile_29_21_to_tile_29_20_1;
	wire horizontal_tile_29_21_to_tile_29_20_2;
	wire horizontal_tile_29_21_to_tile_29_20_3;

	wire horizontal_tile_30_20_to_tile_30_21_0;
	wire horizontal_tile_30_20_to_tile_30_21_1;
	wire horizontal_tile_30_20_to_tile_30_21_2;
	wire horizontal_tile_30_20_to_tile_30_21_3;
	wire horizontal_tile_30_21_to_tile_30_20_0;
	wire horizontal_tile_30_21_to_tile_30_20_1;
	wire horizontal_tile_30_21_to_tile_30_20_2;
	wire horizontal_tile_30_21_to_tile_30_20_3;

	wire horizontal_tile_31_20_to_tile_31_21_0;
	wire horizontal_tile_31_20_to_tile_31_21_1;
	wire horizontal_tile_31_20_to_tile_31_21_2;
	wire horizontal_tile_31_20_to_tile_31_21_3;
	wire horizontal_tile_31_21_to_tile_31_20_0;
	wire horizontal_tile_31_21_to_tile_31_20_1;
	wire horizontal_tile_31_21_to_tile_31_20_2;
	wire horizontal_tile_31_21_to_tile_31_20_3;

	wire horizontal_tile_0_21_to_tile_0_22_0;
	wire horizontal_tile_0_21_to_tile_0_22_1;
	wire horizontal_tile_0_21_to_tile_0_22_2;
	wire horizontal_tile_0_21_to_tile_0_22_3;
	wire horizontal_tile_0_22_to_tile_0_21_0;
	wire horizontal_tile_0_22_to_tile_0_21_1;
	wire horizontal_tile_0_22_to_tile_0_21_2;
	wire horizontal_tile_0_22_to_tile_0_21_3;

	wire horizontal_tile_1_21_to_tile_1_22_0;
	wire horizontal_tile_1_21_to_tile_1_22_1;
	wire horizontal_tile_1_21_to_tile_1_22_2;
	wire horizontal_tile_1_21_to_tile_1_22_3;
	wire horizontal_tile_1_22_to_tile_1_21_0;
	wire horizontal_tile_1_22_to_tile_1_21_1;
	wire horizontal_tile_1_22_to_tile_1_21_2;
	wire horizontal_tile_1_22_to_tile_1_21_3;

	wire horizontal_tile_2_21_to_tile_2_22_0;
	wire horizontal_tile_2_21_to_tile_2_22_1;
	wire horizontal_tile_2_21_to_tile_2_22_2;
	wire horizontal_tile_2_21_to_tile_2_22_3;
	wire horizontal_tile_2_22_to_tile_2_21_0;
	wire horizontal_tile_2_22_to_tile_2_21_1;
	wire horizontal_tile_2_22_to_tile_2_21_2;
	wire horizontal_tile_2_22_to_tile_2_21_3;

	wire horizontal_tile_3_21_to_tile_3_22_0;
	wire horizontal_tile_3_21_to_tile_3_22_1;
	wire horizontal_tile_3_21_to_tile_3_22_2;
	wire horizontal_tile_3_21_to_tile_3_22_3;
	wire horizontal_tile_3_22_to_tile_3_21_0;
	wire horizontal_tile_3_22_to_tile_3_21_1;
	wire horizontal_tile_3_22_to_tile_3_21_2;
	wire horizontal_tile_3_22_to_tile_3_21_3;

	wire horizontal_tile_4_21_to_tile_4_22_0;
	wire horizontal_tile_4_21_to_tile_4_22_1;
	wire horizontal_tile_4_21_to_tile_4_22_2;
	wire horizontal_tile_4_21_to_tile_4_22_3;
	wire horizontal_tile_4_22_to_tile_4_21_0;
	wire horizontal_tile_4_22_to_tile_4_21_1;
	wire horizontal_tile_4_22_to_tile_4_21_2;
	wire horizontal_tile_4_22_to_tile_4_21_3;

	wire horizontal_tile_5_21_to_tile_5_22_0;
	wire horizontal_tile_5_21_to_tile_5_22_1;
	wire horizontal_tile_5_21_to_tile_5_22_2;
	wire horizontal_tile_5_21_to_tile_5_22_3;
	wire horizontal_tile_5_22_to_tile_5_21_0;
	wire horizontal_tile_5_22_to_tile_5_21_1;
	wire horizontal_tile_5_22_to_tile_5_21_2;
	wire horizontal_tile_5_22_to_tile_5_21_3;

	wire horizontal_tile_6_21_to_tile_6_22_0;
	wire horizontal_tile_6_21_to_tile_6_22_1;
	wire horizontal_tile_6_21_to_tile_6_22_2;
	wire horizontal_tile_6_21_to_tile_6_22_3;
	wire horizontal_tile_6_22_to_tile_6_21_0;
	wire horizontal_tile_6_22_to_tile_6_21_1;
	wire horizontal_tile_6_22_to_tile_6_21_2;
	wire horizontal_tile_6_22_to_tile_6_21_3;

	wire horizontal_tile_7_21_to_tile_7_22_0;
	wire horizontal_tile_7_21_to_tile_7_22_1;
	wire horizontal_tile_7_21_to_tile_7_22_2;
	wire horizontal_tile_7_21_to_tile_7_22_3;
	wire horizontal_tile_7_22_to_tile_7_21_0;
	wire horizontal_tile_7_22_to_tile_7_21_1;
	wire horizontal_tile_7_22_to_tile_7_21_2;
	wire horizontal_tile_7_22_to_tile_7_21_3;

	wire horizontal_tile_8_21_to_tile_8_22_0;
	wire horizontal_tile_8_21_to_tile_8_22_1;
	wire horizontal_tile_8_21_to_tile_8_22_2;
	wire horizontal_tile_8_21_to_tile_8_22_3;
	wire horizontal_tile_8_22_to_tile_8_21_0;
	wire horizontal_tile_8_22_to_tile_8_21_1;
	wire horizontal_tile_8_22_to_tile_8_21_2;
	wire horizontal_tile_8_22_to_tile_8_21_3;

	wire horizontal_tile_9_21_to_tile_9_22_0;
	wire horizontal_tile_9_21_to_tile_9_22_1;
	wire horizontal_tile_9_21_to_tile_9_22_2;
	wire horizontal_tile_9_21_to_tile_9_22_3;
	wire horizontal_tile_9_22_to_tile_9_21_0;
	wire horizontal_tile_9_22_to_tile_9_21_1;
	wire horizontal_tile_9_22_to_tile_9_21_2;
	wire horizontal_tile_9_22_to_tile_9_21_3;

	wire horizontal_tile_10_21_to_tile_10_22_0;
	wire horizontal_tile_10_21_to_tile_10_22_1;
	wire horizontal_tile_10_21_to_tile_10_22_2;
	wire horizontal_tile_10_21_to_tile_10_22_3;
	wire horizontal_tile_10_22_to_tile_10_21_0;
	wire horizontal_tile_10_22_to_tile_10_21_1;
	wire horizontal_tile_10_22_to_tile_10_21_2;
	wire horizontal_tile_10_22_to_tile_10_21_3;

	wire horizontal_tile_11_21_to_tile_11_22_0;
	wire horizontal_tile_11_21_to_tile_11_22_1;
	wire horizontal_tile_11_21_to_tile_11_22_2;
	wire horizontal_tile_11_21_to_tile_11_22_3;
	wire horizontal_tile_11_22_to_tile_11_21_0;
	wire horizontal_tile_11_22_to_tile_11_21_1;
	wire horizontal_tile_11_22_to_tile_11_21_2;
	wire horizontal_tile_11_22_to_tile_11_21_3;

	wire horizontal_tile_12_21_to_tile_12_22_0;
	wire horizontal_tile_12_21_to_tile_12_22_1;
	wire horizontal_tile_12_21_to_tile_12_22_2;
	wire horizontal_tile_12_21_to_tile_12_22_3;
	wire horizontal_tile_12_22_to_tile_12_21_0;
	wire horizontal_tile_12_22_to_tile_12_21_1;
	wire horizontal_tile_12_22_to_tile_12_21_2;
	wire horizontal_tile_12_22_to_tile_12_21_3;

	wire horizontal_tile_13_21_to_tile_13_22_0;
	wire horizontal_tile_13_21_to_tile_13_22_1;
	wire horizontal_tile_13_21_to_tile_13_22_2;
	wire horizontal_tile_13_21_to_tile_13_22_3;
	wire horizontal_tile_13_22_to_tile_13_21_0;
	wire horizontal_tile_13_22_to_tile_13_21_1;
	wire horizontal_tile_13_22_to_tile_13_21_2;
	wire horizontal_tile_13_22_to_tile_13_21_3;

	wire horizontal_tile_14_21_to_tile_14_22_0;
	wire horizontal_tile_14_21_to_tile_14_22_1;
	wire horizontal_tile_14_21_to_tile_14_22_2;
	wire horizontal_tile_14_21_to_tile_14_22_3;
	wire horizontal_tile_14_22_to_tile_14_21_0;
	wire horizontal_tile_14_22_to_tile_14_21_1;
	wire horizontal_tile_14_22_to_tile_14_21_2;
	wire horizontal_tile_14_22_to_tile_14_21_3;

	wire horizontal_tile_15_21_to_tile_15_22_0;
	wire horizontal_tile_15_21_to_tile_15_22_1;
	wire horizontal_tile_15_21_to_tile_15_22_2;
	wire horizontal_tile_15_21_to_tile_15_22_3;
	wire horizontal_tile_15_22_to_tile_15_21_0;
	wire horizontal_tile_15_22_to_tile_15_21_1;
	wire horizontal_tile_15_22_to_tile_15_21_2;
	wire horizontal_tile_15_22_to_tile_15_21_3;

	wire horizontal_tile_16_21_to_tile_16_22_0;
	wire horizontal_tile_16_21_to_tile_16_22_1;
	wire horizontal_tile_16_21_to_tile_16_22_2;
	wire horizontal_tile_16_21_to_tile_16_22_3;
	wire horizontal_tile_16_22_to_tile_16_21_0;
	wire horizontal_tile_16_22_to_tile_16_21_1;
	wire horizontal_tile_16_22_to_tile_16_21_2;
	wire horizontal_tile_16_22_to_tile_16_21_3;

	wire horizontal_tile_17_21_to_tile_17_22_0;
	wire horizontal_tile_17_21_to_tile_17_22_1;
	wire horizontal_tile_17_21_to_tile_17_22_2;
	wire horizontal_tile_17_21_to_tile_17_22_3;
	wire horizontal_tile_17_22_to_tile_17_21_0;
	wire horizontal_tile_17_22_to_tile_17_21_1;
	wire horizontal_tile_17_22_to_tile_17_21_2;
	wire horizontal_tile_17_22_to_tile_17_21_3;

	wire horizontal_tile_18_21_to_tile_18_22_0;
	wire horizontal_tile_18_21_to_tile_18_22_1;
	wire horizontal_tile_18_21_to_tile_18_22_2;
	wire horizontal_tile_18_21_to_tile_18_22_3;
	wire horizontal_tile_18_22_to_tile_18_21_0;
	wire horizontal_tile_18_22_to_tile_18_21_1;
	wire horizontal_tile_18_22_to_tile_18_21_2;
	wire horizontal_tile_18_22_to_tile_18_21_3;

	wire horizontal_tile_19_21_to_tile_19_22_0;
	wire horizontal_tile_19_21_to_tile_19_22_1;
	wire horizontal_tile_19_21_to_tile_19_22_2;
	wire horizontal_tile_19_21_to_tile_19_22_3;
	wire horizontal_tile_19_22_to_tile_19_21_0;
	wire horizontal_tile_19_22_to_tile_19_21_1;
	wire horizontal_tile_19_22_to_tile_19_21_2;
	wire horizontal_tile_19_22_to_tile_19_21_3;

	wire horizontal_tile_20_21_to_tile_20_22_0;
	wire horizontal_tile_20_21_to_tile_20_22_1;
	wire horizontal_tile_20_21_to_tile_20_22_2;
	wire horizontal_tile_20_21_to_tile_20_22_3;
	wire horizontal_tile_20_22_to_tile_20_21_0;
	wire horizontal_tile_20_22_to_tile_20_21_1;
	wire horizontal_tile_20_22_to_tile_20_21_2;
	wire horizontal_tile_20_22_to_tile_20_21_3;

	wire horizontal_tile_21_21_to_tile_21_22_0;
	wire horizontal_tile_21_21_to_tile_21_22_1;
	wire horizontal_tile_21_21_to_tile_21_22_2;
	wire horizontal_tile_21_21_to_tile_21_22_3;
	wire horizontal_tile_21_22_to_tile_21_21_0;
	wire horizontal_tile_21_22_to_tile_21_21_1;
	wire horizontal_tile_21_22_to_tile_21_21_2;
	wire horizontal_tile_21_22_to_tile_21_21_3;

	wire horizontal_tile_22_21_to_tile_22_22_0;
	wire horizontal_tile_22_21_to_tile_22_22_1;
	wire horizontal_tile_22_21_to_tile_22_22_2;
	wire horizontal_tile_22_21_to_tile_22_22_3;
	wire horizontal_tile_22_22_to_tile_22_21_0;
	wire horizontal_tile_22_22_to_tile_22_21_1;
	wire horizontal_tile_22_22_to_tile_22_21_2;
	wire horizontal_tile_22_22_to_tile_22_21_3;

	wire horizontal_tile_23_21_to_tile_23_22_0;
	wire horizontal_tile_23_21_to_tile_23_22_1;
	wire horizontal_tile_23_21_to_tile_23_22_2;
	wire horizontal_tile_23_21_to_tile_23_22_3;
	wire horizontal_tile_23_22_to_tile_23_21_0;
	wire horizontal_tile_23_22_to_tile_23_21_1;
	wire horizontal_tile_23_22_to_tile_23_21_2;
	wire horizontal_tile_23_22_to_tile_23_21_3;

	wire horizontal_tile_24_21_to_tile_24_22_0;
	wire horizontal_tile_24_21_to_tile_24_22_1;
	wire horizontal_tile_24_21_to_tile_24_22_2;
	wire horizontal_tile_24_21_to_tile_24_22_3;
	wire horizontal_tile_24_22_to_tile_24_21_0;
	wire horizontal_tile_24_22_to_tile_24_21_1;
	wire horizontal_tile_24_22_to_tile_24_21_2;
	wire horizontal_tile_24_22_to_tile_24_21_3;

	wire horizontal_tile_25_21_to_tile_25_22_0;
	wire horizontal_tile_25_21_to_tile_25_22_1;
	wire horizontal_tile_25_21_to_tile_25_22_2;
	wire horizontal_tile_25_21_to_tile_25_22_3;
	wire horizontal_tile_25_22_to_tile_25_21_0;
	wire horizontal_tile_25_22_to_tile_25_21_1;
	wire horizontal_tile_25_22_to_tile_25_21_2;
	wire horizontal_tile_25_22_to_tile_25_21_3;

	wire horizontal_tile_26_21_to_tile_26_22_0;
	wire horizontal_tile_26_21_to_tile_26_22_1;
	wire horizontal_tile_26_21_to_tile_26_22_2;
	wire horizontal_tile_26_21_to_tile_26_22_3;
	wire horizontal_tile_26_22_to_tile_26_21_0;
	wire horizontal_tile_26_22_to_tile_26_21_1;
	wire horizontal_tile_26_22_to_tile_26_21_2;
	wire horizontal_tile_26_22_to_tile_26_21_3;

	wire horizontal_tile_27_21_to_tile_27_22_0;
	wire horizontal_tile_27_21_to_tile_27_22_1;
	wire horizontal_tile_27_21_to_tile_27_22_2;
	wire horizontal_tile_27_21_to_tile_27_22_3;
	wire horizontal_tile_27_22_to_tile_27_21_0;
	wire horizontal_tile_27_22_to_tile_27_21_1;
	wire horizontal_tile_27_22_to_tile_27_21_2;
	wire horizontal_tile_27_22_to_tile_27_21_3;

	wire horizontal_tile_28_21_to_tile_28_22_0;
	wire horizontal_tile_28_21_to_tile_28_22_1;
	wire horizontal_tile_28_21_to_tile_28_22_2;
	wire horizontal_tile_28_21_to_tile_28_22_3;
	wire horizontal_tile_28_22_to_tile_28_21_0;
	wire horizontal_tile_28_22_to_tile_28_21_1;
	wire horizontal_tile_28_22_to_tile_28_21_2;
	wire horizontal_tile_28_22_to_tile_28_21_3;

	wire horizontal_tile_29_21_to_tile_29_22_0;
	wire horizontal_tile_29_21_to_tile_29_22_1;
	wire horizontal_tile_29_21_to_tile_29_22_2;
	wire horizontal_tile_29_21_to_tile_29_22_3;
	wire horizontal_tile_29_22_to_tile_29_21_0;
	wire horizontal_tile_29_22_to_tile_29_21_1;
	wire horizontal_tile_29_22_to_tile_29_21_2;
	wire horizontal_tile_29_22_to_tile_29_21_3;

	wire horizontal_tile_30_21_to_tile_30_22_0;
	wire horizontal_tile_30_21_to_tile_30_22_1;
	wire horizontal_tile_30_21_to_tile_30_22_2;
	wire horizontal_tile_30_21_to_tile_30_22_3;
	wire horizontal_tile_30_22_to_tile_30_21_0;
	wire horizontal_tile_30_22_to_tile_30_21_1;
	wire horizontal_tile_30_22_to_tile_30_21_2;
	wire horizontal_tile_30_22_to_tile_30_21_3;

	wire horizontal_tile_31_21_to_tile_31_22_0;
	wire horizontal_tile_31_21_to_tile_31_22_1;
	wire horizontal_tile_31_21_to_tile_31_22_2;
	wire horizontal_tile_31_21_to_tile_31_22_3;
	wire horizontal_tile_31_22_to_tile_31_21_0;
	wire horizontal_tile_31_22_to_tile_31_21_1;
	wire horizontal_tile_31_22_to_tile_31_21_2;
	wire horizontal_tile_31_22_to_tile_31_21_3;

	wire horizontal_tile_0_22_to_tile_0_23_0;
	wire horizontal_tile_0_22_to_tile_0_23_1;
	wire horizontal_tile_0_22_to_tile_0_23_2;
	wire horizontal_tile_0_22_to_tile_0_23_3;
	wire horizontal_tile_0_23_to_tile_0_22_0;
	wire horizontal_tile_0_23_to_tile_0_22_1;
	wire horizontal_tile_0_23_to_tile_0_22_2;
	wire horizontal_tile_0_23_to_tile_0_22_3;

	wire horizontal_tile_1_22_to_tile_1_23_0;
	wire horizontal_tile_1_22_to_tile_1_23_1;
	wire horizontal_tile_1_22_to_tile_1_23_2;
	wire horizontal_tile_1_22_to_tile_1_23_3;
	wire horizontal_tile_1_23_to_tile_1_22_0;
	wire horizontal_tile_1_23_to_tile_1_22_1;
	wire horizontal_tile_1_23_to_tile_1_22_2;
	wire horizontal_tile_1_23_to_tile_1_22_3;

	wire horizontal_tile_2_22_to_tile_2_23_0;
	wire horizontal_tile_2_22_to_tile_2_23_1;
	wire horizontal_tile_2_22_to_tile_2_23_2;
	wire horizontal_tile_2_22_to_tile_2_23_3;
	wire horizontal_tile_2_23_to_tile_2_22_0;
	wire horizontal_tile_2_23_to_tile_2_22_1;
	wire horizontal_tile_2_23_to_tile_2_22_2;
	wire horizontal_tile_2_23_to_tile_2_22_3;

	wire horizontal_tile_3_22_to_tile_3_23_0;
	wire horizontal_tile_3_22_to_tile_3_23_1;
	wire horizontal_tile_3_22_to_tile_3_23_2;
	wire horizontal_tile_3_22_to_tile_3_23_3;
	wire horizontal_tile_3_23_to_tile_3_22_0;
	wire horizontal_tile_3_23_to_tile_3_22_1;
	wire horizontal_tile_3_23_to_tile_3_22_2;
	wire horizontal_tile_3_23_to_tile_3_22_3;

	wire horizontal_tile_4_22_to_tile_4_23_0;
	wire horizontal_tile_4_22_to_tile_4_23_1;
	wire horizontal_tile_4_22_to_tile_4_23_2;
	wire horizontal_tile_4_22_to_tile_4_23_3;
	wire horizontal_tile_4_23_to_tile_4_22_0;
	wire horizontal_tile_4_23_to_tile_4_22_1;
	wire horizontal_tile_4_23_to_tile_4_22_2;
	wire horizontal_tile_4_23_to_tile_4_22_3;

	wire horizontal_tile_5_22_to_tile_5_23_0;
	wire horizontal_tile_5_22_to_tile_5_23_1;
	wire horizontal_tile_5_22_to_tile_5_23_2;
	wire horizontal_tile_5_22_to_tile_5_23_3;
	wire horizontal_tile_5_23_to_tile_5_22_0;
	wire horizontal_tile_5_23_to_tile_5_22_1;
	wire horizontal_tile_5_23_to_tile_5_22_2;
	wire horizontal_tile_5_23_to_tile_5_22_3;

	wire horizontal_tile_6_22_to_tile_6_23_0;
	wire horizontal_tile_6_22_to_tile_6_23_1;
	wire horizontal_tile_6_22_to_tile_6_23_2;
	wire horizontal_tile_6_22_to_tile_6_23_3;
	wire horizontal_tile_6_23_to_tile_6_22_0;
	wire horizontal_tile_6_23_to_tile_6_22_1;
	wire horizontal_tile_6_23_to_tile_6_22_2;
	wire horizontal_tile_6_23_to_tile_6_22_3;

	wire horizontal_tile_7_22_to_tile_7_23_0;
	wire horizontal_tile_7_22_to_tile_7_23_1;
	wire horizontal_tile_7_22_to_tile_7_23_2;
	wire horizontal_tile_7_22_to_tile_7_23_3;
	wire horizontal_tile_7_23_to_tile_7_22_0;
	wire horizontal_tile_7_23_to_tile_7_22_1;
	wire horizontal_tile_7_23_to_tile_7_22_2;
	wire horizontal_tile_7_23_to_tile_7_22_3;

	wire horizontal_tile_8_22_to_tile_8_23_0;
	wire horizontal_tile_8_22_to_tile_8_23_1;
	wire horizontal_tile_8_22_to_tile_8_23_2;
	wire horizontal_tile_8_22_to_tile_8_23_3;
	wire horizontal_tile_8_23_to_tile_8_22_0;
	wire horizontal_tile_8_23_to_tile_8_22_1;
	wire horizontal_tile_8_23_to_tile_8_22_2;
	wire horizontal_tile_8_23_to_tile_8_22_3;

	wire horizontal_tile_9_22_to_tile_9_23_0;
	wire horizontal_tile_9_22_to_tile_9_23_1;
	wire horizontal_tile_9_22_to_tile_9_23_2;
	wire horizontal_tile_9_22_to_tile_9_23_3;
	wire horizontal_tile_9_23_to_tile_9_22_0;
	wire horizontal_tile_9_23_to_tile_9_22_1;
	wire horizontal_tile_9_23_to_tile_9_22_2;
	wire horizontal_tile_9_23_to_tile_9_22_3;

	wire horizontal_tile_10_22_to_tile_10_23_0;
	wire horizontal_tile_10_22_to_tile_10_23_1;
	wire horizontal_tile_10_22_to_tile_10_23_2;
	wire horizontal_tile_10_22_to_tile_10_23_3;
	wire horizontal_tile_10_23_to_tile_10_22_0;
	wire horizontal_tile_10_23_to_tile_10_22_1;
	wire horizontal_tile_10_23_to_tile_10_22_2;
	wire horizontal_tile_10_23_to_tile_10_22_3;

	wire horizontal_tile_11_22_to_tile_11_23_0;
	wire horizontal_tile_11_22_to_tile_11_23_1;
	wire horizontal_tile_11_22_to_tile_11_23_2;
	wire horizontal_tile_11_22_to_tile_11_23_3;
	wire horizontal_tile_11_23_to_tile_11_22_0;
	wire horizontal_tile_11_23_to_tile_11_22_1;
	wire horizontal_tile_11_23_to_tile_11_22_2;
	wire horizontal_tile_11_23_to_tile_11_22_3;

	wire horizontal_tile_12_22_to_tile_12_23_0;
	wire horizontal_tile_12_22_to_tile_12_23_1;
	wire horizontal_tile_12_22_to_tile_12_23_2;
	wire horizontal_tile_12_22_to_tile_12_23_3;
	wire horizontal_tile_12_23_to_tile_12_22_0;
	wire horizontal_tile_12_23_to_tile_12_22_1;
	wire horizontal_tile_12_23_to_tile_12_22_2;
	wire horizontal_tile_12_23_to_tile_12_22_3;

	wire horizontal_tile_13_22_to_tile_13_23_0;
	wire horizontal_tile_13_22_to_tile_13_23_1;
	wire horizontal_tile_13_22_to_tile_13_23_2;
	wire horizontal_tile_13_22_to_tile_13_23_3;
	wire horizontal_tile_13_23_to_tile_13_22_0;
	wire horizontal_tile_13_23_to_tile_13_22_1;
	wire horizontal_tile_13_23_to_tile_13_22_2;
	wire horizontal_tile_13_23_to_tile_13_22_3;

	wire horizontal_tile_14_22_to_tile_14_23_0;
	wire horizontal_tile_14_22_to_tile_14_23_1;
	wire horizontal_tile_14_22_to_tile_14_23_2;
	wire horizontal_tile_14_22_to_tile_14_23_3;
	wire horizontal_tile_14_23_to_tile_14_22_0;
	wire horizontal_tile_14_23_to_tile_14_22_1;
	wire horizontal_tile_14_23_to_tile_14_22_2;
	wire horizontal_tile_14_23_to_tile_14_22_3;

	wire horizontal_tile_15_22_to_tile_15_23_0;
	wire horizontal_tile_15_22_to_tile_15_23_1;
	wire horizontal_tile_15_22_to_tile_15_23_2;
	wire horizontal_tile_15_22_to_tile_15_23_3;
	wire horizontal_tile_15_23_to_tile_15_22_0;
	wire horizontal_tile_15_23_to_tile_15_22_1;
	wire horizontal_tile_15_23_to_tile_15_22_2;
	wire horizontal_tile_15_23_to_tile_15_22_3;

	wire horizontal_tile_16_22_to_tile_16_23_0;
	wire horizontal_tile_16_22_to_tile_16_23_1;
	wire horizontal_tile_16_22_to_tile_16_23_2;
	wire horizontal_tile_16_22_to_tile_16_23_3;
	wire horizontal_tile_16_23_to_tile_16_22_0;
	wire horizontal_tile_16_23_to_tile_16_22_1;
	wire horizontal_tile_16_23_to_tile_16_22_2;
	wire horizontal_tile_16_23_to_tile_16_22_3;

	wire horizontal_tile_17_22_to_tile_17_23_0;
	wire horizontal_tile_17_22_to_tile_17_23_1;
	wire horizontal_tile_17_22_to_tile_17_23_2;
	wire horizontal_tile_17_22_to_tile_17_23_3;
	wire horizontal_tile_17_23_to_tile_17_22_0;
	wire horizontal_tile_17_23_to_tile_17_22_1;
	wire horizontal_tile_17_23_to_tile_17_22_2;
	wire horizontal_tile_17_23_to_tile_17_22_3;

	wire horizontal_tile_18_22_to_tile_18_23_0;
	wire horizontal_tile_18_22_to_tile_18_23_1;
	wire horizontal_tile_18_22_to_tile_18_23_2;
	wire horizontal_tile_18_22_to_tile_18_23_3;
	wire horizontal_tile_18_23_to_tile_18_22_0;
	wire horizontal_tile_18_23_to_tile_18_22_1;
	wire horizontal_tile_18_23_to_tile_18_22_2;
	wire horizontal_tile_18_23_to_tile_18_22_3;

	wire horizontal_tile_19_22_to_tile_19_23_0;
	wire horizontal_tile_19_22_to_tile_19_23_1;
	wire horizontal_tile_19_22_to_tile_19_23_2;
	wire horizontal_tile_19_22_to_tile_19_23_3;
	wire horizontal_tile_19_23_to_tile_19_22_0;
	wire horizontal_tile_19_23_to_tile_19_22_1;
	wire horizontal_tile_19_23_to_tile_19_22_2;
	wire horizontal_tile_19_23_to_tile_19_22_3;

	wire horizontal_tile_20_22_to_tile_20_23_0;
	wire horizontal_tile_20_22_to_tile_20_23_1;
	wire horizontal_tile_20_22_to_tile_20_23_2;
	wire horizontal_tile_20_22_to_tile_20_23_3;
	wire horizontal_tile_20_23_to_tile_20_22_0;
	wire horizontal_tile_20_23_to_tile_20_22_1;
	wire horizontal_tile_20_23_to_tile_20_22_2;
	wire horizontal_tile_20_23_to_tile_20_22_3;

	wire horizontal_tile_21_22_to_tile_21_23_0;
	wire horizontal_tile_21_22_to_tile_21_23_1;
	wire horizontal_tile_21_22_to_tile_21_23_2;
	wire horizontal_tile_21_22_to_tile_21_23_3;
	wire horizontal_tile_21_23_to_tile_21_22_0;
	wire horizontal_tile_21_23_to_tile_21_22_1;
	wire horizontal_tile_21_23_to_tile_21_22_2;
	wire horizontal_tile_21_23_to_tile_21_22_3;

	wire horizontal_tile_22_22_to_tile_22_23_0;
	wire horizontal_tile_22_22_to_tile_22_23_1;
	wire horizontal_tile_22_22_to_tile_22_23_2;
	wire horizontal_tile_22_22_to_tile_22_23_3;
	wire horizontal_tile_22_23_to_tile_22_22_0;
	wire horizontal_tile_22_23_to_tile_22_22_1;
	wire horizontal_tile_22_23_to_tile_22_22_2;
	wire horizontal_tile_22_23_to_tile_22_22_3;

	wire horizontal_tile_23_22_to_tile_23_23_0;
	wire horizontal_tile_23_22_to_tile_23_23_1;
	wire horizontal_tile_23_22_to_tile_23_23_2;
	wire horizontal_tile_23_22_to_tile_23_23_3;
	wire horizontal_tile_23_23_to_tile_23_22_0;
	wire horizontal_tile_23_23_to_tile_23_22_1;
	wire horizontal_tile_23_23_to_tile_23_22_2;
	wire horizontal_tile_23_23_to_tile_23_22_3;

	wire horizontal_tile_24_22_to_tile_24_23_0;
	wire horizontal_tile_24_22_to_tile_24_23_1;
	wire horizontal_tile_24_22_to_tile_24_23_2;
	wire horizontal_tile_24_22_to_tile_24_23_3;
	wire horizontal_tile_24_23_to_tile_24_22_0;
	wire horizontal_tile_24_23_to_tile_24_22_1;
	wire horizontal_tile_24_23_to_tile_24_22_2;
	wire horizontal_tile_24_23_to_tile_24_22_3;

	wire horizontal_tile_25_22_to_tile_25_23_0;
	wire horizontal_tile_25_22_to_tile_25_23_1;
	wire horizontal_tile_25_22_to_tile_25_23_2;
	wire horizontal_tile_25_22_to_tile_25_23_3;
	wire horizontal_tile_25_23_to_tile_25_22_0;
	wire horizontal_tile_25_23_to_tile_25_22_1;
	wire horizontal_tile_25_23_to_tile_25_22_2;
	wire horizontal_tile_25_23_to_tile_25_22_3;

	wire horizontal_tile_26_22_to_tile_26_23_0;
	wire horizontal_tile_26_22_to_tile_26_23_1;
	wire horizontal_tile_26_22_to_tile_26_23_2;
	wire horizontal_tile_26_22_to_tile_26_23_3;
	wire horizontal_tile_26_23_to_tile_26_22_0;
	wire horizontal_tile_26_23_to_tile_26_22_1;
	wire horizontal_tile_26_23_to_tile_26_22_2;
	wire horizontal_tile_26_23_to_tile_26_22_3;

	wire horizontal_tile_27_22_to_tile_27_23_0;
	wire horizontal_tile_27_22_to_tile_27_23_1;
	wire horizontal_tile_27_22_to_tile_27_23_2;
	wire horizontal_tile_27_22_to_tile_27_23_3;
	wire horizontal_tile_27_23_to_tile_27_22_0;
	wire horizontal_tile_27_23_to_tile_27_22_1;
	wire horizontal_tile_27_23_to_tile_27_22_2;
	wire horizontal_tile_27_23_to_tile_27_22_3;

	wire horizontal_tile_28_22_to_tile_28_23_0;
	wire horizontal_tile_28_22_to_tile_28_23_1;
	wire horizontal_tile_28_22_to_tile_28_23_2;
	wire horizontal_tile_28_22_to_tile_28_23_3;
	wire horizontal_tile_28_23_to_tile_28_22_0;
	wire horizontal_tile_28_23_to_tile_28_22_1;
	wire horizontal_tile_28_23_to_tile_28_22_2;
	wire horizontal_tile_28_23_to_tile_28_22_3;

	wire horizontal_tile_29_22_to_tile_29_23_0;
	wire horizontal_tile_29_22_to_tile_29_23_1;
	wire horizontal_tile_29_22_to_tile_29_23_2;
	wire horizontal_tile_29_22_to_tile_29_23_3;
	wire horizontal_tile_29_23_to_tile_29_22_0;
	wire horizontal_tile_29_23_to_tile_29_22_1;
	wire horizontal_tile_29_23_to_tile_29_22_2;
	wire horizontal_tile_29_23_to_tile_29_22_3;

	wire horizontal_tile_30_22_to_tile_30_23_0;
	wire horizontal_tile_30_22_to_tile_30_23_1;
	wire horizontal_tile_30_22_to_tile_30_23_2;
	wire horizontal_tile_30_22_to_tile_30_23_3;
	wire horizontal_tile_30_23_to_tile_30_22_0;
	wire horizontal_tile_30_23_to_tile_30_22_1;
	wire horizontal_tile_30_23_to_tile_30_22_2;
	wire horizontal_tile_30_23_to_tile_30_22_3;

	wire horizontal_tile_31_22_to_tile_31_23_0;
	wire horizontal_tile_31_22_to_tile_31_23_1;
	wire horizontal_tile_31_22_to_tile_31_23_2;
	wire horizontal_tile_31_22_to_tile_31_23_3;
	wire horizontal_tile_31_23_to_tile_31_22_0;
	wire horizontal_tile_31_23_to_tile_31_22_1;
	wire horizontal_tile_31_23_to_tile_31_22_2;
	wire horizontal_tile_31_23_to_tile_31_22_3;

	wire horizontal_tile_0_23_to_tile_0_24_0;
	wire horizontal_tile_0_23_to_tile_0_24_1;
	wire horizontal_tile_0_23_to_tile_0_24_2;
	wire horizontal_tile_0_23_to_tile_0_24_3;
	wire horizontal_tile_0_24_to_tile_0_23_0;
	wire horizontal_tile_0_24_to_tile_0_23_1;
	wire horizontal_tile_0_24_to_tile_0_23_2;
	wire horizontal_tile_0_24_to_tile_0_23_3;

	wire horizontal_tile_1_23_to_tile_1_24_0;
	wire horizontal_tile_1_23_to_tile_1_24_1;
	wire horizontal_tile_1_23_to_tile_1_24_2;
	wire horizontal_tile_1_23_to_tile_1_24_3;
	wire horizontal_tile_1_24_to_tile_1_23_0;
	wire horizontal_tile_1_24_to_tile_1_23_1;
	wire horizontal_tile_1_24_to_tile_1_23_2;
	wire horizontal_tile_1_24_to_tile_1_23_3;

	wire horizontal_tile_2_23_to_tile_2_24_0;
	wire horizontal_tile_2_23_to_tile_2_24_1;
	wire horizontal_tile_2_23_to_tile_2_24_2;
	wire horizontal_tile_2_23_to_tile_2_24_3;
	wire horizontal_tile_2_24_to_tile_2_23_0;
	wire horizontal_tile_2_24_to_tile_2_23_1;
	wire horizontal_tile_2_24_to_tile_2_23_2;
	wire horizontal_tile_2_24_to_tile_2_23_3;

	wire horizontal_tile_3_23_to_tile_3_24_0;
	wire horizontal_tile_3_23_to_tile_3_24_1;
	wire horizontal_tile_3_23_to_tile_3_24_2;
	wire horizontal_tile_3_23_to_tile_3_24_3;
	wire horizontal_tile_3_24_to_tile_3_23_0;
	wire horizontal_tile_3_24_to_tile_3_23_1;
	wire horizontal_tile_3_24_to_tile_3_23_2;
	wire horizontal_tile_3_24_to_tile_3_23_3;

	wire horizontal_tile_4_23_to_tile_4_24_0;
	wire horizontal_tile_4_23_to_tile_4_24_1;
	wire horizontal_tile_4_23_to_tile_4_24_2;
	wire horizontal_tile_4_23_to_tile_4_24_3;
	wire horizontal_tile_4_24_to_tile_4_23_0;
	wire horizontal_tile_4_24_to_tile_4_23_1;
	wire horizontal_tile_4_24_to_tile_4_23_2;
	wire horizontal_tile_4_24_to_tile_4_23_3;

	wire horizontal_tile_5_23_to_tile_5_24_0;
	wire horizontal_tile_5_23_to_tile_5_24_1;
	wire horizontal_tile_5_23_to_tile_5_24_2;
	wire horizontal_tile_5_23_to_tile_5_24_3;
	wire horizontal_tile_5_24_to_tile_5_23_0;
	wire horizontal_tile_5_24_to_tile_5_23_1;
	wire horizontal_tile_5_24_to_tile_5_23_2;
	wire horizontal_tile_5_24_to_tile_5_23_3;

	wire horizontal_tile_6_23_to_tile_6_24_0;
	wire horizontal_tile_6_23_to_tile_6_24_1;
	wire horizontal_tile_6_23_to_tile_6_24_2;
	wire horizontal_tile_6_23_to_tile_6_24_3;
	wire horizontal_tile_6_24_to_tile_6_23_0;
	wire horizontal_tile_6_24_to_tile_6_23_1;
	wire horizontal_tile_6_24_to_tile_6_23_2;
	wire horizontal_tile_6_24_to_tile_6_23_3;

	wire horizontal_tile_7_23_to_tile_7_24_0;
	wire horizontal_tile_7_23_to_tile_7_24_1;
	wire horizontal_tile_7_23_to_tile_7_24_2;
	wire horizontal_tile_7_23_to_tile_7_24_3;
	wire horizontal_tile_7_24_to_tile_7_23_0;
	wire horizontal_tile_7_24_to_tile_7_23_1;
	wire horizontal_tile_7_24_to_tile_7_23_2;
	wire horizontal_tile_7_24_to_tile_7_23_3;

	wire horizontal_tile_8_23_to_tile_8_24_0;
	wire horizontal_tile_8_23_to_tile_8_24_1;
	wire horizontal_tile_8_23_to_tile_8_24_2;
	wire horizontal_tile_8_23_to_tile_8_24_3;
	wire horizontal_tile_8_24_to_tile_8_23_0;
	wire horizontal_tile_8_24_to_tile_8_23_1;
	wire horizontal_tile_8_24_to_tile_8_23_2;
	wire horizontal_tile_8_24_to_tile_8_23_3;

	wire horizontal_tile_9_23_to_tile_9_24_0;
	wire horizontal_tile_9_23_to_tile_9_24_1;
	wire horizontal_tile_9_23_to_tile_9_24_2;
	wire horizontal_tile_9_23_to_tile_9_24_3;
	wire horizontal_tile_9_24_to_tile_9_23_0;
	wire horizontal_tile_9_24_to_tile_9_23_1;
	wire horizontal_tile_9_24_to_tile_9_23_2;
	wire horizontal_tile_9_24_to_tile_9_23_3;

	wire horizontal_tile_10_23_to_tile_10_24_0;
	wire horizontal_tile_10_23_to_tile_10_24_1;
	wire horizontal_tile_10_23_to_tile_10_24_2;
	wire horizontal_tile_10_23_to_tile_10_24_3;
	wire horizontal_tile_10_24_to_tile_10_23_0;
	wire horizontal_tile_10_24_to_tile_10_23_1;
	wire horizontal_tile_10_24_to_tile_10_23_2;
	wire horizontal_tile_10_24_to_tile_10_23_3;

	wire horizontal_tile_11_23_to_tile_11_24_0;
	wire horizontal_tile_11_23_to_tile_11_24_1;
	wire horizontal_tile_11_23_to_tile_11_24_2;
	wire horizontal_tile_11_23_to_tile_11_24_3;
	wire horizontal_tile_11_24_to_tile_11_23_0;
	wire horizontal_tile_11_24_to_tile_11_23_1;
	wire horizontal_tile_11_24_to_tile_11_23_2;
	wire horizontal_tile_11_24_to_tile_11_23_3;

	wire horizontal_tile_12_23_to_tile_12_24_0;
	wire horizontal_tile_12_23_to_tile_12_24_1;
	wire horizontal_tile_12_23_to_tile_12_24_2;
	wire horizontal_tile_12_23_to_tile_12_24_3;
	wire horizontal_tile_12_24_to_tile_12_23_0;
	wire horizontal_tile_12_24_to_tile_12_23_1;
	wire horizontal_tile_12_24_to_tile_12_23_2;
	wire horizontal_tile_12_24_to_tile_12_23_3;

	wire horizontal_tile_13_23_to_tile_13_24_0;
	wire horizontal_tile_13_23_to_tile_13_24_1;
	wire horizontal_tile_13_23_to_tile_13_24_2;
	wire horizontal_tile_13_23_to_tile_13_24_3;
	wire horizontal_tile_13_24_to_tile_13_23_0;
	wire horizontal_tile_13_24_to_tile_13_23_1;
	wire horizontal_tile_13_24_to_tile_13_23_2;
	wire horizontal_tile_13_24_to_tile_13_23_3;

	wire horizontal_tile_14_23_to_tile_14_24_0;
	wire horizontal_tile_14_23_to_tile_14_24_1;
	wire horizontal_tile_14_23_to_tile_14_24_2;
	wire horizontal_tile_14_23_to_tile_14_24_3;
	wire horizontal_tile_14_24_to_tile_14_23_0;
	wire horizontal_tile_14_24_to_tile_14_23_1;
	wire horizontal_tile_14_24_to_tile_14_23_2;
	wire horizontal_tile_14_24_to_tile_14_23_3;

	wire horizontal_tile_15_23_to_tile_15_24_0;
	wire horizontal_tile_15_23_to_tile_15_24_1;
	wire horizontal_tile_15_23_to_tile_15_24_2;
	wire horizontal_tile_15_23_to_tile_15_24_3;
	wire horizontal_tile_15_24_to_tile_15_23_0;
	wire horizontal_tile_15_24_to_tile_15_23_1;
	wire horizontal_tile_15_24_to_tile_15_23_2;
	wire horizontal_tile_15_24_to_tile_15_23_3;

	wire horizontal_tile_16_23_to_tile_16_24_0;
	wire horizontal_tile_16_23_to_tile_16_24_1;
	wire horizontal_tile_16_23_to_tile_16_24_2;
	wire horizontal_tile_16_23_to_tile_16_24_3;
	wire horizontal_tile_16_24_to_tile_16_23_0;
	wire horizontal_tile_16_24_to_tile_16_23_1;
	wire horizontal_tile_16_24_to_tile_16_23_2;
	wire horizontal_tile_16_24_to_tile_16_23_3;

	wire horizontal_tile_17_23_to_tile_17_24_0;
	wire horizontal_tile_17_23_to_tile_17_24_1;
	wire horizontal_tile_17_23_to_tile_17_24_2;
	wire horizontal_tile_17_23_to_tile_17_24_3;
	wire horizontal_tile_17_24_to_tile_17_23_0;
	wire horizontal_tile_17_24_to_tile_17_23_1;
	wire horizontal_tile_17_24_to_tile_17_23_2;
	wire horizontal_tile_17_24_to_tile_17_23_3;

	wire horizontal_tile_18_23_to_tile_18_24_0;
	wire horizontal_tile_18_23_to_tile_18_24_1;
	wire horizontal_tile_18_23_to_tile_18_24_2;
	wire horizontal_tile_18_23_to_tile_18_24_3;
	wire horizontal_tile_18_24_to_tile_18_23_0;
	wire horizontal_tile_18_24_to_tile_18_23_1;
	wire horizontal_tile_18_24_to_tile_18_23_2;
	wire horizontal_tile_18_24_to_tile_18_23_3;

	wire horizontal_tile_19_23_to_tile_19_24_0;
	wire horizontal_tile_19_23_to_tile_19_24_1;
	wire horizontal_tile_19_23_to_tile_19_24_2;
	wire horizontal_tile_19_23_to_tile_19_24_3;
	wire horizontal_tile_19_24_to_tile_19_23_0;
	wire horizontal_tile_19_24_to_tile_19_23_1;
	wire horizontal_tile_19_24_to_tile_19_23_2;
	wire horizontal_tile_19_24_to_tile_19_23_3;

	wire horizontal_tile_20_23_to_tile_20_24_0;
	wire horizontal_tile_20_23_to_tile_20_24_1;
	wire horizontal_tile_20_23_to_tile_20_24_2;
	wire horizontal_tile_20_23_to_tile_20_24_3;
	wire horizontal_tile_20_24_to_tile_20_23_0;
	wire horizontal_tile_20_24_to_tile_20_23_1;
	wire horizontal_tile_20_24_to_tile_20_23_2;
	wire horizontal_tile_20_24_to_tile_20_23_3;

	wire horizontal_tile_21_23_to_tile_21_24_0;
	wire horizontal_tile_21_23_to_tile_21_24_1;
	wire horizontal_tile_21_23_to_tile_21_24_2;
	wire horizontal_tile_21_23_to_tile_21_24_3;
	wire horizontal_tile_21_24_to_tile_21_23_0;
	wire horizontal_tile_21_24_to_tile_21_23_1;
	wire horizontal_tile_21_24_to_tile_21_23_2;
	wire horizontal_tile_21_24_to_tile_21_23_3;

	wire horizontal_tile_22_23_to_tile_22_24_0;
	wire horizontal_tile_22_23_to_tile_22_24_1;
	wire horizontal_tile_22_23_to_tile_22_24_2;
	wire horizontal_tile_22_23_to_tile_22_24_3;
	wire horizontal_tile_22_24_to_tile_22_23_0;
	wire horizontal_tile_22_24_to_tile_22_23_1;
	wire horizontal_tile_22_24_to_tile_22_23_2;
	wire horizontal_tile_22_24_to_tile_22_23_3;

	wire horizontal_tile_23_23_to_tile_23_24_0;
	wire horizontal_tile_23_23_to_tile_23_24_1;
	wire horizontal_tile_23_23_to_tile_23_24_2;
	wire horizontal_tile_23_23_to_tile_23_24_3;
	wire horizontal_tile_23_24_to_tile_23_23_0;
	wire horizontal_tile_23_24_to_tile_23_23_1;
	wire horizontal_tile_23_24_to_tile_23_23_2;
	wire horizontal_tile_23_24_to_tile_23_23_3;

	wire horizontal_tile_24_23_to_tile_24_24_0;
	wire horizontal_tile_24_23_to_tile_24_24_1;
	wire horizontal_tile_24_23_to_tile_24_24_2;
	wire horizontal_tile_24_23_to_tile_24_24_3;
	wire horizontal_tile_24_24_to_tile_24_23_0;
	wire horizontal_tile_24_24_to_tile_24_23_1;
	wire horizontal_tile_24_24_to_tile_24_23_2;
	wire horizontal_tile_24_24_to_tile_24_23_3;

	wire horizontal_tile_25_23_to_tile_25_24_0;
	wire horizontal_tile_25_23_to_tile_25_24_1;
	wire horizontal_tile_25_23_to_tile_25_24_2;
	wire horizontal_tile_25_23_to_tile_25_24_3;
	wire horizontal_tile_25_24_to_tile_25_23_0;
	wire horizontal_tile_25_24_to_tile_25_23_1;
	wire horizontal_tile_25_24_to_tile_25_23_2;
	wire horizontal_tile_25_24_to_tile_25_23_3;

	wire horizontal_tile_26_23_to_tile_26_24_0;
	wire horizontal_tile_26_23_to_tile_26_24_1;
	wire horizontal_tile_26_23_to_tile_26_24_2;
	wire horizontal_tile_26_23_to_tile_26_24_3;
	wire horizontal_tile_26_24_to_tile_26_23_0;
	wire horizontal_tile_26_24_to_tile_26_23_1;
	wire horizontal_tile_26_24_to_tile_26_23_2;
	wire horizontal_tile_26_24_to_tile_26_23_3;

	wire horizontal_tile_27_23_to_tile_27_24_0;
	wire horizontal_tile_27_23_to_tile_27_24_1;
	wire horizontal_tile_27_23_to_tile_27_24_2;
	wire horizontal_tile_27_23_to_tile_27_24_3;
	wire horizontal_tile_27_24_to_tile_27_23_0;
	wire horizontal_tile_27_24_to_tile_27_23_1;
	wire horizontal_tile_27_24_to_tile_27_23_2;
	wire horizontal_tile_27_24_to_tile_27_23_3;

	wire horizontal_tile_28_23_to_tile_28_24_0;
	wire horizontal_tile_28_23_to_tile_28_24_1;
	wire horizontal_tile_28_23_to_tile_28_24_2;
	wire horizontal_tile_28_23_to_tile_28_24_3;
	wire horizontal_tile_28_24_to_tile_28_23_0;
	wire horizontal_tile_28_24_to_tile_28_23_1;
	wire horizontal_tile_28_24_to_tile_28_23_2;
	wire horizontal_tile_28_24_to_tile_28_23_3;

	wire horizontal_tile_29_23_to_tile_29_24_0;
	wire horizontal_tile_29_23_to_tile_29_24_1;
	wire horizontal_tile_29_23_to_tile_29_24_2;
	wire horizontal_tile_29_23_to_tile_29_24_3;
	wire horizontal_tile_29_24_to_tile_29_23_0;
	wire horizontal_tile_29_24_to_tile_29_23_1;
	wire horizontal_tile_29_24_to_tile_29_23_2;
	wire horizontal_tile_29_24_to_tile_29_23_3;

	wire horizontal_tile_30_23_to_tile_30_24_0;
	wire horizontal_tile_30_23_to_tile_30_24_1;
	wire horizontal_tile_30_23_to_tile_30_24_2;
	wire horizontal_tile_30_23_to_tile_30_24_3;
	wire horizontal_tile_30_24_to_tile_30_23_0;
	wire horizontal_tile_30_24_to_tile_30_23_1;
	wire horizontal_tile_30_24_to_tile_30_23_2;
	wire horizontal_tile_30_24_to_tile_30_23_3;

	wire horizontal_tile_31_23_to_tile_31_24_0;
	wire horizontal_tile_31_23_to_tile_31_24_1;
	wire horizontal_tile_31_23_to_tile_31_24_2;
	wire horizontal_tile_31_23_to_tile_31_24_3;
	wire horizontal_tile_31_24_to_tile_31_23_0;
	wire horizontal_tile_31_24_to_tile_31_23_1;
	wire horizontal_tile_31_24_to_tile_31_23_2;
	wire horizontal_tile_31_24_to_tile_31_23_3;

	wire horizontal_tile_0_24_to_tile_0_25_0;
	wire horizontal_tile_0_24_to_tile_0_25_1;
	wire horizontal_tile_0_24_to_tile_0_25_2;
	wire horizontal_tile_0_24_to_tile_0_25_3;
	wire horizontal_tile_0_25_to_tile_0_24_0;
	wire horizontal_tile_0_25_to_tile_0_24_1;
	wire horizontal_tile_0_25_to_tile_0_24_2;
	wire horizontal_tile_0_25_to_tile_0_24_3;

	wire horizontal_tile_1_24_to_tile_1_25_0;
	wire horizontal_tile_1_24_to_tile_1_25_1;
	wire horizontal_tile_1_24_to_tile_1_25_2;
	wire horizontal_tile_1_24_to_tile_1_25_3;
	wire horizontal_tile_1_25_to_tile_1_24_0;
	wire horizontal_tile_1_25_to_tile_1_24_1;
	wire horizontal_tile_1_25_to_tile_1_24_2;
	wire horizontal_tile_1_25_to_tile_1_24_3;

	wire horizontal_tile_2_24_to_tile_2_25_0;
	wire horizontal_tile_2_24_to_tile_2_25_1;
	wire horizontal_tile_2_24_to_tile_2_25_2;
	wire horizontal_tile_2_24_to_tile_2_25_3;
	wire horizontal_tile_2_25_to_tile_2_24_0;
	wire horizontal_tile_2_25_to_tile_2_24_1;
	wire horizontal_tile_2_25_to_tile_2_24_2;
	wire horizontal_tile_2_25_to_tile_2_24_3;

	wire horizontal_tile_3_24_to_tile_3_25_0;
	wire horizontal_tile_3_24_to_tile_3_25_1;
	wire horizontal_tile_3_24_to_tile_3_25_2;
	wire horizontal_tile_3_24_to_tile_3_25_3;
	wire horizontal_tile_3_25_to_tile_3_24_0;
	wire horizontal_tile_3_25_to_tile_3_24_1;
	wire horizontal_tile_3_25_to_tile_3_24_2;
	wire horizontal_tile_3_25_to_tile_3_24_3;

	wire horizontal_tile_4_24_to_tile_4_25_0;
	wire horizontal_tile_4_24_to_tile_4_25_1;
	wire horizontal_tile_4_24_to_tile_4_25_2;
	wire horizontal_tile_4_24_to_tile_4_25_3;
	wire horizontal_tile_4_25_to_tile_4_24_0;
	wire horizontal_tile_4_25_to_tile_4_24_1;
	wire horizontal_tile_4_25_to_tile_4_24_2;
	wire horizontal_tile_4_25_to_tile_4_24_3;

	wire horizontal_tile_5_24_to_tile_5_25_0;
	wire horizontal_tile_5_24_to_tile_5_25_1;
	wire horizontal_tile_5_24_to_tile_5_25_2;
	wire horizontal_tile_5_24_to_tile_5_25_3;
	wire horizontal_tile_5_25_to_tile_5_24_0;
	wire horizontal_tile_5_25_to_tile_5_24_1;
	wire horizontal_tile_5_25_to_tile_5_24_2;
	wire horizontal_tile_5_25_to_tile_5_24_3;

	wire horizontal_tile_6_24_to_tile_6_25_0;
	wire horizontal_tile_6_24_to_tile_6_25_1;
	wire horizontal_tile_6_24_to_tile_6_25_2;
	wire horizontal_tile_6_24_to_tile_6_25_3;
	wire horizontal_tile_6_25_to_tile_6_24_0;
	wire horizontal_tile_6_25_to_tile_6_24_1;
	wire horizontal_tile_6_25_to_tile_6_24_2;
	wire horizontal_tile_6_25_to_tile_6_24_3;

	wire horizontal_tile_7_24_to_tile_7_25_0;
	wire horizontal_tile_7_24_to_tile_7_25_1;
	wire horizontal_tile_7_24_to_tile_7_25_2;
	wire horizontal_tile_7_24_to_tile_7_25_3;
	wire horizontal_tile_7_25_to_tile_7_24_0;
	wire horizontal_tile_7_25_to_tile_7_24_1;
	wire horizontal_tile_7_25_to_tile_7_24_2;
	wire horizontal_tile_7_25_to_tile_7_24_3;

	wire horizontal_tile_8_24_to_tile_8_25_0;
	wire horizontal_tile_8_24_to_tile_8_25_1;
	wire horizontal_tile_8_24_to_tile_8_25_2;
	wire horizontal_tile_8_24_to_tile_8_25_3;
	wire horizontal_tile_8_25_to_tile_8_24_0;
	wire horizontal_tile_8_25_to_tile_8_24_1;
	wire horizontal_tile_8_25_to_tile_8_24_2;
	wire horizontal_tile_8_25_to_tile_8_24_3;

	wire horizontal_tile_9_24_to_tile_9_25_0;
	wire horizontal_tile_9_24_to_tile_9_25_1;
	wire horizontal_tile_9_24_to_tile_9_25_2;
	wire horizontal_tile_9_24_to_tile_9_25_3;
	wire horizontal_tile_9_25_to_tile_9_24_0;
	wire horizontal_tile_9_25_to_tile_9_24_1;
	wire horizontal_tile_9_25_to_tile_9_24_2;
	wire horizontal_tile_9_25_to_tile_9_24_3;

	wire horizontal_tile_10_24_to_tile_10_25_0;
	wire horizontal_tile_10_24_to_tile_10_25_1;
	wire horizontal_tile_10_24_to_tile_10_25_2;
	wire horizontal_tile_10_24_to_tile_10_25_3;
	wire horizontal_tile_10_25_to_tile_10_24_0;
	wire horizontal_tile_10_25_to_tile_10_24_1;
	wire horizontal_tile_10_25_to_tile_10_24_2;
	wire horizontal_tile_10_25_to_tile_10_24_3;

	wire horizontal_tile_11_24_to_tile_11_25_0;
	wire horizontal_tile_11_24_to_tile_11_25_1;
	wire horizontal_tile_11_24_to_tile_11_25_2;
	wire horizontal_tile_11_24_to_tile_11_25_3;
	wire horizontal_tile_11_25_to_tile_11_24_0;
	wire horizontal_tile_11_25_to_tile_11_24_1;
	wire horizontal_tile_11_25_to_tile_11_24_2;
	wire horizontal_tile_11_25_to_tile_11_24_3;

	wire horizontal_tile_12_24_to_tile_12_25_0;
	wire horizontal_tile_12_24_to_tile_12_25_1;
	wire horizontal_tile_12_24_to_tile_12_25_2;
	wire horizontal_tile_12_24_to_tile_12_25_3;
	wire horizontal_tile_12_25_to_tile_12_24_0;
	wire horizontal_tile_12_25_to_tile_12_24_1;
	wire horizontal_tile_12_25_to_tile_12_24_2;
	wire horizontal_tile_12_25_to_tile_12_24_3;

	wire horizontal_tile_13_24_to_tile_13_25_0;
	wire horizontal_tile_13_24_to_tile_13_25_1;
	wire horizontal_tile_13_24_to_tile_13_25_2;
	wire horizontal_tile_13_24_to_tile_13_25_3;
	wire horizontal_tile_13_25_to_tile_13_24_0;
	wire horizontal_tile_13_25_to_tile_13_24_1;
	wire horizontal_tile_13_25_to_tile_13_24_2;
	wire horizontal_tile_13_25_to_tile_13_24_3;

	wire horizontal_tile_14_24_to_tile_14_25_0;
	wire horizontal_tile_14_24_to_tile_14_25_1;
	wire horizontal_tile_14_24_to_tile_14_25_2;
	wire horizontal_tile_14_24_to_tile_14_25_3;
	wire horizontal_tile_14_25_to_tile_14_24_0;
	wire horizontal_tile_14_25_to_tile_14_24_1;
	wire horizontal_tile_14_25_to_tile_14_24_2;
	wire horizontal_tile_14_25_to_tile_14_24_3;

	wire horizontal_tile_15_24_to_tile_15_25_0;
	wire horizontal_tile_15_24_to_tile_15_25_1;
	wire horizontal_tile_15_24_to_tile_15_25_2;
	wire horizontal_tile_15_24_to_tile_15_25_3;
	wire horizontal_tile_15_25_to_tile_15_24_0;
	wire horizontal_tile_15_25_to_tile_15_24_1;
	wire horizontal_tile_15_25_to_tile_15_24_2;
	wire horizontal_tile_15_25_to_tile_15_24_3;

	wire horizontal_tile_16_24_to_tile_16_25_0;
	wire horizontal_tile_16_24_to_tile_16_25_1;
	wire horizontal_tile_16_24_to_tile_16_25_2;
	wire horizontal_tile_16_24_to_tile_16_25_3;
	wire horizontal_tile_16_25_to_tile_16_24_0;
	wire horizontal_tile_16_25_to_tile_16_24_1;
	wire horizontal_tile_16_25_to_tile_16_24_2;
	wire horizontal_tile_16_25_to_tile_16_24_3;

	wire horizontal_tile_17_24_to_tile_17_25_0;
	wire horizontal_tile_17_24_to_tile_17_25_1;
	wire horizontal_tile_17_24_to_tile_17_25_2;
	wire horizontal_tile_17_24_to_tile_17_25_3;
	wire horizontal_tile_17_25_to_tile_17_24_0;
	wire horizontal_tile_17_25_to_tile_17_24_1;
	wire horizontal_tile_17_25_to_tile_17_24_2;
	wire horizontal_tile_17_25_to_tile_17_24_3;

	wire horizontal_tile_18_24_to_tile_18_25_0;
	wire horizontal_tile_18_24_to_tile_18_25_1;
	wire horizontal_tile_18_24_to_tile_18_25_2;
	wire horizontal_tile_18_24_to_tile_18_25_3;
	wire horizontal_tile_18_25_to_tile_18_24_0;
	wire horizontal_tile_18_25_to_tile_18_24_1;
	wire horizontal_tile_18_25_to_tile_18_24_2;
	wire horizontal_tile_18_25_to_tile_18_24_3;

	wire horizontal_tile_19_24_to_tile_19_25_0;
	wire horizontal_tile_19_24_to_tile_19_25_1;
	wire horizontal_tile_19_24_to_tile_19_25_2;
	wire horizontal_tile_19_24_to_tile_19_25_3;
	wire horizontal_tile_19_25_to_tile_19_24_0;
	wire horizontal_tile_19_25_to_tile_19_24_1;
	wire horizontal_tile_19_25_to_tile_19_24_2;
	wire horizontal_tile_19_25_to_tile_19_24_3;

	wire horizontal_tile_20_24_to_tile_20_25_0;
	wire horizontal_tile_20_24_to_tile_20_25_1;
	wire horizontal_tile_20_24_to_tile_20_25_2;
	wire horizontal_tile_20_24_to_tile_20_25_3;
	wire horizontal_tile_20_25_to_tile_20_24_0;
	wire horizontal_tile_20_25_to_tile_20_24_1;
	wire horizontal_tile_20_25_to_tile_20_24_2;
	wire horizontal_tile_20_25_to_tile_20_24_3;

	wire horizontal_tile_21_24_to_tile_21_25_0;
	wire horizontal_tile_21_24_to_tile_21_25_1;
	wire horizontal_tile_21_24_to_tile_21_25_2;
	wire horizontal_tile_21_24_to_tile_21_25_3;
	wire horizontal_tile_21_25_to_tile_21_24_0;
	wire horizontal_tile_21_25_to_tile_21_24_1;
	wire horizontal_tile_21_25_to_tile_21_24_2;
	wire horizontal_tile_21_25_to_tile_21_24_3;

	wire horizontal_tile_22_24_to_tile_22_25_0;
	wire horizontal_tile_22_24_to_tile_22_25_1;
	wire horizontal_tile_22_24_to_tile_22_25_2;
	wire horizontal_tile_22_24_to_tile_22_25_3;
	wire horizontal_tile_22_25_to_tile_22_24_0;
	wire horizontal_tile_22_25_to_tile_22_24_1;
	wire horizontal_tile_22_25_to_tile_22_24_2;
	wire horizontal_tile_22_25_to_tile_22_24_3;

	wire horizontal_tile_23_24_to_tile_23_25_0;
	wire horizontal_tile_23_24_to_tile_23_25_1;
	wire horizontal_tile_23_24_to_tile_23_25_2;
	wire horizontal_tile_23_24_to_tile_23_25_3;
	wire horizontal_tile_23_25_to_tile_23_24_0;
	wire horizontal_tile_23_25_to_tile_23_24_1;
	wire horizontal_tile_23_25_to_tile_23_24_2;
	wire horizontal_tile_23_25_to_tile_23_24_3;

	wire horizontal_tile_24_24_to_tile_24_25_0;
	wire horizontal_tile_24_24_to_tile_24_25_1;
	wire horizontal_tile_24_24_to_tile_24_25_2;
	wire horizontal_tile_24_24_to_tile_24_25_3;
	wire horizontal_tile_24_25_to_tile_24_24_0;
	wire horizontal_tile_24_25_to_tile_24_24_1;
	wire horizontal_tile_24_25_to_tile_24_24_2;
	wire horizontal_tile_24_25_to_tile_24_24_3;

	wire horizontal_tile_25_24_to_tile_25_25_0;
	wire horizontal_tile_25_24_to_tile_25_25_1;
	wire horizontal_tile_25_24_to_tile_25_25_2;
	wire horizontal_tile_25_24_to_tile_25_25_3;
	wire horizontal_tile_25_25_to_tile_25_24_0;
	wire horizontal_tile_25_25_to_tile_25_24_1;
	wire horizontal_tile_25_25_to_tile_25_24_2;
	wire horizontal_tile_25_25_to_tile_25_24_3;

	wire horizontal_tile_26_24_to_tile_26_25_0;
	wire horizontal_tile_26_24_to_tile_26_25_1;
	wire horizontal_tile_26_24_to_tile_26_25_2;
	wire horizontal_tile_26_24_to_tile_26_25_3;
	wire horizontal_tile_26_25_to_tile_26_24_0;
	wire horizontal_tile_26_25_to_tile_26_24_1;
	wire horizontal_tile_26_25_to_tile_26_24_2;
	wire horizontal_tile_26_25_to_tile_26_24_3;

	wire horizontal_tile_27_24_to_tile_27_25_0;
	wire horizontal_tile_27_24_to_tile_27_25_1;
	wire horizontal_tile_27_24_to_tile_27_25_2;
	wire horizontal_tile_27_24_to_tile_27_25_3;
	wire horizontal_tile_27_25_to_tile_27_24_0;
	wire horizontal_tile_27_25_to_tile_27_24_1;
	wire horizontal_tile_27_25_to_tile_27_24_2;
	wire horizontal_tile_27_25_to_tile_27_24_3;

	wire horizontal_tile_28_24_to_tile_28_25_0;
	wire horizontal_tile_28_24_to_tile_28_25_1;
	wire horizontal_tile_28_24_to_tile_28_25_2;
	wire horizontal_tile_28_24_to_tile_28_25_3;
	wire horizontal_tile_28_25_to_tile_28_24_0;
	wire horizontal_tile_28_25_to_tile_28_24_1;
	wire horizontal_tile_28_25_to_tile_28_24_2;
	wire horizontal_tile_28_25_to_tile_28_24_3;

	wire horizontal_tile_29_24_to_tile_29_25_0;
	wire horizontal_tile_29_24_to_tile_29_25_1;
	wire horizontal_tile_29_24_to_tile_29_25_2;
	wire horizontal_tile_29_24_to_tile_29_25_3;
	wire horizontal_tile_29_25_to_tile_29_24_0;
	wire horizontal_tile_29_25_to_tile_29_24_1;
	wire horizontal_tile_29_25_to_tile_29_24_2;
	wire horizontal_tile_29_25_to_tile_29_24_3;

	wire horizontal_tile_30_24_to_tile_30_25_0;
	wire horizontal_tile_30_24_to_tile_30_25_1;
	wire horizontal_tile_30_24_to_tile_30_25_2;
	wire horizontal_tile_30_24_to_tile_30_25_3;
	wire horizontal_tile_30_25_to_tile_30_24_0;
	wire horizontal_tile_30_25_to_tile_30_24_1;
	wire horizontal_tile_30_25_to_tile_30_24_2;
	wire horizontal_tile_30_25_to_tile_30_24_3;

	wire horizontal_tile_31_24_to_tile_31_25_0;
	wire horizontal_tile_31_24_to_tile_31_25_1;
	wire horizontal_tile_31_24_to_tile_31_25_2;
	wire horizontal_tile_31_24_to_tile_31_25_3;
	wire horizontal_tile_31_25_to_tile_31_24_0;
	wire horizontal_tile_31_25_to_tile_31_24_1;
	wire horizontal_tile_31_25_to_tile_31_24_2;
	wire horizontal_tile_31_25_to_tile_31_24_3;

	wire horizontal_tile_0_25_to_tile_0_26_0;
	wire horizontal_tile_0_25_to_tile_0_26_1;
	wire horizontal_tile_0_25_to_tile_0_26_2;
	wire horizontal_tile_0_25_to_tile_0_26_3;
	wire horizontal_tile_0_26_to_tile_0_25_0;
	wire horizontal_tile_0_26_to_tile_0_25_1;
	wire horizontal_tile_0_26_to_tile_0_25_2;
	wire horizontal_tile_0_26_to_tile_0_25_3;

	wire horizontal_tile_1_25_to_tile_1_26_0;
	wire horizontal_tile_1_25_to_tile_1_26_1;
	wire horizontal_tile_1_25_to_tile_1_26_2;
	wire horizontal_tile_1_25_to_tile_1_26_3;
	wire horizontal_tile_1_26_to_tile_1_25_0;
	wire horizontal_tile_1_26_to_tile_1_25_1;
	wire horizontal_tile_1_26_to_tile_1_25_2;
	wire horizontal_tile_1_26_to_tile_1_25_3;

	wire horizontal_tile_2_25_to_tile_2_26_0;
	wire horizontal_tile_2_25_to_tile_2_26_1;
	wire horizontal_tile_2_25_to_tile_2_26_2;
	wire horizontal_tile_2_25_to_tile_2_26_3;
	wire horizontal_tile_2_26_to_tile_2_25_0;
	wire horizontal_tile_2_26_to_tile_2_25_1;
	wire horizontal_tile_2_26_to_tile_2_25_2;
	wire horizontal_tile_2_26_to_tile_2_25_3;

	wire horizontal_tile_3_25_to_tile_3_26_0;
	wire horizontal_tile_3_25_to_tile_3_26_1;
	wire horizontal_tile_3_25_to_tile_3_26_2;
	wire horizontal_tile_3_25_to_tile_3_26_3;
	wire horizontal_tile_3_26_to_tile_3_25_0;
	wire horizontal_tile_3_26_to_tile_3_25_1;
	wire horizontal_tile_3_26_to_tile_3_25_2;
	wire horizontal_tile_3_26_to_tile_3_25_3;

	wire horizontal_tile_4_25_to_tile_4_26_0;
	wire horizontal_tile_4_25_to_tile_4_26_1;
	wire horizontal_tile_4_25_to_tile_4_26_2;
	wire horizontal_tile_4_25_to_tile_4_26_3;
	wire horizontal_tile_4_26_to_tile_4_25_0;
	wire horizontal_tile_4_26_to_tile_4_25_1;
	wire horizontal_tile_4_26_to_tile_4_25_2;
	wire horizontal_tile_4_26_to_tile_4_25_3;

	wire horizontal_tile_5_25_to_tile_5_26_0;
	wire horizontal_tile_5_25_to_tile_5_26_1;
	wire horizontal_tile_5_25_to_tile_5_26_2;
	wire horizontal_tile_5_25_to_tile_5_26_3;
	wire horizontal_tile_5_26_to_tile_5_25_0;
	wire horizontal_tile_5_26_to_tile_5_25_1;
	wire horizontal_tile_5_26_to_tile_5_25_2;
	wire horizontal_tile_5_26_to_tile_5_25_3;

	wire horizontal_tile_6_25_to_tile_6_26_0;
	wire horizontal_tile_6_25_to_tile_6_26_1;
	wire horizontal_tile_6_25_to_tile_6_26_2;
	wire horizontal_tile_6_25_to_tile_6_26_3;
	wire horizontal_tile_6_26_to_tile_6_25_0;
	wire horizontal_tile_6_26_to_tile_6_25_1;
	wire horizontal_tile_6_26_to_tile_6_25_2;
	wire horizontal_tile_6_26_to_tile_6_25_3;

	wire horizontal_tile_7_25_to_tile_7_26_0;
	wire horizontal_tile_7_25_to_tile_7_26_1;
	wire horizontal_tile_7_25_to_tile_7_26_2;
	wire horizontal_tile_7_25_to_tile_7_26_3;
	wire horizontal_tile_7_26_to_tile_7_25_0;
	wire horizontal_tile_7_26_to_tile_7_25_1;
	wire horizontal_tile_7_26_to_tile_7_25_2;
	wire horizontal_tile_7_26_to_tile_7_25_3;

	wire horizontal_tile_8_25_to_tile_8_26_0;
	wire horizontal_tile_8_25_to_tile_8_26_1;
	wire horizontal_tile_8_25_to_tile_8_26_2;
	wire horizontal_tile_8_25_to_tile_8_26_3;
	wire horizontal_tile_8_26_to_tile_8_25_0;
	wire horizontal_tile_8_26_to_tile_8_25_1;
	wire horizontal_tile_8_26_to_tile_8_25_2;
	wire horizontal_tile_8_26_to_tile_8_25_3;

	wire horizontal_tile_9_25_to_tile_9_26_0;
	wire horizontal_tile_9_25_to_tile_9_26_1;
	wire horizontal_tile_9_25_to_tile_9_26_2;
	wire horizontal_tile_9_25_to_tile_9_26_3;
	wire horizontal_tile_9_26_to_tile_9_25_0;
	wire horizontal_tile_9_26_to_tile_9_25_1;
	wire horizontal_tile_9_26_to_tile_9_25_2;
	wire horizontal_tile_9_26_to_tile_9_25_3;

	wire horizontal_tile_10_25_to_tile_10_26_0;
	wire horizontal_tile_10_25_to_tile_10_26_1;
	wire horizontal_tile_10_25_to_tile_10_26_2;
	wire horizontal_tile_10_25_to_tile_10_26_3;
	wire horizontal_tile_10_26_to_tile_10_25_0;
	wire horizontal_tile_10_26_to_tile_10_25_1;
	wire horizontal_tile_10_26_to_tile_10_25_2;
	wire horizontal_tile_10_26_to_tile_10_25_3;

	wire horizontal_tile_11_25_to_tile_11_26_0;
	wire horizontal_tile_11_25_to_tile_11_26_1;
	wire horizontal_tile_11_25_to_tile_11_26_2;
	wire horizontal_tile_11_25_to_tile_11_26_3;
	wire horizontal_tile_11_26_to_tile_11_25_0;
	wire horizontal_tile_11_26_to_tile_11_25_1;
	wire horizontal_tile_11_26_to_tile_11_25_2;
	wire horizontal_tile_11_26_to_tile_11_25_3;

	wire horizontal_tile_12_25_to_tile_12_26_0;
	wire horizontal_tile_12_25_to_tile_12_26_1;
	wire horizontal_tile_12_25_to_tile_12_26_2;
	wire horizontal_tile_12_25_to_tile_12_26_3;
	wire horizontal_tile_12_26_to_tile_12_25_0;
	wire horizontal_tile_12_26_to_tile_12_25_1;
	wire horizontal_tile_12_26_to_tile_12_25_2;
	wire horizontal_tile_12_26_to_tile_12_25_3;

	wire horizontal_tile_13_25_to_tile_13_26_0;
	wire horizontal_tile_13_25_to_tile_13_26_1;
	wire horizontal_tile_13_25_to_tile_13_26_2;
	wire horizontal_tile_13_25_to_tile_13_26_3;
	wire horizontal_tile_13_26_to_tile_13_25_0;
	wire horizontal_tile_13_26_to_tile_13_25_1;
	wire horizontal_tile_13_26_to_tile_13_25_2;
	wire horizontal_tile_13_26_to_tile_13_25_3;

	wire horizontal_tile_14_25_to_tile_14_26_0;
	wire horizontal_tile_14_25_to_tile_14_26_1;
	wire horizontal_tile_14_25_to_tile_14_26_2;
	wire horizontal_tile_14_25_to_tile_14_26_3;
	wire horizontal_tile_14_26_to_tile_14_25_0;
	wire horizontal_tile_14_26_to_tile_14_25_1;
	wire horizontal_tile_14_26_to_tile_14_25_2;
	wire horizontal_tile_14_26_to_tile_14_25_3;

	wire horizontal_tile_15_25_to_tile_15_26_0;
	wire horizontal_tile_15_25_to_tile_15_26_1;
	wire horizontal_tile_15_25_to_tile_15_26_2;
	wire horizontal_tile_15_25_to_tile_15_26_3;
	wire horizontal_tile_15_26_to_tile_15_25_0;
	wire horizontal_tile_15_26_to_tile_15_25_1;
	wire horizontal_tile_15_26_to_tile_15_25_2;
	wire horizontal_tile_15_26_to_tile_15_25_3;

	wire horizontal_tile_16_25_to_tile_16_26_0;
	wire horizontal_tile_16_25_to_tile_16_26_1;
	wire horizontal_tile_16_25_to_tile_16_26_2;
	wire horizontal_tile_16_25_to_tile_16_26_3;
	wire horizontal_tile_16_26_to_tile_16_25_0;
	wire horizontal_tile_16_26_to_tile_16_25_1;
	wire horizontal_tile_16_26_to_tile_16_25_2;
	wire horizontal_tile_16_26_to_tile_16_25_3;

	wire horizontal_tile_17_25_to_tile_17_26_0;
	wire horizontal_tile_17_25_to_tile_17_26_1;
	wire horizontal_tile_17_25_to_tile_17_26_2;
	wire horizontal_tile_17_25_to_tile_17_26_3;
	wire horizontal_tile_17_26_to_tile_17_25_0;
	wire horizontal_tile_17_26_to_tile_17_25_1;
	wire horizontal_tile_17_26_to_tile_17_25_2;
	wire horizontal_tile_17_26_to_tile_17_25_3;

	wire horizontal_tile_18_25_to_tile_18_26_0;
	wire horizontal_tile_18_25_to_tile_18_26_1;
	wire horizontal_tile_18_25_to_tile_18_26_2;
	wire horizontal_tile_18_25_to_tile_18_26_3;
	wire horizontal_tile_18_26_to_tile_18_25_0;
	wire horizontal_tile_18_26_to_tile_18_25_1;
	wire horizontal_tile_18_26_to_tile_18_25_2;
	wire horizontal_tile_18_26_to_tile_18_25_3;

	wire horizontal_tile_19_25_to_tile_19_26_0;
	wire horizontal_tile_19_25_to_tile_19_26_1;
	wire horizontal_tile_19_25_to_tile_19_26_2;
	wire horizontal_tile_19_25_to_tile_19_26_3;
	wire horizontal_tile_19_26_to_tile_19_25_0;
	wire horizontal_tile_19_26_to_tile_19_25_1;
	wire horizontal_tile_19_26_to_tile_19_25_2;
	wire horizontal_tile_19_26_to_tile_19_25_3;

	wire horizontal_tile_20_25_to_tile_20_26_0;
	wire horizontal_tile_20_25_to_tile_20_26_1;
	wire horizontal_tile_20_25_to_tile_20_26_2;
	wire horizontal_tile_20_25_to_tile_20_26_3;
	wire horizontal_tile_20_26_to_tile_20_25_0;
	wire horizontal_tile_20_26_to_tile_20_25_1;
	wire horizontal_tile_20_26_to_tile_20_25_2;
	wire horizontal_tile_20_26_to_tile_20_25_3;

	wire horizontal_tile_21_25_to_tile_21_26_0;
	wire horizontal_tile_21_25_to_tile_21_26_1;
	wire horizontal_tile_21_25_to_tile_21_26_2;
	wire horizontal_tile_21_25_to_tile_21_26_3;
	wire horizontal_tile_21_26_to_tile_21_25_0;
	wire horizontal_tile_21_26_to_tile_21_25_1;
	wire horizontal_tile_21_26_to_tile_21_25_2;
	wire horizontal_tile_21_26_to_tile_21_25_3;

	wire horizontal_tile_22_25_to_tile_22_26_0;
	wire horizontal_tile_22_25_to_tile_22_26_1;
	wire horizontal_tile_22_25_to_tile_22_26_2;
	wire horizontal_tile_22_25_to_tile_22_26_3;
	wire horizontal_tile_22_26_to_tile_22_25_0;
	wire horizontal_tile_22_26_to_tile_22_25_1;
	wire horizontal_tile_22_26_to_tile_22_25_2;
	wire horizontal_tile_22_26_to_tile_22_25_3;

	wire horizontal_tile_23_25_to_tile_23_26_0;
	wire horizontal_tile_23_25_to_tile_23_26_1;
	wire horizontal_tile_23_25_to_tile_23_26_2;
	wire horizontal_tile_23_25_to_tile_23_26_3;
	wire horizontal_tile_23_26_to_tile_23_25_0;
	wire horizontal_tile_23_26_to_tile_23_25_1;
	wire horizontal_tile_23_26_to_tile_23_25_2;
	wire horizontal_tile_23_26_to_tile_23_25_3;

	wire horizontal_tile_24_25_to_tile_24_26_0;
	wire horizontal_tile_24_25_to_tile_24_26_1;
	wire horizontal_tile_24_25_to_tile_24_26_2;
	wire horizontal_tile_24_25_to_tile_24_26_3;
	wire horizontal_tile_24_26_to_tile_24_25_0;
	wire horizontal_tile_24_26_to_tile_24_25_1;
	wire horizontal_tile_24_26_to_tile_24_25_2;
	wire horizontal_tile_24_26_to_tile_24_25_3;

	wire horizontal_tile_25_25_to_tile_25_26_0;
	wire horizontal_tile_25_25_to_tile_25_26_1;
	wire horizontal_tile_25_25_to_tile_25_26_2;
	wire horizontal_tile_25_25_to_tile_25_26_3;
	wire horizontal_tile_25_26_to_tile_25_25_0;
	wire horizontal_tile_25_26_to_tile_25_25_1;
	wire horizontal_tile_25_26_to_tile_25_25_2;
	wire horizontal_tile_25_26_to_tile_25_25_3;

	wire horizontal_tile_26_25_to_tile_26_26_0;
	wire horizontal_tile_26_25_to_tile_26_26_1;
	wire horizontal_tile_26_25_to_tile_26_26_2;
	wire horizontal_tile_26_25_to_tile_26_26_3;
	wire horizontal_tile_26_26_to_tile_26_25_0;
	wire horizontal_tile_26_26_to_tile_26_25_1;
	wire horizontal_tile_26_26_to_tile_26_25_2;
	wire horizontal_tile_26_26_to_tile_26_25_3;

	wire horizontal_tile_27_25_to_tile_27_26_0;
	wire horizontal_tile_27_25_to_tile_27_26_1;
	wire horizontal_tile_27_25_to_tile_27_26_2;
	wire horizontal_tile_27_25_to_tile_27_26_3;
	wire horizontal_tile_27_26_to_tile_27_25_0;
	wire horizontal_tile_27_26_to_tile_27_25_1;
	wire horizontal_tile_27_26_to_tile_27_25_2;
	wire horizontal_tile_27_26_to_tile_27_25_3;

	wire horizontal_tile_28_25_to_tile_28_26_0;
	wire horizontal_tile_28_25_to_tile_28_26_1;
	wire horizontal_tile_28_25_to_tile_28_26_2;
	wire horizontal_tile_28_25_to_tile_28_26_3;
	wire horizontal_tile_28_26_to_tile_28_25_0;
	wire horizontal_tile_28_26_to_tile_28_25_1;
	wire horizontal_tile_28_26_to_tile_28_25_2;
	wire horizontal_tile_28_26_to_tile_28_25_3;

	wire horizontal_tile_29_25_to_tile_29_26_0;
	wire horizontal_tile_29_25_to_tile_29_26_1;
	wire horizontal_tile_29_25_to_tile_29_26_2;
	wire horizontal_tile_29_25_to_tile_29_26_3;
	wire horizontal_tile_29_26_to_tile_29_25_0;
	wire horizontal_tile_29_26_to_tile_29_25_1;
	wire horizontal_tile_29_26_to_tile_29_25_2;
	wire horizontal_tile_29_26_to_tile_29_25_3;

	wire horizontal_tile_30_25_to_tile_30_26_0;
	wire horizontal_tile_30_25_to_tile_30_26_1;
	wire horizontal_tile_30_25_to_tile_30_26_2;
	wire horizontal_tile_30_25_to_tile_30_26_3;
	wire horizontal_tile_30_26_to_tile_30_25_0;
	wire horizontal_tile_30_26_to_tile_30_25_1;
	wire horizontal_tile_30_26_to_tile_30_25_2;
	wire horizontal_tile_30_26_to_tile_30_25_3;

	wire horizontal_tile_31_25_to_tile_31_26_0;
	wire horizontal_tile_31_25_to_tile_31_26_1;
	wire horizontal_tile_31_25_to_tile_31_26_2;
	wire horizontal_tile_31_25_to_tile_31_26_3;
	wire horizontal_tile_31_26_to_tile_31_25_0;
	wire horizontal_tile_31_26_to_tile_31_25_1;
	wire horizontal_tile_31_26_to_tile_31_25_2;
	wire horizontal_tile_31_26_to_tile_31_25_3;

	wire horizontal_tile_0_26_to_tile_0_27_0;
	wire horizontal_tile_0_26_to_tile_0_27_1;
	wire horizontal_tile_0_26_to_tile_0_27_2;
	wire horizontal_tile_0_26_to_tile_0_27_3;
	wire horizontal_tile_0_27_to_tile_0_26_0;
	wire horizontal_tile_0_27_to_tile_0_26_1;
	wire horizontal_tile_0_27_to_tile_0_26_2;
	wire horizontal_tile_0_27_to_tile_0_26_3;

	wire horizontal_tile_1_26_to_tile_1_27_0;
	wire horizontal_tile_1_26_to_tile_1_27_1;
	wire horizontal_tile_1_26_to_tile_1_27_2;
	wire horizontal_tile_1_26_to_tile_1_27_3;
	wire horizontal_tile_1_27_to_tile_1_26_0;
	wire horizontal_tile_1_27_to_tile_1_26_1;
	wire horizontal_tile_1_27_to_tile_1_26_2;
	wire horizontal_tile_1_27_to_tile_1_26_3;

	wire horizontal_tile_2_26_to_tile_2_27_0;
	wire horizontal_tile_2_26_to_tile_2_27_1;
	wire horizontal_tile_2_26_to_tile_2_27_2;
	wire horizontal_tile_2_26_to_tile_2_27_3;
	wire horizontal_tile_2_27_to_tile_2_26_0;
	wire horizontal_tile_2_27_to_tile_2_26_1;
	wire horizontal_tile_2_27_to_tile_2_26_2;
	wire horizontal_tile_2_27_to_tile_2_26_3;

	wire horizontal_tile_3_26_to_tile_3_27_0;
	wire horizontal_tile_3_26_to_tile_3_27_1;
	wire horizontal_tile_3_26_to_tile_3_27_2;
	wire horizontal_tile_3_26_to_tile_3_27_3;
	wire horizontal_tile_3_27_to_tile_3_26_0;
	wire horizontal_tile_3_27_to_tile_3_26_1;
	wire horizontal_tile_3_27_to_tile_3_26_2;
	wire horizontal_tile_3_27_to_tile_3_26_3;

	wire horizontal_tile_4_26_to_tile_4_27_0;
	wire horizontal_tile_4_26_to_tile_4_27_1;
	wire horizontal_tile_4_26_to_tile_4_27_2;
	wire horizontal_tile_4_26_to_tile_4_27_3;
	wire horizontal_tile_4_27_to_tile_4_26_0;
	wire horizontal_tile_4_27_to_tile_4_26_1;
	wire horizontal_tile_4_27_to_tile_4_26_2;
	wire horizontal_tile_4_27_to_tile_4_26_3;

	wire horizontal_tile_5_26_to_tile_5_27_0;
	wire horizontal_tile_5_26_to_tile_5_27_1;
	wire horizontal_tile_5_26_to_tile_5_27_2;
	wire horizontal_tile_5_26_to_tile_5_27_3;
	wire horizontal_tile_5_27_to_tile_5_26_0;
	wire horizontal_tile_5_27_to_tile_5_26_1;
	wire horizontal_tile_5_27_to_tile_5_26_2;
	wire horizontal_tile_5_27_to_tile_5_26_3;

	wire horizontal_tile_6_26_to_tile_6_27_0;
	wire horizontal_tile_6_26_to_tile_6_27_1;
	wire horizontal_tile_6_26_to_tile_6_27_2;
	wire horizontal_tile_6_26_to_tile_6_27_3;
	wire horizontal_tile_6_27_to_tile_6_26_0;
	wire horizontal_tile_6_27_to_tile_6_26_1;
	wire horizontal_tile_6_27_to_tile_6_26_2;
	wire horizontal_tile_6_27_to_tile_6_26_3;

	wire horizontal_tile_7_26_to_tile_7_27_0;
	wire horizontal_tile_7_26_to_tile_7_27_1;
	wire horizontal_tile_7_26_to_tile_7_27_2;
	wire horizontal_tile_7_26_to_tile_7_27_3;
	wire horizontal_tile_7_27_to_tile_7_26_0;
	wire horizontal_tile_7_27_to_tile_7_26_1;
	wire horizontal_tile_7_27_to_tile_7_26_2;
	wire horizontal_tile_7_27_to_tile_7_26_3;

	wire horizontal_tile_8_26_to_tile_8_27_0;
	wire horizontal_tile_8_26_to_tile_8_27_1;
	wire horizontal_tile_8_26_to_tile_8_27_2;
	wire horizontal_tile_8_26_to_tile_8_27_3;
	wire horizontal_tile_8_27_to_tile_8_26_0;
	wire horizontal_tile_8_27_to_tile_8_26_1;
	wire horizontal_tile_8_27_to_tile_8_26_2;
	wire horizontal_tile_8_27_to_tile_8_26_3;

	wire horizontal_tile_9_26_to_tile_9_27_0;
	wire horizontal_tile_9_26_to_tile_9_27_1;
	wire horizontal_tile_9_26_to_tile_9_27_2;
	wire horizontal_tile_9_26_to_tile_9_27_3;
	wire horizontal_tile_9_27_to_tile_9_26_0;
	wire horizontal_tile_9_27_to_tile_9_26_1;
	wire horizontal_tile_9_27_to_tile_9_26_2;
	wire horizontal_tile_9_27_to_tile_9_26_3;

	wire horizontal_tile_10_26_to_tile_10_27_0;
	wire horizontal_tile_10_26_to_tile_10_27_1;
	wire horizontal_tile_10_26_to_tile_10_27_2;
	wire horizontal_tile_10_26_to_tile_10_27_3;
	wire horizontal_tile_10_27_to_tile_10_26_0;
	wire horizontal_tile_10_27_to_tile_10_26_1;
	wire horizontal_tile_10_27_to_tile_10_26_2;
	wire horizontal_tile_10_27_to_tile_10_26_3;

	wire horizontal_tile_11_26_to_tile_11_27_0;
	wire horizontal_tile_11_26_to_tile_11_27_1;
	wire horizontal_tile_11_26_to_tile_11_27_2;
	wire horizontal_tile_11_26_to_tile_11_27_3;
	wire horizontal_tile_11_27_to_tile_11_26_0;
	wire horizontal_tile_11_27_to_tile_11_26_1;
	wire horizontal_tile_11_27_to_tile_11_26_2;
	wire horizontal_tile_11_27_to_tile_11_26_3;

	wire horizontal_tile_12_26_to_tile_12_27_0;
	wire horizontal_tile_12_26_to_tile_12_27_1;
	wire horizontal_tile_12_26_to_tile_12_27_2;
	wire horizontal_tile_12_26_to_tile_12_27_3;
	wire horizontal_tile_12_27_to_tile_12_26_0;
	wire horizontal_tile_12_27_to_tile_12_26_1;
	wire horizontal_tile_12_27_to_tile_12_26_2;
	wire horizontal_tile_12_27_to_tile_12_26_3;

	wire horizontal_tile_13_26_to_tile_13_27_0;
	wire horizontal_tile_13_26_to_tile_13_27_1;
	wire horizontal_tile_13_26_to_tile_13_27_2;
	wire horizontal_tile_13_26_to_tile_13_27_3;
	wire horizontal_tile_13_27_to_tile_13_26_0;
	wire horizontal_tile_13_27_to_tile_13_26_1;
	wire horizontal_tile_13_27_to_tile_13_26_2;
	wire horizontal_tile_13_27_to_tile_13_26_3;

	wire horizontal_tile_14_26_to_tile_14_27_0;
	wire horizontal_tile_14_26_to_tile_14_27_1;
	wire horizontal_tile_14_26_to_tile_14_27_2;
	wire horizontal_tile_14_26_to_tile_14_27_3;
	wire horizontal_tile_14_27_to_tile_14_26_0;
	wire horizontal_tile_14_27_to_tile_14_26_1;
	wire horizontal_tile_14_27_to_tile_14_26_2;
	wire horizontal_tile_14_27_to_tile_14_26_3;

	wire horizontal_tile_15_26_to_tile_15_27_0;
	wire horizontal_tile_15_26_to_tile_15_27_1;
	wire horizontal_tile_15_26_to_tile_15_27_2;
	wire horizontal_tile_15_26_to_tile_15_27_3;
	wire horizontal_tile_15_27_to_tile_15_26_0;
	wire horizontal_tile_15_27_to_tile_15_26_1;
	wire horizontal_tile_15_27_to_tile_15_26_2;
	wire horizontal_tile_15_27_to_tile_15_26_3;

	wire horizontal_tile_16_26_to_tile_16_27_0;
	wire horizontal_tile_16_26_to_tile_16_27_1;
	wire horizontal_tile_16_26_to_tile_16_27_2;
	wire horizontal_tile_16_26_to_tile_16_27_3;
	wire horizontal_tile_16_27_to_tile_16_26_0;
	wire horizontal_tile_16_27_to_tile_16_26_1;
	wire horizontal_tile_16_27_to_tile_16_26_2;
	wire horizontal_tile_16_27_to_tile_16_26_3;

	wire horizontal_tile_17_26_to_tile_17_27_0;
	wire horizontal_tile_17_26_to_tile_17_27_1;
	wire horizontal_tile_17_26_to_tile_17_27_2;
	wire horizontal_tile_17_26_to_tile_17_27_3;
	wire horizontal_tile_17_27_to_tile_17_26_0;
	wire horizontal_tile_17_27_to_tile_17_26_1;
	wire horizontal_tile_17_27_to_tile_17_26_2;
	wire horizontal_tile_17_27_to_tile_17_26_3;

	wire horizontal_tile_18_26_to_tile_18_27_0;
	wire horizontal_tile_18_26_to_tile_18_27_1;
	wire horizontal_tile_18_26_to_tile_18_27_2;
	wire horizontal_tile_18_26_to_tile_18_27_3;
	wire horizontal_tile_18_27_to_tile_18_26_0;
	wire horizontal_tile_18_27_to_tile_18_26_1;
	wire horizontal_tile_18_27_to_tile_18_26_2;
	wire horizontal_tile_18_27_to_tile_18_26_3;

	wire horizontal_tile_19_26_to_tile_19_27_0;
	wire horizontal_tile_19_26_to_tile_19_27_1;
	wire horizontal_tile_19_26_to_tile_19_27_2;
	wire horizontal_tile_19_26_to_tile_19_27_3;
	wire horizontal_tile_19_27_to_tile_19_26_0;
	wire horizontal_tile_19_27_to_tile_19_26_1;
	wire horizontal_tile_19_27_to_tile_19_26_2;
	wire horizontal_tile_19_27_to_tile_19_26_3;

	wire horizontal_tile_20_26_to_tile_20_27_0;
	wire horizontal_tile_20_26_to_tile_20_27_1;
	wire horizontal_tile_20_26_to_tile_20_27_2;
	wire horizontal_tile_20_26_to_tile_20_27_3;
	wire horizontal_tile_20_27_to_tile_20_26_0;
	wire horizontal_tile_20_27_to_tile_20_26_1;
	wire horizontal_tile_20_27_to_tile_20_26_2;
	wire horizontal_tile_20_27_to_tile_20_26_3;

	wire horizontal_tile_21_26_to_tile_21_27_0;
	wire horizontal_tile_21_26_to_tile_21_27_1;
	wire horizontal_tile_21_26_to_tile_21_27_2;
	wire horizontal_tile_21_26_to_tile_21_27_3;
	wire horizontal_tile_21_27_to_tile_21_26_0;
	wire horizontal_tile_21_27_to_tile_21_26_1;
	wire horizontal_tile_21_27_to_tile_21_26_2;
	wire horizontal_tile_21_27_to_tile_21_26_3;

	wire horizontal_tile_22_26_to_tile_22_27_0;
	wire horizontal_tile_22_26_to_tile_22_27_1;
	wire horizontal_tile_22_26_to_tile_22_27_2;
	wire horizontal_tile_22_26_to_tile_22_27_3;
	wire horizontal_tile_22_27_to_tile_22_26_0;
	wire horizontal_tile_22_27_to_tile_22_26_1;
	wire horizontal_tile_22_27_to_tile_22_26_2;
	wire horizontal_tile_22_27_to_tile_22_26_3;

	wire horizontal_tile_23_26_to_tile_23_27_0;
	wire horizontal_tile_23_26_to_tile_23_27_1;
	wire horizontal_tile_23_26_to_tile_23_27_2;
	wire horizontal_tile_23_26_to_tile_23_27_3;
	wire horizontal_tile_23_27_to_tile_23_26_0;
	wire horizontal_tile_23_27_to_tile_23_26_1;
	wire horizontal_tile_23_27_to_tile_23_26_2;
	wire horizontal_tile_23_27_to_tile_23_26_3;

	wire horizontal_tile_24_26_to_tile_24_27_0;
	wire horizontal_tile_24_26_to_tile_24_27_1;
	wire horizontal_tile_24_26_to_tile_24_27_2;
	wire horizontal_tile_24_26_to_tile_24_27_3;
	wire horizontal_tile_24_27_to_tile_24_26_0;
	wire horizontal_tile_24_27_to_tile_24_26_1;
	wire horizontal_tile_24_27_to_tile_24_26_2;
	wire horizontal_tile_24_27_to_tile_24_26_3;

	wire horizontal_tile_25_26_to_tile_25_27_0;
	wire horizontal_tile_25_26_to_tile_25_27_1;
	wire horizontal_tile_25_26_to_tile_25_27_2;
	wire horizontal_tile_25_26_to_tile_25_27_3;
	wire horizontal_tile_25_27_to_tile_25_26_0;
	wire horizontal_tile_25_27_to_tile_25_26_1;
	wire horizontal_tile_25_27_to_tile_25_26_2;
	wire horizontal_tile_25_27_to_tile_25_26_3;

	wire horizontal_tile_26_26_to_tile_26_27_0;
	wire horizontal_tile_26_26_to_tile_26_27_1;
	wire horizontal_tile_26_26_to_tile_26_27_2;
	wire horizontal_tile_26_26_to_tile_26_27_3;
	wire horizontal_tile_26_27_to_tile_26_26_0;
	wire horizontal_tile_26_27_to_tile_26_26_1;
	wire horizontal_tile_26_27_to_tile_26_26_2;
	wire horizontal_tile_26_27_to_tile_26_26_3;

	wire horizontal_tile_27_26_to_tile_27_27_0;
	wire horizontal_tile_27_26_to_tile_27_27_1;
	wire horizontal_tile_27_26_to_tile_27_27_2;
	wire horizontal_tile_27_26_to_tile_27_27_3;
	wire horizontal_tile_27_27_to_tile_27_26_0;
	wire horizontal_tile_27_27_to_tile_27_26_1;
	wire horizontal_tile_27_27_to_tile_27_26_2;
	wire horizontal_tile_27_27_to_tile_27_26_3;

	wire horizontal_tile_28_26_to_tile_28_27_0;
	wire horizontal_tile_28_26_to_tile_28_27_1;
	wire horizontal_tile_28_26_to_tile_28_27_2;
	wire horizontal_tile_28_26_to_tile_28_27_3;
	wire horizontal_tile_28_27_to_tile_28_26_0;
	wire horizontal_tile_28_27_to_tile_28_26_1;
	wire horizontal_tile_28_27_to_tile_28_26_2;
	wire horizontal_tile_28_27_to_tile_28_26_3;

	wire horizontal_tile_29_26_to_tile_29_27_0;
	wire horizontal_tile_29_26_to_tile_29_27_1;
	wire horizontal_tile_29_26_to_tile_29_27_2;
	wire horizontal_tile_29_26_to_tile_29_27_3;
	wire horizontal_tile_29_27_to_tile_29_26_0;
	wire horizontal_tile_29_27_to_tile_29_26_1;
	wire horizontal_tile_29_27_to_tile_29_26_2;
	wire horizontal_tile_29_27_to_tile_29_26_3;

	wire horizontal_tile_30_26_to_tile_30_27_0;
	wire horizontal_tile_30_26_to_tile_30_27_1;
	wire horizontal_tile_30_26_to_tile_30_27_2;
	wire horizontal_tile_30_26_to_tile_30_27_3;
	wire horizontal_tile_30_27_to_tile_30_26_0;
	wire horizontal_tile_30_27_to_tile_30_26_1;
	wire horizontal_tile_30_27_to_tile_30_26_2;
	wire horizontal_tile_30_27_to_tile_30_26_3;

	wire horizontal_tile_31_26_to_tile_31_27_0;
	wire horizontal_tile_31_26_to_tile_31_27_1;
	wire horizontal_tile_31_26_to_tile_31_27_2;
	wire horizontal_tile_31_26_to_tile_31_27_3;
	wire horizontal_tile_31_27_to_tile_31_26_0;
	wire horizontal_tile_31_27_to_tile_31_26_1;
	wire horizontal_tile_31_27_to_tile_31_26_2;
	wire horizontal_tile_31_27_to_tile_31_26_3;

	wire horizontal_tile_0_27_to_tile_0_28_0;
	wire horizontal_tile_0_27_to_tile_0_28_1;
	wire horizontal_tile_0_27_to_tile_0_28_2;
	wire horizontal_tile_0_27_to_tile_0_28_3;
	wire horizontal_tile_0_28_to_tile_0_27_0;
	wire horizontal_tile_0_28_to_tile_0_27_1;
	wire horizontal_tile_0_28_to_tile_0_27_2;
	wire horizontal_tile_0_28_to_tile_0_27_3;

	wire horizontal_tile_1_27_to_tile_1_28_0;
	wire horizontal_tile_1_27_to_tile_1_28_1;
	wire horizontal_tile_1_27_to_tile_1_28_2;
	wire horizontal_tile_1_27_to_tile_1_28_3;
	wire horizontal_tile_1_28_to_tile_1_27_0;
	wire horizontal_tile_1_28_to_tile_1_27_1;
	wire horizontal_tile_1_28_to_tile_1_27_2;
	wire horizontal_tile_1_28_to_tile_1_27_3;

	wire horizontal_tile_2_27_to_tile_2_28_0;
	wire horizontal_tile_2_27_to_tile_2_28_1;
	wire horizontal_tile_2_27_to_tile_2_28_2;
	wire horizontal_tile_2_27_to_tile_2_28_3;
	wire horizontal_tile_2_28_to_tile_2_27_0;
	wire horizontal_tile_2_28_to_tile_2_27_1;
	wire horizontal_tile_2_28_to_tile_2_27_2;
	wire horizontal_tile_2_28_to_tile_2_27_3;

	wire horizontal_tile_3_27_to_tile_3_28_0;
	wire horizontal_tile_3_27_to_tile_3_28_1;
	wire horizontal_tile_3_27_to_tile_3_28_2;
	wire horizontal_tile_3_27_to_tile_3_28_3;
	wire horizontal_tile_3_28_to_tile_3_27_0;
	wire horizontal_tile_3_28_to_tile_3_27_1;
	wire horizontal_tile_3_28_to_tile_3_27_2;
	wire horizontal_tile_3_28_to_tile_3_27_3;

	wire horizontal_tile_4_27_to_tile_4_28_0;
	wire horizontal_tile_4_27_to_tile_4_28_1;
	wire horizontal_tile_4_27_to_tile_4_28_2;
	wire horizontal_tile_4_27_to_tile_4_28_3;
	wire horizontal_tile_4_28_to_tile_4_27_0;
	wire horizontal_tile_4_28_to_tile_4_27_1;
	wire horizontal_tile_4_28_to_tile_4_27_2;
	wire horizontal_tile_4_28_to_tile_4_27_3;

	wire horizontal_tile_5_27_to_tile_5_28_0;
	wire horizontal_tile_5_27_to_tile_5_28_1;
	wire horizontal_tile_5_27_to_tile_5_28_2;
	wire horizontal_tile_5_27_to_tile_5_28_3;
	wire horizontal_tile_5_28_to_tile_5_27_0;
	wire horizontal_tile_5_28_to_tile_5_27_1;
	wire horizontal_tile_5_28_to_tile_5_27_2;
	wire horizontal_tile_5_28_to_tile_5_27_3;

	wire horizontal_tile_6_27_to_tile_6_28_0;
	wire horizontal_tile_6_27_to_tile_6_28_1;
	wire horizontal_tile_6_27_to_tile_6_28_2;
	wire horizontal_tile_6_27_to_tile_6_28_3;
	wire horizontal_tile_6_28_to_tile_6_27_0;
	wire horizontal_tile_6_28_to_tile_6_27_1;
	wire horizontal_tile_6_28_to_tile_6_27_2;
	wire horizontal_tile_6_28_to_tile_6_27_3;

	wire horizontal_tile_7_27_to_tile_7_28_0;
	wire horizontal_tile_7_27_to_tile_7_28_1;
	wire horizontal_tile_7_27_to_tile_7_28_2;
	wire horizontal_tile_7_27_to_tile_7_28_3;
	wire horizontal_tile_7_28_to_tile_7_27_0;
	wire horizontal_tile_7_28_to_tile_7_27_1;
	wire horizontal_tile_7_28_to_tile_7_27_2;
	wire horizontal_tile_7_28_to_tile_7_27_3;

	wire horizontal_tile_8_27_to_tile_8_28_0;
	wire horizontal_tile_8_27_to_tile_8_28_1;
	wire horizontal_tile_8_27_to_tile_8_28_2;
	wire horizontal_tile_8_27_to_tile_8_28_3;
	wire horizontal_tile_8_28_to_tile_8_27_0;
	wire horizontal_tile_8_28_to_tile_8_27_1;
	wire horizontal_tile_8_28_to_tile_8_27_2;
	wire horizontal_tile_8_28_to_tile_8_27_3;

	wire horizontal_tile_9_27_to_tile_9_28_0;
	wire horizontal_tile_9_27_to_tile_9_28_1;
	wire horizontal_tile_9_27_to_tile_9_28_2;
	wire horizontal_tile_9_27_to_tile_9_28_3;
	wire horizontal_tile_9_28_to_tile_9_27_0;
	wire horizontal_tile_9_28_to_tile_9_27_1;
	wire horizontal_tile_9_28_to_tile_9_27_2;
	wire horizontal_tile_9_28_to_tile_9_27_3;

	wire horizontal_tile_10_27_to_tile_10_28_0;
	wire horizontal_tile_10_27_to_tile_10_28_1;
	wire horizontal_tile_10_27_to_tile_10_28_2;
	wire horizontal_tile_10_27_to_tile_10_28_3;
	wire horizontal_tile_10_28_to_tile_10_27_0;
	wire horizontal_tile_10_28_to_tile_10_27_1;
	wire horizontal_tile_10_28_to_tile_10_27_2;
	wire horizontal_tile_10_28_to_tile_10_27_3;

	wire horizontal_tile_11_27_to_tile_11_28_0;
	wire horizontal_tile_11_27_to_tile_11_28_1;
	wire horizontal_tile_11_27_to_tile_11_28_2;
	wire horizontal_tile_11_27_to_tile_11_28_3;
	wire horizontal_tile_11_28_to_tile_11_27_0;
	wire horizontal_tile_11_28_to_tile_11_27_1;
	wire horizontal_tile_11_28_to_tile_11_27_2;
	wire horizontal_tile_11_28_to_tile_11_27_3;

	wire horizontal_tile_12_27_to_tile_12_28_0;
	wire horizontal_tile_12_27_to_tile_12_28_1;
	wire horizontal_tile_12_27_to_tile_12_28_2;
	wire horizontal_tile_12_27_to_tile_12_28_3;
	wire horizontal_tile_12_28_to_tile_12_27_0;
	wire horizontal_tile_12_28_to_tile_12_27_1;
	wire horizontal_tile_12_28_to_tile_12_27_2;
	wire horizontal_tile_12_28_to_tile_12_27_3;

	wire horizontal_tile_13_27_to_tile_13_28_0;
	wire horizontal_tile_13_27_to_tile_13_28_1;
	wire horizontal_tile_13_27_to_tile_13_28_2;
	wire horizontal_tile_13_27_to_tile_13_28_3;
	wire horizontal_tile_13_28_to_tile_13_27_0;
	wire horizontal_tile_13_28_to_tile_13_27_1;
	wire horizontal_tile_13_28_to_tile_13_27_2;
	wire horizontal_tile_13_28_to_tile_13_27_3;

	wire horizontal_tile_14_27_to_tile_14_28_0;
	wire horizontal_tile_14_27_to_tile_14_28_1;
	wire horizontal_tile_14_27_to_tile_14_28_2;
	wire horizontal_tile_14_27_to_tile_14_28_3;
	wire horizontal_tile_14_28_to_tile_14_27_0;
	wire horizontal_tile_14_28_to_tile_14_27_1;
	wire horizontal_tile_14_28_to_tile_14_27_2;
	wire horizontal_tile_14_28_to_tile_14_27_3;

	wire horizontal_tile_15_27_to_tile_15_28_0;
	wire horizontal_tile_15_27_to_tile_15_28_1;
	wire horizontal_tile_15_27_to_tile_15_28_2;
	wire horizontal_tile_15_27_to_tile_15_28_3;
	wire horizontal_tile_15_28_to_tile_15_27_0;
	wire horizontal_tile_15_28_to_tile_15_27_1;
	wire horizontal_tile_15_28_to_tile_15_27_2;
	wire horizontal_tile_15_28_to_tile_15_27_3;

	wire horizontal_tile_16_27_to_tile_16_28_0;
	wire horizontal_tile_16_27_to_tile_16_28_1;
	wire horizontal_tile_16_27_to_tile_16_28_2;
	wire horizontal_tile_16_27_to_tile_16_28_3;
	wire horizontal_tile_16_28_to_tile_16_27_0;
	wire horizontal_tile_16_28_to_tile_16_27_1;
	wire horizontal_tile_16_28_to_tile_16_27_2;
	wire horizontal_tile_16_28_to_tile_16_27_3;

	wire horizontal_tile_17_27_to_tile_17_28_0;
	wire horizontal_tile_17_27_to_tile_17_28_1;
	wire horizontal_tile_17_27_to_tile_17_28_2;
	wire horizontal_tile_17_27_to_tile_17_28_3;
	wire horizontal_tile_17_28_to_tile_17_27_0;
	wire horizontal_tile_17_28_to_tile_17_27_1;
	wire horizontal_tile_17_28_to_tile_17_27_2;
	wire horizontal_tile_17_28_to_tile_17_27_3;

	wire horizontal_tile_18_27_to_tile_18_28_0;
	wire horizontal_tile_18_27_to_tile_18_28_1;
	wire horizontal_tile_18_27_to_tile_18_28_2;
	wire horizontal_tile_18_27_to_tile_18_28_3;
	wire horizontal_tile_18_28_to_tile_18_27_0;
	wire horizontal_tile_18_28_to_tile_18_27_1;
	wire horizontal_tile_18_28_to_tile_18_27_2;
	wire horizontal_tile_18_28_to_tile_18_27_3;

	wire horizontal_tile_19_27_to_tile_19_28_0;
	wire horizontal_tile_19_27_to_tile_19_28_1;
	wire horizontal_tile_19_27_to_tile_19_28_2;
	wire horizontal_tile_19_27_to_tile_19_28_3;
	wire horizontal_tile_19_28_to_tile_19_27_0;
	wire horizontal_tile_19_28_to_tile_19_27_1;
	wire horizontal_tile_19_28_to_tile_19_27_2;
	wire horizontal_tile_19_28_to_tile_19_27_3;

	wire horizontal_tile_20_27_to_tile_20_28_0;
	wire horizontal_tile_20_27_to_tile_20_28_1;
	wire horizontal_tile_20_27_to_tile_20_28_2;
	wire horizontal_tile_20_27_to_tile_20_28_3;
	wire horizontal_tile_20_28_to_tile_20_27_0;
	wire horizontal_tile_20_28_to_tile_20_27_1;
	wire horizontal_tile_20_28_to_tile_20_27_2;
	wire horizontal_tile_20_28_to_tile_20_27_3;

	wire horizontal_tile_21_27_to_tile_21_28_0;
	wire horizontal_tile_21_27_to_tile_21_28_1;
	wire horizontal_tile_21_27_to_tile_21_28_2;
	wire horizontal_tile_21_27_to_tile_21_28_3;
	wire horizontal_tile_21_28_to_tile_21_27_0;
	wire horizontal_tile_21_28_to_tile_21_27_1;
	wire horizontal_tile_21_28_to_tile_21_27_2;
	wire horizontal_tile_21_28_to_tile_21_27_3;

	wire horizontal_tile_22_27_to_tile_22_28_0;
	wire horizontal_tile_22_27_to_tile_22_28_1;
	wire horizontal_tile_22_27_to_tile_22_28_2;
	wire horizontal_tile_22_27_to_tile_22_28_3;
	wire horizontal_tile_22_28_to_tile_22_27_0;
	wire horizontal_tile_22_28_to_tile_22_27_1;
	wire horizontal_tile_22_28_to_tile_22_27_2;
	wire horizontal_tile_22_28_to_tile_22_27_3;

	wire horizontal_tile_23_27_to_tile_23_28_0;
	wire horizontal_tile_23_27_to_tile_23_28_1;
	wire horizontal_tile_23_27_to_tile_23_28_2;
	wire horizontal_tile_23_27_to_tile_23_28_3;
	wire horizontal_tile_23_28_to_tile_23_27_0;
	wire horizontal_tile_23_28_to_tile_23_27_1;
	wire horizontal_tile_23_28_to_tile_23_27_2;
	wire horizontal_tile_23_28_to_tile_23_27_3;

	wire horizontal_tile_24_27_to_tile_24_28_0;
	wire horizontal_tile_24_27_to_tile_24_28_1;
	wire horizontal_tile_24_27_to_tile_24_28_2;
	wire horizontal_tile_24_27_to_tile_24_28_3;
	wire horizontal_tile_24_28_to_tile_24_27_0;
	wire horizontal_tile_24_28_to_tile_24_27_1;
	wire horizontal_tile_24_28_to_tile_24_27_2;
	wire horizontal_tile_24_28_to_tile_24_27_3;

	wire horizontal_tile_25_27_to_tile_25_28_0;
	wire horizontal_tile_25_27_to_tile_25_28_1;
	wire horizontal_tile_25_27_to_tile_25_28_2;
	wire horizontal_tile_25_27_to_tile_25_28_3;
	wire horizontal_tile_25_28_to_tile_25_27_0;
	wire horizontal_tile_25_28_to_tile_25_27_1;
	wire horizontal_tile_25_28_to_tile_25_27_2;
	wire horizontal_tile_25_28_to_tile_25_27_3;

	wire horizontal_tile_26_27_to_tile_26_28_0;
	wire horizontal_tile_26_27_to_tile_26_28_1;
	wire horizontal_tile_26_27_to_tile_26_28_2;
	wire horizontal_tile_26_27_to_tile_26_28_3;
	wire horizontal_tile_26_28_to_tile_26_27_0;
	wire horizontal_tile_26_28_to_tile_26_27_1;
	wire horizontal_tile_26_28_to_tile_26_27_2;
	wire horizontal_tile_26_28_to_tile_26_27_3;

	wire horizontal_tile_27_27_to_tile_27_28_0;
	wire horizontal_tile_27_27_to_tile_27_28_1;
	wire horizontal_tile_27_27_to_tile_27_28_2;
	wire horizontal_tile_27_27_to_tile_27_28_3;
	wire horizontal_tile_27_28_to_tile_27_27_0;
	wire horizontal_tile_27_28_to_tile_27_27_1;
	wire horizontal_tile_27_28_to_tile_27_27_2;
	wire horizontal_tile_27_28_to_tile_27_27_3;

	wire horizontal_tile_28_27_to_tile_28_28_0;
	wire horizontal_tile_28_27_to_tile_28_28_1;
	wire horizontal_tile_28_27_to_tile_28_28_2;
	wire horizontal_tile_28_27_to_tile_28_28_3;
	wire horizontal_tile_28_28_to_tile_28_27_0;
	wire horizontal_tile_28_28_to_tile_28_27_1;
	wire horizontal_tile_28_28_to_tile_28_27_2;
	wire horizontal_tile_28_28_to_tile_28_27_3;

	wire horizontal_tile_29_27_to_tile_29_28_0;
	wire horizontal_tile_29_27_to_tile_29_28_1;
	wire horizontal_tile_29_27_to_tile_29_28_2;
	wire horizontal_tile_29_27_to_tile_29_28_3;
	wire horizontal_tile_29_28_to_tile_29_27_0;
	wire horizontal_tile_29_28_to_tile_29_27_1;
	wire horizontal_tile_29_28_to_tile_29_27_2;
	wire horizontal_tile_29_28_to_tile_29_27_3;

	wire horizontal_tile_30_27_to_tile_30_28_0;
	wire horizontal_tile_30_27_to_tile_30_28_1;
	wire horizontal_tile_30_27_to_tile_30_28_2;
	wire horizontal_tile_30_27_to_tile_30_28_3;
	wire horizontal_tile_30_28_to_tile_30_27_0;
	wire horizontal_tile_30_28_to_tile_30_27_1;
	wire horizontal_tile_30_28_to_tile_30_27_2;
	wire horizontal_tile_30_28_to_tile_30_27_3;

	wire horizontal_tile_31_27_to_tile_31_28_0;
	wire horizontal_tile_31_27_to_tile_31_28_1;
	wire horizontal_tile_31_27_to_tile_31_28_2;
	wire horizontal_tile_31_27_to_tile_31_28_3;
	wire horizontal_tile_31_28_to_tile_31_27_0;
	wire horizontal_tile_31_28_to_tile_31_27_1;
	wire horizontal_tile_31_28_to_tile_31_27_2;
	wire horizontal_tile_31_28_to_tile_31_27_3;

	wire horizontal_tile_0_28_to_tile_0_29_0;
	wire horizontal_tile_0_28_to_tile_0_29_1;
	wire horizontal_tile_0_28_to_tile_0_29_2;
	wire horizontal_tile_0_28_to_tile_0_29_3;
	wire horizontal_tile_0_29_to_tile_0_28_0;
	wire horizontal_tile_0_29_to_tile_0_28_1;
	wire horizontal_tile_0_29_to_tile_0_28_2;
	wire horizontal_tile_0_29_to_tile_0_28_3;

	wire horizontal_tile_1_28_to_tile_1_29_0;
	wire horizontal_tile_1_28_to_tile_1_29_1;
	wire horizontal_tile_1_28_to_tile_1_29_2;
	wire horizontal_tile_1_28_to_tile_1_29_3;
	wire horizontal_tile_1_29_to_tile_1_28_0;
	wire horizontal_tile_1_29_to_tile_1_28_1;
	wire horizontal_tile_1_29_to_tile_1_28_2;
	wire horizontal_tile_1_29_to_tile_1_28_3;

	wire horizontal_tile_2_28_to_tile_2_29_0;
	wire horizontal_tile_2_28_to_tile_2_29_1;
	wire horizontal_tile_2_28_to_tile_2_29_2;
	wire horizontal_tile_2_28_to_tile_2_29_3;
	wire horizontal_tile_2_29_to_tile_2_28_0;
	wire horizontal_tile_2_29_to_tile_2_28_1;
	wire horizontal_tile_2_29_to_tile_2_28_2;
	wire horizontal_tile_2_29_to_tile_2_28_3;

	wire horizontal_tile_3_28_to_tile_3_29_0;
	wire horizontal_tile_3_28_to_tile_3_29_1;
	wire horizontal_tile_3_28_to_tile_3_29_2;
	wire horizontal_tile_3_28_to_tile_3_29_3;
	wire horizontal_tile_3_29_to_tile_3_28_0;
	wire horizontal_tile_3_29_to_tile_3_28_1;
	wire horizontal_tile_3_29_to_tile_3_28_2;
	wire horizontal_tile_3_29_to_tile_3_28_3;

	wire horizontal_tile_4_28_to_tile_4_29_0;
	wire horizontal_tile_4_28_to_tile_4_29_1;
	wire horizontal_tile_4_28_to_tile_4_29_2;
	wire horizontal_tile_4_28_to_tile_4_29_3;
	wire horizontal_tile_4_29_to_tile_4_28_0;
	wire horizontal_tile_4_29_to_tile_4_28_1;
	wire horizontal_tile_4_29_to_tile_4_28_2;
	wire horizontal_tile_4_29_to_tile_4_28_3;

	wire horizontal_tile_5_28_to_tile_5_29_0;
	wire horizontal_tile_5_28_to_tile_5_29_1;
	wire horizontal_tile_5_28_to_tile_5_29_2;
	wire horizontal_tile_5_28_to_tile_5_29_3;
	wire horizontal_tile_5_29_to_tile_5_28_0;
	wire horizontal_tile_5_29_to_tile_5_28_1;
	wire horizontal_tile_5_29_to_tile_5_28_2;
	wire horizontal_tile_5_29_to_tile_5_28_3;

	wire horizontal_tile_6_28_to_tile_6_29_0;
	wire horizontal_tile_6_28_to_tile_6_29_1;
	wire horizontal_tile_6_28_to_tile_6_29_2;
	wire horizontal_tile_6_28_to_tile_6_29_3;
	wire horizontal_tile_6_29_to_tile_6_28_0;
	wire horizontal_tile_6_29_to_tile_6_28_1;
	wire horizontal_tile_6_29_to_tile_6_28_2;
	wire horizontal_tile_6_29_to_tile_6_28_3;

	wire horizontal_tile_7_28_to_tile_7_29_0;
	wire horizontal_tile_7_28_to_tile_7_29_1;
	wire horizontal_tile_7_28_to_tile_7_29_2;
	wire horizontal_tile_7_28_to_tile_7_29_3;
	wire horizontal_tile_7_29_to_tile_7_28_0;
	wire horizontal_tile_7_29_to_tile_7_28_1;
	wire horizontal_tile_7_29_to_tile_7_28_2;
	wire horizontal_tile_7_29_to_tile_7_28_3;

	wire horizontal_tile_8_28_to_tile_8_29_0;
	wire horizontal_tile_8_28_to_tile_8_29_1;
	wire horizontal_tile_8_28_to_tile_8_29_2;
	wire horizontal_tile_8_28_to_tile_8_29_3;
	wire horizontal_tile_8_29_to_tile_8_28_0;
	wire horizontal_tile_8_29_to_tile_8_28_1;
	wire horizontal_tile_8_29_to_tile_8_28_2;
	wire horizontal_tile_8_29_to_tile_8_28_3;

	wire horizontal_tile_9_28_to_tile_9_29_0;
	wire horizontal_tile_9_28_to_tile_9_29_1;
	wire horizontal_tile_9_28_to_tile_9_29_2;
	wire horizontal_tile_9_28_to_tile_9_29_3;
	wire horizontal_tile_9_29_to_tile_9_28_0;
	wire horizontal_tile_9_29_to_tile_9_28_1;
	wire horizontal_tile_9_29_to_tile_9_28_2;
	wire horizontal_tile_9_29_to_tile_9_28_3;

	wire horizontal_tile_10_28_to_tile_10_29_0;
	wire horizontal_tile_10_28_to_tile_10_29_1;
	wire horizontal_tile_10_28_to_tile_10_29_2;
	wire horizontal_tile_10_28_to_tile_10_29_3;
	wire horizontal_tile_10_29_to_tile_10_28_0;
	wire horizontal_tile_10_29_to_tile_10_28_1;
	wire horizontal_tile_10_29_to_tile_10_28_2;
	wire horizontal_tile_10_29_to_tile_10_28_3;

	wire horizontal_tile_11_28_to_tile_11_29_0;
	wire horizontal_tile_11_28_to_tile_11_29_1;
	wire horizontal_tile_11_28_to_tile_11_29_2;
	wire horizontal_tile_11_28_to_tile_11_29_3;
	wire horizontal_tile_11_29_to_tile_11_28_0;
	wire horizontal_tile_11_29_to_tile_11_28_1;
	wire horizontal_tile_11_29_to_tile_11_28_2;
	wire horizontal_tile_11_29_to_tile_11_28_3;

	wire horizontal_tile_12_28_to_tile_12_29_0;
	wire horizontal_tile_12_28_to_tile_12_29_1;
	wire horizontal_tile_12_28_to_tile_12_29_2;
	wire horizontal_tile_12_28_to_tile_12_29_3;
	wire horizontal_tile_12_29_to_tile_12_28_0;
	wire horizontal_tile_12_29_to_tile_12_28_1;
	wire horizontal_tile_12_29_to_tile_12_28_2;
	wire horizontal_tile_12_29_to_tile_12_28_3;

	wire horizontal_tile_13_28_to_tile_13_29_0;
	wire horizontal_tile_13_28_to_tile_13_29_1;
	wire horizontal_tile_13_28_to_tile_13_29_2;
	wire horizontal_tile_13_28_to_tile_13_29_3;
	wire horizontal_tile_13_29_to_tile_13_28_0;
	wire horizontal_tile_13_29_to_tile_13_28_1;
	wire horizontal_tile_13_29_to_tile_13_28_2;
	wire horizontal_tile_13_29_to_tile_13_28_3;

	wire horizontal_tile_14_28_to_tile_14_29_0;
	wire horizontal_tile_14_28_to_tile_14_29_1;
	wire horizontal_tile_14_28_to_tile_14_29_2;
	wire horizontal_tile_14_28_to_tile_14_29_3;
	wire horizontal_tile_14_29_to_tile_14_28_0;
	wire horizontal_tile_14_29_to_tile_14_28_1;
	wire horizontal_tile_14_29_to_tile_14_28_2;
	wire horizontal_tile_14_29_to_tile_14_28_3;

	wire horizontal_tile_15_28_to_tile_15_29_0;
	wire horizontal_tile_15_28_to_tile_15_29_1;
	wire horizontal_tile_15_28_to_tile_15_29_2;
	wire horizontal_tile_15_28_to_tile_15_29_3;
	wire horizontal_tile_15_29_to_tile_15_28_0;
	wire horizontal_tile_15_29_to_tile_15_28_1;
	wire horizontal_tile_15_29_to_tile_15_28_2;
	wire horizontal_tile_15_29_to_tile_15_28_3;

	wire horizontal_tile_16_28_to_tile_16_29_0;
	wire horizontal_tile_16_28_to_tile_16_29_1;
	wire horizontal_tile_16_28_to_tile_16_29_2;
	wire horizontal_tile_16_28_to_tile_16_29_3;
	wire horizontal_tile_16_29_to_tile_16_28_0;
	wire horizontal_tile_16_29_to_tile_16_28_1;
	wire horizontal_tile_16_29_to_tile_16_28_2;
	wire horizontal_tile_16_29_to_tile_16_28_3;

	wire horizontal_tile_17_28_to_tile_17_29_0;
	wire horizontal_tile_17_28_to_tile_17_29_1;
	wire horizontal_tile_17_28_to_tile_17_29_2;
	wire horizontal_tile_17_28_to_tile_17_29_3;
	wire horizontal_tile_17_29_to_tile_17_28_0;
	wire horizontal_tile_17_29_to_tile_17_28_1;
	wire horizontal_tile_17_29_to_tile_17_28_2;
	wire horizontal_tile_17_29_to_tile_17_28_3;

	wire horizontal_tile_18_28_to_tile_18_29_0;
	wire horizontal_tile_18_28_to_tile_18_29_1;
	wire horizontal_tile_18_28_to_tile_18_29_2;
	wire horizontal_tile_18_28_to_tile_18_29_3;
	wire horizontal_tile_18_29_to_tile_18_28_0;
	wire horizontal_tile_18_29_to_tile_18_28_1;
	wire horizontal_tile_18_29_to_tile_18_28_2;
	wire horizontal_tile_18_29_to_tile_18_28_3;

	wire horizontal_tile_19_28_to_tile_19_29_0;
	wire horizontal_tile_19_28_to_tile_19_29_1;
	wire horizontal_tile_19_28_to_tile_19_29_2;
	wire horizontal_tile_19_28_to_tile_19_29_3;
	wire horizontal_tile_19_29_to_tile_19_28_0;
	wire horizontal_tile_19_29_to_tile_19_28_1;
	wire horizontal_tile_19_29_to_tile_19_28_2;
	wire horizontal_tile_19_29_to_tile_19_28_3;

	wire horizontal_tile_20_28_to_tile_20_29_0;
	wire horizontal_tile_20_28_to_tile_20_29_1;
	wire horizontal_tile_20_28_to_tile_20_29_2;
	wire horizontal_tile_20_28_to_tile_20_29_3;
	wire horizontal_tile_20_29_to_tile_20_28_0;
	wire horizontal_tile_20_29_to_tile_20_28_1;
	wire horizontal_tile_20_29_to_tile_20_28_2;
	wire horizontal_tile_20_29_to_tile_20_28_3;

	wire horizontal_tile_21_28_to_tile_21_29_0;
	wire horizontal_tile_21_28_to_tile_21_29_1;
	wire horizontal_tile_21_28_to_tile_21_29_2;
	wire horizontal_tile_21_28_to_tile_21_29_3;
	wire horizontal_tile_21_29_to_tile_21_28_0;
	wire horizontal_tile_21_29_to_tile_21_28_1;
	wire horizontal_tile_21_29_to_tile_21_28_2;
	wire horizontal_tile_21_29_to_tile_21_28_3;

	wire horizontal_tile_22_28_to_tile_22_29_0;
	wire horizontal_tile_22_28_to_tile_22_29_1;
	wire horizontal_tile_22_28_to_tile_22_29_2;
	wire horizontal_tile_22_28_to_tile_22_29_3;
	wire horizontal_tile_22_29_to_tile_22_28_0;
	wire horizontal_tile_22_29_to_tile_22_28_1;
	wire horizontal_tile_22_29_to_tile_22_28_2;
	wire horizontal_tile_22_29_to_tile_22_28_3;

	wire horizontal_tile_23_28_to_tile_23_29_0;
	wire horizontal_tile_23_28_to_tile_23_29_1;
	wire horizontal_tile_23_28_to_tile_23_29_2;
	wire horizontal_tile_23_28_to_tile_23_29_3;
	wire horizontal_tile_23_29_to_tile_23_28_0;
	wire horizontal_tile_23_29_to_tile_23_28_1;
	wire horizontal_tile_23_29_to_tile_23_28_2;
	wire horizontal_tile_23_29_to_tile_23_28_3;

	wire horizontal_tile_24_28_to_tile_24_29_0;
	wire horizontal_tile_24_28_to_tile_24_29_1;
	wire horizontal_tile_24_28_to_tile_24_29_2;
	wire horizontal_tile_24_28_to_tile_24_29_3;
	wire horizontal_tile_24_29_to_tile_24_28_0;
	wire horizontal_tile_24_29_to_tile_24_28_1;
	wire horizontal_tile_24_29_to_tile_24_28_2;
	wire horizontal_tile_24_29_to_tile_24_28_3;

	wire horizontal_tile_25_28_to_tile_25_29_0;
	wire horizontal_tile_25_28_to_tile_25_29_1;
	wire horizontal_tile_25_28_to_tile_25_29_2;
	wire horizontal_tile_25_28_to_tile_25_29_3;
	wire horizontal_tile_25_29_to_tile_25_28_0;
	wire horizontal_tile_25_29_to_tile_25_28_1;
	wire horizontal_tile_25_29_to_tile_25_28_2;
	wire horizontal_tile_25_29_to_tile_25_28_3;

	wire horizontal_tile_26_28_to_tile_26_29_0;
	wire horizontal_tile_26_28_to_tile_26_29_1;
	wire horizontal_tile_26_28_to_tile_26_29_2;
	wire horizontal_tile_26_28_to_tile_26_29_3;
	wire horizontal_tile_26_29_to_tile_26_28_0;
	wire horizontal_tile_26_29_to_tile_26_28_1;
	wire horizontal_tile_26_29_to_tile_26_28_2;
	wire horizontal_tile_26_29_to_tile_26_28_3;

	wire horizontal_tile_27_28_to_tile_27_29_0;
	wire horizontal_tile_27_28_to_tile_27_29_1;
	wire horizontal_tile_27_28_to_tile_27_29_2;
	wire horizontal_tile_27_28_to_tile_27_29_3;
	wire horizontal_tile_27_29_to_tile_27_28_0;
	wire horizontal_tile_27_29_to_tile_27_28_1;
	wire horizontal_tile_27_29_to_tile_27_28_2;
	wire horizontal_tile_27_29_to_tile_27_28_3;

	wire horizontal_tile_28_28_to_tile_28_29_0;
	wire horizontal_tile_28_28_to_tile_28_29_1;
	wire horizontal_tile_28_28_to_tile_28_29_2;
	wire horizontal_tile_28_28_to_tile_28_29_3;
	wire horizontal_tile_28_29_to_tile_28_28_0;
	wire horizontal_tile_28_29_to_tile_28_28_1;
	wire horizontal_tile_28_29_to_tile_28_28_2;
	wire horizontal_tile_28_29_to_tile_28_28_3;

	wire horizontal_tile_29_28_to_tile_29_29_0;
	wire horizontal_tile_29_28_to_tile_29_29_1;
	wire horizontal_tile_29_28_to_tile_29_29_2;
	wire horizontal_tile_29_28_to_tile_29_29_3;
	wire horizontal_tile_29_29_to_tile_29_28_0;
	wire horizontal_tile_29_29_to_tile_29_28_1;
	wire horizontal_tile_29_29_to_tile_29_28_2;
	wire horizontal_tile_29_29_to_tile_29_28_3;

	wire horizontal_tile_30_28_to_tile_30_29_0;
	wire horizontal_tile_30_28_to_tile_30_29_1;
	wire horizontal_tile_30_28_to_tile_30_29_2;
	wire horizontal_tile_30_28_to_tile_30_29_3;
	wire horizontal_tile_30_29_to_tile_30_28_0;
	wire horizontal_tile_30_29_to_tile_30_28_1;
	wire horizontal_tile_30_29_to_tile_30_28_2;
	wire horizontal_tile_30_29_to_tile_30_28_3;

	wire horizontal_tile_31_28_to_tile_31_29_0;
	wire horizontal_tile_31_28_to_tile_31_29_1;
	wire horizontal_tile_31_28_to_tile_31_29_2;
	wire horizontal_tile_31_28_to_tile_31_29_3;
	wire horizontal_tile_31_29_to_tile_31_28_0;
	wire horizontal_tile_31_29_to_tile_31_28_1;
	wire horizontal_tile_31_29_to_tile_31_28_2;
	wire horizontal_tile_31_29_to_tile_31_28_3;

	wire horizontal_tile_0_29_to_tile_0_30_0;
	wire horizontal_tile_0_29_to_tile_0_30_1;
	wire horizontal_tile_0_29_to_tile_0_30_2;
	wire horizontal_tile_0_29_to_tile_0_30_3;
	wire horizontal_tile_0_30_to_tile_0_29_0;
	wire horizontal_tile_0_30_to_tile_0_29_1;
	wire horizontal_tile_0_30_to_tile_0_29_2;
	wire horizontal_tile_0_30_to_tile_0_29_3;

	wire horizontal_tile_1_29_to_tile_1_30_0;
	wire horizontal_tile_1_29_to_tile_1_30_1;
	wire horizontal_tile_1_29_to_tile_1_30_2;
	wire horizontal_tile_1_29_to_tile_1_30_3;
	wire horizontal_tile_1_30_to_tile_1_29_0;
	wire horizontal_tile_1_30_to_tile_1_29_1;
	wire horizontal_tile_1_30_to_tile_1_29_2;
	wire horizontal_tile_1_30_to_tile_1_29_3;

	wire horizontal_tile_2_29_to_tile_2_30_0;
	wire horizontal_tile_2_29_to_tile_2_30_1;
	wire horizontal_tile_2_29_to_tile_2_30_2;
	wire horizontal_tile_2_29_to_tile_2_30_3;
	wire horizontal_tile_2_30_to_tile_2_29_0;
	wire horizontal_tile_2_30_to_tile_2_29_1;
	wire horizontal_tile_2_30_to_tile_2_29_2;
	wire horizontal_tile_2_30_to_tile_2_29_3;

	wire horizontal_tile_3_29_to_tile_3_30_0;
	wire horizontal_tile_3_29_to_tile_3_30_1;
	wire horizontal_tile_3_29_to_tile_3_30_2;
	wire horizontal_tile_3_29_to_tile_3_30_3;
	wire horizontal_tile_3_30_to_tile_3_29_0;
	wire horizontal_tile_3_30_to_tile_3_29_1;
	wire horizontal_tile_3_30_to_tile_3_29_2;
	wire horizontal_tile_3_30_to_tile_3_29_3;

	wire horizontal_tile_4_29_to_tile_4_30_0;
	wire horizontal_tile_4_29_to_tile_4_30_1;
	wire horizontal_tile_4_29_to_tile_4_30_2;
	wire horizontal_tile_4_29_to_tile_4_30_3;
	wire horizontal_tile_4_30_to_tile_4_29_0;
	wire horizontal_tile_4_30_to_tile_4_29_1;
	wire horizontal_tile_4_30_to_tile_4_29_2;
	wire horizontal_tile_4_30_to_tile_4_29_3;

	wire horizontal_tile_5_29_to_tile_5_30_0;
	wire horizontal_tile_5_29_to_tile_5_30_1;
	wire horizontal_tile_5_29_to_tile_5_30_2;
	wire horizontal_tile_5_29_to_tile_5_30_3;
	wire horizontal_tile_5_30_to_tile_5_29_0;
	wire horizontal_tile_5_30_to_tile_5_29_1;
	wire horizontal_tile_5_30_to_tile_5_29_2;
	wire horizontal_tile_5_30_to_tile_5_29_3;

	wire horizontal_tile_6_29_to_tile_6_30_0;
	wire horizontal_tile_6_29_to_tile_6_30_1;
	wire horizontal_tile_6_29_to_tile_6_30_2;
	wire horizontal_tile_6_29_to_tile_6_30_3;
	wire horizontal_tile_6_30_to_tile_6_29_0;
	wire horizontal_tile_6_30_to_tile_6_29_1;
	wire horizontal_tile_6_30_to_tile_6_29_2;
	wire horizontal_tile_6_30_to_tile_6_29_3;

	wire horizontal_tile_7_29_to_tile_7_30_0;
	wire horizontal_tile_7_29_to_tile_7_30_1;
	wire horizontal_tile_7_29_to_tile_7_30_2;
	wire horizontal_tile_7_29_to_tile_7_30_3;
	wire horizontal_tile_7_30_to_tile_7_29_0;
	wire horizontal_tile_7_30_to_tile_7_29_1;
	wire horizontal_tile_7_30_to_tile_7_29_2;
	wire horizontal_tile_7_30_to_tile_7_29_3;

	wire horizontal_tile_8_29_to_tile_8_30_0;
	wire horizontal_tile_8_29_to_tile_8_30_1;
	wire horizontal_tile_8_29_to_tile_8_30_2;
	wire horizontal_tile_8_29_to_tile_8_30_3;
	wire horizontal_tile_8_30_to_tile_8_29_0;
	wire horizontal_tile_8_30_to_tile_8_29_1;
	wire horizontal_tile_8_30_to_tile_8_29_2;
	wire horizontal_tile_8_30_to_tile_8_29_3;

	wire horizontal_tile_9_29_to_tile_9_30_0;
	wire horizontal_tile_9_29_to_tile_9_30_1;
	wire horizontal_tile_9_29_to_tile_9_30_2;
	wire horizontal_tile_9_29_to_tile_9_30_3;
	wire horizontal_tile_9_30_to_tile_9_29_0;
	wire horizontal_tile_9_30_to_tile_9_29_1;
	wire horizontal_tile_9_30_to_tile_9_29_2;
	wire horizontal_tile_9_30_to_tile_9_29_3;

	wire horizontal_tile_10_29_to_tile_10_30_0;
	wire horizontal_tile_10_29_to_tile_10_30_1;
	wire horizontal_tile_10_29_to_tile_10_30_2;
	wire horizontal_tile_10_29_to_tile_10_30_3;
	wire horizontal_tile_10_30_to_tile_10_29_0;
	wire horizontal_tile_10_30_to_tile_10_29_1;
	wire horizontal_tile_10_30_to_tile_10_29_2;
	wire horizontal_tile_10_30_to_tile_10_29_3;

	wire horizontal_tile_11_29_to_tile_11_30_0;
	wire horizontal_tile_11_29_to_tile_11_30_1;
	wire horizontal_tile_11_29_to_tile_11_30_2;
	wire horizontal_tile_11_29_to_tile_11_30_3;
	wire horizontal_tile_11_30_to_tile_11_29_0;
	wire horizontal_tile_11_30_to_tile_11_29_1;
	wire horizontal_tile_11_30_to_tile_11_29_2;
	wire horizontal_tile_11_30_to_tile_11_29_3;

	wire horizontal_tile_12_29_to_tile_12_30_0;
	wire horizontal_tile_12_29_to_tile_12_30_1;
	wire horizontal_tile_12_29_to_tile_12_30_2;
	wire horizontal_tile_12_29_to_tile_12_30_3;
	wire horizontal_tile_12_30_to_tile_12_29_0;
	wire horizontal_tile_12_30_to_tile_12_29_1;
	wire horizontal_tile_12_30_to_tile_12_29_2;
	wire horizontal_tile_12_30_to_tile_12_29_3;

	wire horizontal_tile_13_29_to_tile_13_30_0;
	wire horizontal_tile_13_29_to_tile_13_30_1;
	wire horizontal_tile_13_29_to_tile_13_30_2;
	wire horizontal_tile_13_29_to_tile_13_30_3;
	wire horizontal_tile_13_30_to_tile_13_29_0;
	wire horizontal_tile_13_30_to_tile_13_29_1;
	wire horizontal_tile_13_30_to_tile_13_29_2;
	wire horizontal_tile_13_30_to_tile_13_29_3;

	wire horizontal_tile_14_29_to_tile_14_30_0;
	wire horizontal_tile_14_29_to_tile_14_30_1;
	wire horizontal_tile_14_29_to_tile_14_30_2;
	wire horizontal_tile_14_29_to_tile_14_30_3;
	wire horizontal_tile_14_30_to_tile_14_29_0;
	wire horizontal_tile_14_30_to_tile_14_29_1;
	wire horizontal_tile_14_30_to_tile_14_29_2;
	wire horizontal_tile_14_30_to_tile_14_29_3;

	wire horizontal_tile_15_29_to_tile_15_30_0;
	wire horizontal_tile_15_29_to_tile_15_30_1;
	wire horizontal_tile_15_29_to_tile_15_30_2;
	wire horizontal_tile_15_29_to_tile_15_30_3;
	wire horizontal_tile_15_30_to_tile_15_29_0;
	wire horizontal_tile_15_30_to_tile_15_29_1;
	wire horizontal_tile_15_30_to_tile_15_29_2;
	wire horizontal_tile_15_30_to_tile_15_29_3;

	wire horizontal_tile_16_29_to_tile_16_30_0;
	wire horizontal_tile_16_29_to_tile_16_30_1;
	wire horizontal_tile_16_29_to_tile_16_30_2;
	wire horizontal_tile_16_29_to_tile_16_30_3;
	wire horizontal_tile_16_30_to_tile_16_29_0;
	wire horizontal_tile_16_30_to_tile_16_29_1;
	wire horizontal_tile_16_30_to_tile_16_29_2;
	wire horizontal_tile_16_30_to_tile_16_29_3;

	wire horizontal_tile_17_29_to_tile_17_30_0;
	wire horizontal_tile_17_29_to_tile_17_30_1;
	wire horizontal_tile_17_29_to_tile_17_30_2;
	wire horizontal_tile_17_29_to_tile_17_30_3;
	wire horizontal_tile_17_30_to_tile_17_29_0;
	wire horizontal_tile_17_30_to_tile_17_29_1;
	wire horizontal_tile_17_30_to_tile_17_29_2;
	wire horizontal_tile_17_30_to_tile_17_29_3;

	wire horizontal_tile_18_29_to_tile_18_30_0;
	wire horizontal_tile_18_29_to_tile_18_30_1;
	wire horizontal_tile_18_29_to_tile_18_30_2;
	wire horizontal_tile_18_29_to_tile_18_30_3;
	wire horizontal_tile_18_30_to_tile_18_29_0;
	wire horizontal_tile_18_30_to_tile_18_29_1;
	wire horizontal_tile_18_30_to_tile_18_29_2;
	wire horizontal_tile_18_30_to_tile_18_29_3;

	wire horizontal_tile_19_29_to_tile_19_30_0;
	wire horizontal_tile_19_29_to_tile_19_30_1;
	wire horizontal_tile_19_29_to_tile_19_30_2;
	wire horizontal_tile_19_29_to_tile_19_30_3;
	wire horizontal_tile_19_30_to_tile_19_29_0;
	wire horizontal_tile_19_30_to_tile_19_29_1;
	wire horizontal_tile_19_30_to_tile_19_29_2;
	wire horizontal_tile_19_30_to_tile_19_29_3;

	wire horizontal_tile_20_29_to_tile_20_30_0;
	wire horizontal_tile_20_29_to_tile_20_30_1;
	wire horizontal_tile_20_29_to_tile_20_30_2;
	wire horizontal_tile_20_29_to_tile_20_30_3;
	wire horizontal_tile_20_30_to_tile_20_29_0;
	wire horizontal_tile_20_30_to_tile_20_29_1;
	wire horizontal_tile_20_30_to_tile_20_29_2;
	wire horizontal_tile_20_30_to_tile_20_29_3;

	wire horizontal_tile_21_29_to_tile_21_30_0;
	wire horizontal_tile_21_29_to_tile_21_30_1;
	wire horizontal_tile_21_29_to_tile_21_30_2;
	wire horizontal_tile_21_29_to_tile_21_30_3;
	wire horizontal_tile_21_30_to_tile_21_29_0;
	wire horizontal_tile_21_30_to_tile_21_29_1;
	wire horizontal_tile_21_30_to_tile_21_29_2;
	wire horizontal_tile_21_30_to_tile_21_29_3;

	wire horizontal_tile_22_29_to_tile_22_30_0;
	wire horizontal_tile_22_29_to_tile_22_30_1;
	wire horizontal_tile_22_29_to_tile_22_30_2;
	wire horizontal_tile_22_29_to_tile_22_30_3;
	wire horizontal_tile_22_30_to_tile_22_29_0;
	wire horizontal_tile_22_30_to_tile_22_29_1;
	wire horizontal_tile_22_30_to_tile_22_29_2;
	wire horizontal_tile_22_30_to_tile_22_29_3;

	wire horizontal_tile_23_29_to_tile_23_30_0;
	wire horizontal_tile_23_29_to_tile_23_30_1;
	wire horizontal_tile_23_29_to_tile_23_30_2;
	wire horizontal_tile_23_29_to_tile_23_30_3;
	wire horizontal_tile_23_30_to_tile_23_29_0;
	wire horizontal_tile_23_30_to_tile_23_29_1;
	wire horizontal_tile_23_30_to_tile_23_29_2;
	wire horizontal_tile_23_30_to_tile_23_29_3;

	wire horizontal_tile_24_29_to_tile_24_30_0;
	wire horizontal_tile_24_29_to_tile_24_30_1;
	wire horizontal_tile_24_29_to_tile_24_30_2;
	wire horizontal_tile_24_29_to_tile_24_30_3;
	wire horizontal_tile_24_30_to_tile_24_29_0;
	wire horizontal_tile_24_30_to_tile_24_29_1;
	wire horizontal_tile_24_30_to_tile_24_29_2;
	wire horizontal_tile_24_30_to_tile_24_29_3;

	wire horizontal_tile_25_29_to_tile_25_30_0;
	wire horizontal_tile_25_29_to_tile_25_30_1;
	wire horizontal_tile_25_29_to_tile_25_30_2;
	wire horizontal_tile_25_29_to_tile_25_30_3;
	wire horizontal_tile_25_30_to_tile_25_29_0;
	wire horizontal_tile_25_30_to_tile_25_29_1;
	wire horizontal_tile_25_30_to_tile_25_29_2;
	wire horizontal_tile_25_30_to_tile_25_29_3;

	wire horizontal_tile_26_29_to_tile_26_30_0;
	wire horizontal_tile_26_29_to_tile_26_30_1;
	wire horizontal_tile_26_29_to_tile_26_30_2;
	wire horizontal_tile_26_29_to_tile_26_30_3;
	wire horizontal_tile_26_30_to_tile_26_29_0;
	wire horizontal_tile_26_30_to_tile_26_29_1;
	wire horizontal_tile_26_30_to_tile_26_29_2;
	wire horizontal_tile_26_30_to_tile_26_29_3;

	wire horizontal_tile_27_29_to_tile_27_30_0;
	wire horizontal_tile_27_29_to_tile_27_30_1;
	wire horizontal_tile_27_29_to_tile_27_30_2;
	wire horizontal_tile_27_29_to_tile_27_30_3;
	wire horizontal_tile_27_30_to_tile_27_29_0;
	wire horizontal_tile_27_30_to_tile_27_29_1;
	wire horizontal_tile_27_30_to_tile_27_29_2;
	wire horizontal_tile_27_30_to_tile_27_29_3;

	wire horizontal_tile_28_29_to_tile_28_30_0;
	wire horizontal_tile_28_29_to_tile_28_30_1;
	wire horizontal_tile_28_29_to_tile_28_30_2;
	wire horizontal_tile_28_29_to_tile_28_30_3;
	wire horizontal_tile_28_30_to_tile_28_29_0;
	wire horizontal_tile_28_30_to_tile_28_29_1;
	wire horizontal_tile_28_30_to_tile_28_29_2;
	wire horizontal_tile_28_30_to_tile_28_29_3;

	wire horizontal_tile_29_29_to_tile_29_30_0;
	wire horizontal_tile_29_29_to_tile_29_30_1;
	wire horizontal_tile_29_29_to_tile_29_30_2;
	wire horizontal_tile_29_29_to_tile_29_30_3;
	wire horizontal_tile_29_30_to_tile_29_29_0;
	wire horizontal_tile_29_30_to_tile_29_29_1;
	wire horizontal_tile_29_30_to_tile_29_29_2;
	wire horizontal_tile_29_30_to_tile_29_29_3;

	wire horizontal_tile_30_29_to_tile_30_30_0;
	wire horizontal_tile_30_29_to_tile_30_30_1;
	wire horizontal_tile_30_29_to_tile_30_30_2;
	wire horizontal_tile_30_29_to_tile_30_30_3;
	wire horizontal_tile_30_30_to_tile_30_29_0;
	wire horizontal_tile_30_30_to_tile_30_29_1;
	wire horizontal_tile_30_30_to_tile_30_29_2;
	wire horizontal_tile_30_30_to_tile_30_29_3;

	wire horizontal_tile_31_29_to_tile_31_30_0;
	wire horizontal_tile_31_29_to_tile_31_30_1;
	wire horizontal_tile_31_29_to_tile_31_30_2;
	wire horizontal_tile_31_29_to_tile_31_30_3;
	wire horizontal_tile_31_30_to_tile_31_29_0;
	wire horizontal_tile_31_30_to_tile_31_29_1;
	wire horizontal_tile_31_30_to_tile_31_29_2;
	wire horizontal_tile_31_30_to_tile_31_29_3;

	wire horizontal_tile_0_30_to_tile_0_31_0;
	wire horizontal_tile_0_30_to_tile_0_31_1;
	wire horizontal_tile_0_30_to_tile_0_31_2;
	wire horizontal_tile_0_30_to_tile_0_31_3;
	wire horizontal_tile_0_31_to_tile_0_30_0;
	wire horizontal_tile_0_31_to_tile_0_30_1;
	wire horizontal_tile_0_31_to_tile_0_30_2;
	wire horizontal_tile_0_31_to_tile_0_30_3;

	wire horizontal_tile_1_30_to_tile_1_31_0;
	wire horizontal_tile_1_30_to_tile_1_31_1;
	wire horizontal_tile_1_30_to_tile_1_31_2;
	wire horizontal_tile_1_30_to_tile_1_31_3;
	wire horizontal_tile_1_31_to_tile_1_30_0;
	wire horizontal_tile_1_31_to_tile_1_30_1;
	wire horizontal_tile_1_31_to_tile_1_30_2;
	wire horizontal_tile_1_31_to_tile_1_30_3;

	wire horizontal_tile_2_30_to_tile_2_31_0;
	wire horizontal_tile_2_30_to_tile_2_31_1;
	wire horizontal_tile_2_30_to_tile_2_31_2;
	wire horizontal_tile_2_30_to_tile_2_31_3;
	wire horizontal_tile_2_31_to_tile_2_30_0;
	wire horizontal_tile_2_31_to_tile_2_30_1;
	wire horizontal_tile_2_31_to_tile_2_30_2;
	wire horizontal_tile_2_31_to_tile_2_30_3;

	wire horizontal_tile_3_30_to_tile_3_31_0;
	wire horizontal_tile_3_30_to_tile_3_31_1;
	wire horizontal_tile_3_30_to_tile_3_31_2;
	wire horizontal_tile_3_30_to_tile_3_31_3;
	wire horizontal_tile_3_31_to_tile_3_30_0;
	wire horizontal_tile_3_31_to_tile_3_30_1;
	wire horizontal_tile_3_31_to_tile_3_30_2;
	wire horizontal_tile_3_31_to_tile_3_30_3;

	wire horizontal_tile_4_30_to_tile_4_31_0;
	wire horizontal_tile_4_30_to_tile_4_31_1;
	wire horizontal_tile_4_30_to_tile_4_31_2;
	wire horizontal_tile_4_30_to_tile_4_31_3;
	wire horizontal_tile_4_31_to_tile_4_30_0;
	wire horizontal_tile_4_31_to_tile_4_30_1;
	wire horizontal_tile_4_31_to_tile_4_30_2;
	wire horizontal_tile_4_31_to_tile_4_30_3;

	wire horizontal_tile_5_30_to_tile_5_31_0;
	wire horizontal_tile_5_30_to_tile_5_31_1;
	wire horizontal_tile_5_30_to_tile_5_31_2;
	wire horizontal_tile_5_30_to_tile_5_31_3;
	wire horizontal_tile_5_31_to_tile_5_30_0;
	wire horizontal_tile_5_31_to_tile_5_30_1;
	wire horizontal_tile_5_31_to_tile_5_30_2;
	wire horizontal_tile_5_31_to_tile_5_30_3;

	wire horizontal_tile_6_30_to_tile_6_31_0;
	wire horizontal_tile_6_30_to_tile_6_31_1;
	wire horizontal_tile_6_30_to_tile_6_31_2;
	wire horizontal_tile_6_30_to_tile_6_31_3;
	wire horizontal_tile_6_31_to_tile_6_30_0;
	wire horizontal_tile_6_31_to_tile_6_30_1;
	wire horizontal_tile_6_31_to_tile_6_30_2;
	wire horizontal_tile_6_31_to_tile_6_30_3;

	wire horizontal_tile_7_30_to_tile_7_31_0;
	wire horizontal_tile_7_30_to_tile_7_31_1;
	wire horizontal_tile_7_30_to_tile_7_31_2;
	wire horizontal_tile_7_30_to_tile_7_31_3;
	wire horizontal_tile_7_31_to_tile_7_30_0;
	wire horizontal_tile_7_31_to_tile_7_30_1;
	wire horizontal_tile_7_31_to_tile_7_30_2;
	wire horizontal_tile_7_31_to_tile_7_30_3;

	wire horizontal_tile_8_30_to_tile_8_31_0;
	wire horizontal_tile_8_30_to_tile_8_31_1;
	wire horizontal_tile_8_30_to_tile_8_31_2;
	wire horizontal_tile_8_30_to_tile_8_31_3;
	wire horizontal_tile_8_31_to_tile_8_30_0;
	wire horizontal_tile_8_31_to_tile_8_30_1;
	wire horizontal_tile_8_31_to_tile_8_30_2;
	wire horizontal_tile_8_31_to_tile_8_30_3;

	wire horizontal_tile_9_30_to_tile_9_31_0;
	wire horizontal_tile_9_30_to_tile_9_31_1;
	wire horizontal_tile_9_30_to_tile_9_31_2;
	wire horizontal_tile_9_30_to_tile_9_31_3;
	wire horizontal_tile_9_31_to_tile_9_30_0;
	wire horizontal_tile_9_31_to_tile_9_30_1;
	wire horizontal_tile_9_31_to_tile_9_30_2;
	wire horizontal_tile_9_31_to_tile_9_30_3;

	wire horizontal_tile_10_30_to_tile_10_31_0;
	wire horizontal_tile_10_30_to_tile_10_31_1;
	wire horizontal_tile_10_30_to_tile_10_31_2;
	wire horizontal_tile_10_30_to_tile_10_31_3;
	wire horizontal_tile_10_31_to_tile_10_30_0;
	wire horizontal_tile_10_31_to_tile_10_30_1;
	wire horizontal_tile_10_31_to_tile_10_30_2;
	wire horizontal_tile_10_31_to_tile_10_30_3;

	wire horizontal_tile_11_30_to_tile_11_31_0;
	wire horizontal_tile_11_30_to_tile_11_31_1;
	wire horizontal_tile_11_30_to_tile_11_31_2;
	wire horizontal_tile_11_30_to_tile_11_31_3;
	wire horizontal_tile_11_31_to_tile_11_30_0;
	wire horizontal_tile_11_31_to_tile_11_30_1;
	wire horizontal_tile_11_31_to_tile_11_30_2;
	wire horizontal_tile_11_31_to_tile_11_30_3;

	wire horizontal_tile_12_30_to_tile_12_31_0;
	wire horizontal_tile_12_30_to_tile_12_31_1;
	wire horizontal_tile_12_30_to_tile_12_31_2;
	wire horizontal_tile_12_30_to_tile_12_31_3;
	wire horizontal_tile_12_31_to_tile_12_30_0;
	wire horizontal_tile_12_31_to_tile_12_30_1;
	wire horizontal_tile_12_31_to_tile_12_30_2;
	wire horizontal_tile_12_31_to_tile_12_30_3;

	wire horizontal_tile_13_30_to_tile_13_31_0;
	wire horizontal_tile_13_30_to_tile_13_31_1;
	wire horizontal_tile_13_30_to_tile_13_31_2;
	wire horizontal_tile_13_30_to_tile_13_31_3;
	wire horizontal_tile_13_31_to_tile_13_30_0;
	wire horizontal_tile_13_31_to_tile_13_30_1;
	wire horizontal_tile_13_31_to_tile_13_30_2;
	wire horizontal_tile_13_31_to_tile_13_30_3;

	wire horizontal_tile_14_30_to_tile_14_31_0;
	wire horizontal_tile_14_30_to_tile_14_31_1;
	wire horizontal_tile_14_30_to_tile_14_31_2;
	wire horizontal_tile_14_30_to_tile_14_31_3;
	wire horizontal_tile_14_31_to_tile_14_30_0;
	wire horizontal_tile_14_31_to_tile_14_30_1;
	wire horizontal_tile_14_31_to_tile_14_30_2;
	wire horizontal_tile_14_31_to_tile_14_30_3;

	wire horizontal_tile_15_30_to_tile_15_31_0;
	wire horizontal_tile_15_30_to_tile_15_31_1;
	wire horizontal_tile_15_30_to_tile_15_31_2;
	wire horizontal_tile_15_30_to_tile_15_31_3;
	wire horizontal_tile_15_31_to_tile_15_30_0;
	wire horizontal_tile_15_31_to_tile_15_30_1;
	wire horizontal_tile_15_31_to_tile_15_30_2;
	wire horizontal_tile_15_31_to_tile_15_30_3;

	wire horizontal_tile_16_30_to_tile_16_31_0;
	wire horizontal_tile_16_30_to_tile_16_31_1;
	wire horizontal_tile_16_30_to_tile_16_31_2;
	wire horizontal_tile_16_30_to_tile_16_31_3;
	wire horizontal_tile_16_31_to_tile_16_30_0;
	wire horizontal_tile_16_31_to_tile_16_30_1;
	wire horizontal_tile_16_31_to_tile_16_30_2;
	wire horizontal_tile_16_31_to_tile_16_30_3;

	wire horizontal_tile_17_30_to_tile_17_31_0;
	wire horizontal_tile_17_30_to_tile_17_31_1;
	wire horizontal_tile_17_30_to_tile_17_31_2;
	wire horizontal_tile_17_30_to_tile_17_31_3;
	wire horizontal_tile_17_31_to_tile_17_30_0;
	wire horizontal_tile_17_31_to_tile_17_30_1;
	wire horizontal_tile_17_31_to_tile_17_30_2;
	wire horizontal_tile_17_31_to_tile_17_30_3;

	wire horizontal_tile_18_30_to_tile_18_31_0;
	wire horizontal_tile_18_30_to_tile_18_31_1;
	wire horizontal_tile_18_30_to_tile_18_31_2;
	wire horizontal_tile_18_30_to_tile_18_31_3;
	wire horizontal_tile_18_31_to_tile_18_30_0;
	wire horizontal_tile_18_31_to_tile_18_30_1;
	wire horizontal_tile_18_31_to_tile_18_30_2;
	wire horizontal_tile_18_31_to_tile_18_30_3;

	wire horizontal_tile_19_30_to_tile_19_31_0;
	wire horizontal_tile_19_30_to_tile_19_31_1;
	wire horizontal_tile_19_30_to_tile_19_31_2;
	wire horizontal_tile_19_30_to_tile_19_31_3;
	wire horizontal_tile_19_31_to_tile_19_30_0;
	wire horizontal_tile_19_31_to_tile_19_30_1;
	wire horizontal_tile_19_31_to_tile_19_30_2;
	wire horizontal_tile_19_31_to_tile_19_30_3;

	wire horizontal_tile_20_30_to_tile_20_31_0;
	wire horizontal_tile_20_30_to_tile_20_31_1;
	wire horizontal_tile_20_30_to_tile_20_31_2;
	wire horizontal_tile_20_30_to_tile_20_31_3;
	wire horizontal_tile_20_31_to_tile_20_30_0;
	wire horizontal_tile_20_31_to_tile_20_30_1;
	wire horizontal_tile_20_31_to_tile_20_30_2;
	wire horizontal_tile_20_31_to_tile_20_30_3;

	wire horizontal_tile_21_30_to_tile_21_31_0;
	wire horizontal_tile_21_30_to_tile_21_31_1;
	wire horizontal_tile_21_30_to_tile_21_31_2;
	wire horizontal_tile_21_30_to_tile_21_31_3;
	wire horizontal_tile_21_31_to_tile_21_30_0;
	wire horizontal_tile_21_31_to_tile_21_30_1;
	wire horizontal_tile_21_31_to_tile_21_30_2;
	wire horizontal_tile_21_31_to_tile_21_30_3;

	wire horizontal_tile_22_30_to_tile_22_31_0;
	wire horizontal_tile_22_30_to_tile_22_31_1;
	wire horizontal_tile_22_30_to_tile_22_31_2;
	wire horizontal_tile_22_30_to_tile_22_31_3;
	wire horizontal_tile_22_31_to_tile_22_30_0;
	wire horizontal_tile_22_31_to_tile_22_30_1;
	wire horizontal_tile_22_31_to_tile_22_30_2;
	wire horizontal_tile_22_31_to_tile_22_30_3;

	wire horizontal_tile_23_30_to_tile_23_31_0;
	wire horizontal_tile_23_30_to_tile_23_31_1;
	wire horizontal_tile_23_30_to_tile_23_31_2;
	wire horizontal_tile_23_30_to_tile_23_31_3;
	wire horizontal_tile_23_31_to_tile_23_30_0;
	wire horizontal_tile_23_31_to_tile_23_30_1;
	wire horizontal_tile_23_31_to_tile_23_30_2;
	wire horizontal_tile_23_31_to_tile_23_30_3;

	wire horizontal_tile_24_30_to_tile_24_31_0;
	wire horizontal_tile_24_30_to_tile_24_31_1;
	wire horizontal_tile_24_30_to_tile_24_31_2;
	wire horizontal_tile_24_30_to_tile_24_31_3;
	wire horizontal_tile_24_31_to_tile_24_30_0;
	wire horizontal_tile_24_31_to_tile_24_30_1;
	wire horizontal_tile_24_31_to_tile_24_30_2;
	wire horizontal_tile_24_31_to_tile_24_30_3;

	wire horizontal_tile_25_30_to_tile_25_31_0;
	wire horizontal_tile_25_30_to_tile_25_31_1;
	wire horizontal_tile_25_30_to_tile_25_31_2;
	wire horizontal_tile_25_30_to_tile_25_31_3;
	wire horizontal_tile_25_31_to_tile_25_30_0;
	wire horizontal_tile_25_31_to_tile_25_30_1;
	wire horizontal_tile_25_31_to_tile_25_30_2;
	wire horizontal_tile_25_31_to_tile_25_30_3;

	wire horizontal_tile_26_30_to_tile_26_31_0;
	wire horizontal_tile_26_30_to_tile_26_31_1;
	wire horizontal_tile_26_30_to_tile_26_31_2;
	wire horizontal_tile_26_30_to_tile_26_31_3;
	wire horizontal_tile_26_31_to_tile_26_30_0;
	wire horizontal_tile_26_31_to_tile_26_30_1;
	wire horizontal_tile_26_31_to_tile_26_30_2;
	wire horizontal_tile_26_31_to_tile_26_30_3;

	wire horizontal_tile_27_30_to_tile_27_31_0;
	wire horizontal_tile_27_30_to_tile_27_31_1;
	wire horizontal_tile_27_30_to_tile_27_31_2;
	wire horizontal_tile_27_30_to_tile_27_31_3;
	wire horizontal_tile_27_31_to_tile_27_30_0;
	wire horizontal_tile_27_31_to_tile_27_30_1;
	wire horizontal_tile_27_31_to_tile_27_30_2;
	wire horizontal_tile_27_31_to_tile_27_30_3;

	wire horizontal_tile_28_30_to_tile_28_31_0;
	wire horizontal_tile_28_30_to_tile_28_31_1;
	wire horizontal_tile_28_30_to_tile_28_31_2;
	wire horizontal_tile_28_30_to_tile_28_31_3;
	wire horizontal_tile_28_31_to_tile_28_30_0;
	wire horizontal_tile_28_31_to_tile_28_30_1;
	wire horizontal_tile_28_31_to_tile_28_30_2;
	wire horizontal_tile_28_31_to_tile_28_30_3;

	wire horizontal_tile_29_30_to_tile_29_31_0;
	wire horizontal_tile_29_30_to_tile_29_31_1;
	wire horizontal_tile_29_30_to_tile_29_31_2;
	wire horizontal_tile_29_30_to_tile_29_31_3;
	wire horizontal_tile_29_31_to_tile_29_30_0;
	wire horizontal_tile_29_31_to_tile_29_30_1;
	wire horizontal_tile_29_31_to_tile_29_30_2;
	wire horizontal_tile_29_31_to_tile_29_30_3;

	wire horizontal_tile_30_30_to_tile_30_31_0;
	wire horizontal_tile_30_30_to_tile_30_31_1;
	wire horizontal_tile_30_30_to_tile_30_31_2;
	wire horizontal_tile_30_30_to_tile_30_31_3;
	wire horizontal_tile_30_31_to_tile_30_30_0;
	wire horizontal_tile_30_31_to_tile_30_30_1;
	wire horizontal_tile_30_31_to_tile_30_30_2;
	wire horizontal_tile_30_31_to_tile_30_30_3;

	wire horizontal_tile_31_30_to_tile_31_31_0;
	wire horizontal_tile_31_30_to_tile_31_31_1;
	wire horizontal_tile_31_30_to_tile_31_31_2;
	wire horizontal_tile_31_30_to_tile_31_31_3;
	wire horizontal_tile_31_31_to_tile_31_30_0;
	wire horizontal_tile_31_31_to_tile_31_30_1;
	wire horizontal_tile_31_31_to_tile_31_30_2;
	wire horizontal_tile_31_31_to_tile_31_30_3;

	// Tile declarations
	pe_tile_top_left pe_tile_0_0(
		.in_wire_3_0(input_to_grid_0),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_0_to_tile_1_0_0),
		.out_wire_1_1(vertical_tile_0_0_to_tile_1_0_1),
		.out_wire_1_2(vertical_tile_0_0_to_tile_1_0_2),
		.out_wire_1_3(vertical_tile_0_0_to_tile_1_0_3),
		.in_wire_1_0(vertical_tile_1_0_to_tile_0_0_0),
		.in_wire_1_1(vertical_tile_1_0_to_tile_0_0_1),
		.in_wire_1_2(vertical_tile_1_0_to_tile_0_0_2),
		.in_wire_1_3(vertical_tile_1_0_to_tile_0_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_0_0_to_tile_0_1_0),
		.out_wire_0_1(horizontal_tile_0_0_to_tile_0_1_1),
		.out_wire_0_2(horizontal_tile_0_0_to_tile_0_1_2),
		.out_wire_0_3(horizontal_tile_0_0_to_tile_0_1_3),
		.in_wire_0_0(horizontal_tile_0_1_to_tile_0_0_0),
		.in_wire_0_1(horizontal_tile_0_1_to_tile_0_0_1),
		.in_wire_0_2(horizontal_tile_0_1_to_tile_0_0_2),
		.in_wire_0_3(horizontal_tile_0_1_to_tile_0_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1)
	);

	pe_tile_top pe_tile_0_1(
		.in_wire_3_0(input_to_grid_1),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_1_to_tile_1_1_0),
		.out_wire_1_1(vertical_tile_0_1_to_tile_1_1_1),
		.out_wire_1_2(vertical_tile_0_1_to_tile_1_1_2),
		.out_wire_1_3(vertical_tile_0_1_to_tile_1_1_3),
		.in_wire_1_0(vertical_tile_1_1_to_tile_0_1_0),
		.in_wire_1_1(vertical_tile_1_1_to_tile_0_1_1),
		.in_wire_1_2(vertical_tile_1_1_to_tile_0_1_2),
		.in_wire_1_3(vertical_tile_1_1_to_tile_0_1_3),
		.out_wire_2_0(horizontal_tile_0_1_to_tile_0_0_0),
		.out_wire_2_1(horizontal_tile_0_1_to_tile_0_0_1),
		.out_wire_2_2(horizontal_tile_0_1_to_tile_0_0_2),
		.out_wire_2_3(horizontal_tile_0_1_to_tile_0_0_3),
		.in_wire_2_0(horizontal_tile_0_0_to_tile_0_1_0),
		.in_wire_2_1(horizontal_tile_0_0_to_tile_0_1_1),
		.in_wire_2_2(horizontal_tile_0_0_to_tile_0_1_2),
		.in_wire_2_3(horizontal_tile_0_0_to_tile_0_1_3),
		.out_wire_0_0(horizontal_tile_0_1_to_tile_0_2_0),
		.out_wire_0_1(horizontal_tile_0_1_to_tile_0_2_1),
		.out_wire_0_2(horizontal_tile_0_1_to_tile_0_2_2),
		.out_wire_0_3(horizontal_tile_0_1_to_tile_0_2_3),
		.in_wire_0_0(horizontal_tile_0_2_to_tile_0_1_0),
		.in_wire_0_1(horizontal_tile_0_2_to_tile_0_1_1),
		.in_wire_0_2(horizontal_tile_0_2_to_tile_0_1_2),
		.in_wire_0_3(horizontal_tile_0_2_to_tile_0_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(2)
	);

	pe_tile_top pe_tile_0_2(
		.in_wire_3_0(input_to_grid_2),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_2_to_tile_1_2_0),
		.out_wire_1_1(vertical_tile_0_2_to_tile_1_2_1),
		.out_wire_1_2(vertical_tile_0_2_to_tile_1_2_2),
		.out_wire_1_3(vertical_tile_0_2_to_tile_1_2_3),
		.in_wire_1_0(vertical_tile_1_2_to_tile_0_2_0),
		.in_wire_1_1(vertical_tile_1_2_to_tile_0_2_1),
		.in_wire_1_2(vertical_tile_1_2_to_tile_0_2_2),
		.in_wire_1_3(vertical_tile_1_2_to_tile_0_2_3),
		.out_wire_2_0(horizontal_tile_0_2_to_tile_0_1_0),
		.out_wire_2_1(horizontal_tile_0_2_to_tile_0_1_1),
		.out_wire_2_2(horizontal_tile_0_2_to_tile_0_1_2),
		.out_wire_2_3(horizontal_tile_0_2_to_tile_0_1_3),
		.in_wire_2_0(horizontal_tile_0_1_to_tile_0_2_0),
		.in_wire_2_1(horizontal_tile_0_1_to_tile_0_2_1),
		.in_wire_2_2(horizontal_tile_0_1_to_tile_0_2_2),
		.in_wire_2_3(horizontal_tile_0_1_to_tile_0_2_3),
		.out_wire_0_0(horizontal_tile_0_2_to_tile_0_3_0),
		.out_wire_0_1(horizontal_tile_0_2_to_tile_0_3_1),
		.out_wire_0_2(horizontal_tile_0_2_to_tile_0_3_2),
		.out_wire_0_3(horizontal_tile_0_2_to_tile_0_3_3),
		.in_wire_0_0(horizontal_tile_0_3_to_tile_0_2_0),
		.in_wire_0_1(horizontal_tile_0_3_to_tile_0_2_1),
		.in_wire_0_2(horizontal_tile_0_3_to_tile_0_2_2),
		.in_wire_0_3(horizontal_tile_0_3_to_tile_0_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(3)
	);

	pe_tile_top pe_tile_0_3(
		.in_wire_3_0(input_to_grid_3),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_3_to_tile_1_3_0),
		.out_wire_1_1(vertical_tile_0_3_to_tile_1_3_1),
		.out_wire_1_2(vertical_tile_0_3_to_tile_1_3_2),
		.out_wire_1_3(vertical_tile_0_3_to_tile_1_3_3),
		.in_wire_1_0(vertical_tile_1_3_to_tile_0_3_0),
		.in_wire_1_1(vertical_tile_1_3_to_tile_0_3_1),
		.in_wire_1_2(vertical_tile_1_3_to_tile_0_3_2),
		.in_wire_1_3(vertical_tile_1_3_to_tile_0_3_3),
		.out_wire_2_0(horizontal_tile_0_3_to_tile_0_2_0),
		.out_wire_2_1(horizontal_tile_0_3_to_tile_0_2_1),
		.out_wire_2_2(horizontal_tile_0_3_to_tile_0_2_2),
		.out_wire_2_3(horizontal_tile_0_3_to_tile_0_2_3),
		.in_wire_2_0(horizontal_tile_0_2_to_tile_0_3_0),
		.in_wire_2_1(horizontal_tile_0_2_to_tile_0_3_1),
		.in_wire_2_2(horizontal_tile_0_2_to_tile_0_3_2),
		.in_wire_2_3(horizontal_tile_0_2_to_tile_0_3_3),
		.out_wire_0_0(horizontal_tile_0_3_to_tile_0_4_0),
		.out_wire_0_1(horizontal_tile_0_3_to_tile_0_4_1),
		.out_wire_0_2(horizontal_tile_0_3_to_tile_0_4_2),
		.out_wire_0_3(horizontal_tile_0_3_to_tile_0_4_3),
		.in_wire_0_0(horizontal_tile_0_4_to_tile_0_3_0),
		.in_wire_0_1(horizontal_tile_0_4_to_tile_0_3_1),
		.in_wire_0_2(horizontal_tile_0_4_to_tile_0_3_2),
		.in_wire_0_3(horizontal_tile_0_4_to_tile_0_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(4)
	);

	pe_tile_top pe_tile_0_4(
		.in_wire_3_0(input_to_grid_4),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_4_to_tile_1_4_0),
		.out_wire_1_1(vertical_tile_0_4_to_tile_1_4_1),
		.out_wire_1_2(vertical_tile_0_4_to_tile_1_4_2),
		.out_wire_1_3(vertical_tile_0_4_to_tile_1_4_3),
		.in_wire_1_0(vertical_tile_1_4_to_tile_0_4_0),
		.in_wire_1_1(vertical_tile_1_4_to_tile_0_4_1),
		.in_wire_1_2(vertical_tile_1_4_to_tile_0_4_2),
		.in_wire_1_3(vertical_tile_1_4_to_tile_0_4_3),
		.out_wire_2_0(horizontal_tile_0_4_to_tile_0_3_0),
		.out_wire_2_1(horizontal_tile_0_4_to_tile_0_3_1),
		.out_wire_2_2(horizontal_tile_0_4_to_tile_0_3_2),
		.out_wire_2_3(horizontal_tile_0_4_to_tile_0_3_3),
		.in_wire_2_0(horizontal_tile_0_3_to_tile_0_4_0),
		.in_wire_2_1(horizontal_tile_0_3_to_tile_0_4_1),
		.in_wire_2_2(horizontal_tile_0_3_to_tile_0_4_2),
		.in_wire_2_3(horizontal_tile_0_3_to_tile_0_4_3),
		.out_wire_0_0(horizontal_tile_0_4_to_tile_0_5_0),
		.out_wire_0_1(horizontal_tile_0_4_to_tile_0_5_1),
		.out_wire_0_2(horizontal_tile_0_4_to_tile_0_5_2),
		.out_wire_0_3(horizontal_tile_0_4_to_tile_0_5_3),
		.in_wire_0_0(horizontal_tile_0_5_to_tile_0_4_0),
		.in_wire_0_1(horizontal_tile_0_5_to_tile_0_4_1),
		.in_wire_0_2(horizontal_tile_0_5_to_tile_0_4_2),
		.in_wire_0_3(horizontal_tile_0_5_to_tile_0_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(5)
	);

	pe_tile_top pe_tile_0_5(
		.in_wire_3_0(input_to_grid_5),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_5_to_tile_1_5_0),
		.out_wire_1_1(vertical_tile_0_5_to_tile_1_5_1),
		.out_wire_1_2(vertical_tile_0_5_to_tile_1_5_2),
		.out_wire_1_3(vertical_tile_0_5_to_tile_1_5_3),
		.in_wire_1_0(vertical_tile_1_5_to_tile_0_5_0),
		.in_wire_1_1(vertical_tile_1_5_to_tile_0_5_1),
		.in_wire_1_2(vertical_tile_1_5_to_tile_0_5_2),
		.in_wire_1_3(vertical_tile_1_5_to_tile_0_5_3),
		.out_wire_2_0(horizontal_tile_0_5_to_tile_0_4_0),
		.out_wire_2_1(horizontal_tile_0_5_to_tile_0_4_1),
		.out_wire_2_2(horizontal_tile_0_5_to_tile_0_4_2),
		.out_wire_2_3(horizontal_tile_0_5_to_tile_0_4_3),
		.in_wire_2_0(horizontal_tile_0_4_to_tile_0_5_0),
		.in_wire_2_1(horizontal_tile_0_4_to_tile_0_5_1),
		.in_wire_2_2(horizontal_tile_0_4_to_tile_0_5_2),
		.in_wire_2_3(horizontal_tile_0_4_to_tile_0_5_3),
		.out_wire_0_0(horizontal_tile_0_5_to_tile_0_6_0),
		.out_wire_0_1(horizontal_tile_0_5_to_tile_0_6_1),
		.out_wire_0_2(horizontal_tile_0_5_to_tile_0_6_2),
		.out_wire_0_3(horizontal_tile_0_5_to_tile_0_6_3),
		.in_wire_0_0(horizontal_tile_0_6_to_tile_0_5_0),
		.in_wire_0_1(horizontal_tile_0_6_to_tile_0_5_1),
		.in_wire_0_2(horizontal_tile_0_6_to_tile_0_5_2),
		.in_wire_0_3(horizontal_tile_0_6_to_tile_0_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(6)
	);

	pe_tile_top pe_tile_0_6(
		.in_wire_3_0(input_to_grid_6),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_6_to_tile_1_6_0),
		.out_wire_1_1(vertical_tile_0_6_to_tile_1_6_1),
		.out_wire_1_2(vertical_tile_0_6_to_tile_1_6_2),
		.out_wire_1_3(vertical_tile_0_6_to_tile_1_6_3),
		.in_wire_1_0(vertical_tile_1_6_to_tile_0_6_0),
		.in_wire_1_1(vertical_tile_1_6_to_tile_0_6_1),
		.in_wire_1_2(vertical_tile_1_6_to_tile_0_6_2),
		.in_wire_1_3(vertical_tile_1_6_to_tile_0_6_3),
		.out_wire_2_0(horizontal_tile_0_6_to_tile_0_5_0),
		.out_wire_2_1(horizontal_tile_0_6_to_tile_0_5_1),
		.out_wire_2_2(horizontal_tile_0_6_to_tile_0_5_2),
		.out_wire_2_3(horizontal_tile_0_6_to_tile_0_5_3),
		.in_wire_2_0(horizontal_tile_0_5_to_tile_0_6_0),
		.in_wire_2_1(horizontal_tile_0_5_to_tile_0_6_1),
		.in_wire_2_2(horizontal_tile_0_5_to_tile_0_6_2),
		.in_wire_2_3(horizontal_tile_0_5_to_tile_0_6_3),
		.out_wire_0_0(horizontal_tile_0_6_to_tile_0_7_0),
		.out_wire_0_1(horizontal_tile_0_6_to_tile_0_7_1),
		.out_wire_0_2(horizontal_tile_0_6_to_tile_0_7_2),
		.out_wire_0_3(horizontal_tile_0_6_to_tile_0_7_3),
		.in_wire_0_0(horizontal_tile_0_7_to_tile_0_6_0),
		.in_wire_0_1(horizontal_tile_0_7_to_tile_0_6_1),
		.in_wire_0_2(horizontal_tile_0_7_to_tile_0_6_2),
		.in_wire_0_3(horizontal_tile_0_7_to_tile_0_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(7)
	);

	pe_tile_top pe_tile_0_7(
		.in_wire_3_0(input_to_grid_7),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_7_to_tile_1_7_0),
		.out_wire_1_1(vertical_tile_0_7_to_tile_1_7_1),
		.out_wire_1_2(vertical_tile_0_7_to_tile_1_7_2),
		.out_wire_1_3(vertical_tile_0_7_to_tile_1_7_3),
		.in_wire_1_0(vertical_tile_1_7_to_tile_0_7_0),
		.in_wire_1_1(vertical_tile_1_7_to_tile_0_7_1),
		.in_wire_1_2(vertical_tile_1_7_to_tile_0_7_2),
		.in_wire_1_3(vertical_tile_1_7_to_tile_0_7_3),
		.out_wire_2_0(horizontal_tile_0_7_to_tile_0_6_0),
		.out_wire_2_1(horizontal_tile_0_7_to_tile_0_6_1),
		.out_wire_2_2(horizontal_tile_0_7_to_tile_0_6_2),
		.out_wire_2_3(horizontal_tile_0_7_to_tile_0_6_3),
		.in_wire_2_0(horizontal_tile_0_6_to_tile_0_7_0),
		.in_wire_2_1(horizontal_tile_0_6_to_tile_0_7_1),
		.in_wire_2_2(horizontal_tile_0_6_to_tile_0_7_2),
		.in_wire_2_3(horizontal_tile_0_6_to_tile_0_7_3),
		.out_wire_0_0(horizontal_tile_0_7_to_tile_0_8_0),
		.out_wire_0_1(horizontal_tile_0_7_to_tile_0_8_1),
		.out_wire_0_2(horizontal_tile_0_7_to_tile_0_8_2),
		.out_wire_0_3(horizontal_tile_0_7_to_tile_0_8_3),
		.in_wire_0_0(horizontal_tile_0_8_to_tile_0_7_0),
		.in_wire_0_1(horizontal_tile_0_8_to_tile_0_7_1),
		.in_wire_0_2(horizontal_tile_0_8_to_tile_0_7_2),
		.in_wire_0_3(horizontal_tile_0_8_to_tile_0_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(8)
	);

	pe_tile_top pe_tile_0_8(
		.in_wire_3_0(input_to_grid_8),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_8_to_tile_1_8_0),
		.out_wire_1_1(vertical_tile_0_8_to_tile_1_8_1),
		.out_wire_1_2(vertical_tile_0_8_to_tile_1_8_2),
		.out_wire_1_3(vertical_tile_0_8_to_tile_1_8_3),
		.in_wire_1_0(vertical_tile_1_8_to_tile_0_8_0),
		.in_wire_1_1(vertical_tile_1_8_to_tile_0_8_1),
		.in_wire_1_2(vertical_tile_1_8_to_tile_0_8_2),
		.in_wire_1_3(vertical_tile_1_8_to_tile_0_8_3),
		.out_wire_2_0(horizontal_tile_0_8_to_tile_0_7_0),
		.out_wire_2_1(horizontal_tile_0_8_to_tile_0_7_1),
		.out_wire_2_2(horizontal_tile_0_8_to_tile_0_7_2),
		.out_wire_2_3(horizontal_tile_0_8_to_tile_0_7_3),
		.in_wire_2_0(horizontal_tile_0_7_to_tile_0_8_0),
		.in_wire_2_1(horizontal_tile_0_7_to_tile_0_8_1),
		.in_wire_2_2(horizontal_tile_0_7_to_tile_0_8_2),
		.in_wire_2_3(horizontal_tile_0_7_to_tile_0_8_3),
		.out_wire_0_0(horizontal_tile_0_8_to_tile_0_9_0),
		.out_wire_0_1(horizontal_tile_0_8_to_tile_0_9_1),
		.out_wire_0_2(horizontal_tile_0_8_to_tile_0_9_2),
		.out_wire_0_3(horizontal_tile_0_8_to_tile_0_9_3),
		.in_wire_0_0(horizontal_tile_0_9_to_tile_0_8_0),
		.in_wire_0_1(horizontal_tile_0_9_to_tile_0_8_1),
		.in_wire_0_2(horizontal_tile_0_9_to_tile_0_8_2),
		.in_wire_0_3(horizontal_tile_0_9_to_tile_0_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(9)
	);

	pe_tile_top pe_tile_0_9(
		.in_wire_3_0(input_to_grid_9),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_9_to_tile_1_9_0),
		.out_wire_1_1(vertical_tile_0_9_to_tile_1_9_1),
		.out_wire_1_2(vertical_tile_0_9_to_tile_1_9_2),
		.out_wire_1_3(vertical_tile_0_9_to_tile_1_9_3),
		.in_wire_1_0(vertical_tile_1_9_to_tile_0_9_0),
		.in_wire_1_1(vertical_tile_1_9_to_tile_0_9_1),
		.in_wire_1_2(vertical_tile_1_9_to_tile_0_9_2),
		.in_wire_1_3(vertical_tile_1_9_to_tile_0_9_3),
		.out_wire_2_0(horizontal_tile_0_9_to_tile_0_8_0),
		.out_wire_2_1(horizontal_tile_0_9_to_tile_0_8_1),
		.out_wire_2_2(horizontal_tile_0_9_to_tile_0_8_2),
		.out_wire_2_3(horizontal_tile_0_9_to_tile_0_8_3),
		.in_wire_2_0(horizontal_tile_0_8_to_tile_0_9_0),
		.in_wire_2_1(horizontal_tile_0_8_to_tile_0_9_1),
		.in_wire_2_2(horizontal_tile_0_8_to_tile_0_9_2),
		.in_wire_2_3(horizontal_tile_0_8_to_tile_0_9_3),
		.out_wire_0_0(horizontal_tile_0_9_to_tile_0_10_0),
		.out_wire_0_1(horizontal_tile_0_9_to_tile_0_10_1),
		.out_wire_0_2(horizontal_tile_0_9_to_tile_0_10_2),
		.out_wire_0_3(horizontal_tile_0_9_to_tile_0_10_3),
		.in_wire_0_0(horizontal_tile_0_10_to_tile_0_9_0),
		.in_wire_0_1(horizontal_tile_0_10_to_tile_0_9_1),
		.in_wire_0_2(horizontal_tile_0_10_to_tile_0_9_2),
		.in_wire_0_3(horizontal_tile_0_10_to_tile_0_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(10)
	);

	pe_tile_top pe_tile_0_10(
		.in_wire_3_0(input_to_grid_10),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_10_to_tile_1_10_0),
		.out_wire_1_1(vertical_tile_0_10_to_tile_1_10_1),
		.out_wire_1_2(vertical_tile_0_10_to_tile_1_10_2),
		.out_wire_1_3(vertical_tile_0_10_to_tile_1_10_3),
		.in_wire_1_0(vertical_tile_1_10_to_tile_0_10_0),
		.in_wire_1_1(vertical_tile_1_10_to_tile_0_10_1),
		.in_wire_1_2(vertical_tile_1_10_to_tile_0_10_2),
		.in_wire_1_3(vertical_tile_1_10_to_tile_0_10_3),
		.out_wire_2_0(horizontal_tile_0_10_to_tile_0_9_0),
		.out_wire_2_1(horizontal_tile_0_10_to_tile_0_9_1),
		.out_wire_2_2(horizontal_tile_0_10_to_tile_0_9_2),
		.out_wire_2_3(horizontal_tile_0_10_to_tile_0_9_3),
		.in_wire_2_0(horizontal_tile_0_9_to_tile_0_10_0),
		.in_wire_2_1(horizontal_tile_0_9_to_tile_0_10_1),
		.in_wire_2_2(horizontal_tile_0_9_to_tile_0_10_2),
		.in_wire_2_3(horizontal_tile_0_9_to_tile_0_10_3),
		.out_wire_0_0(horizontal_tile_0_10_to_tile_0_11_0),
		.out_wire_0_1(horizontal_tile_0_10_to_tile_0_11_1),
		.out_wire_0_2(horizontal_tile_0_10_to_tile_0_11_2),
		.out_wire_0_3(horizontal_tile_0_10_to_tile_0_11_3),
		.in_wire_0_0(horizontal_tile_0_11_to_tile_0_10_0),
		.in_wire_0_1(horizontal_tile_0_11_to_tile_0_10_1),
		.in_wire_0_2(horizontal_tile_0_11_to_tile_0_10_2),
		.in_wire_0_3(horizontal_tile_0_11_to_tile_0_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(11)
	);

	pe_tile_top pe_tile_0_11(
		.in_wire_3_0(input_to_grid_11),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_11_to_tile_1_11_0),
		.out_wire_1_1(vertical_tile_0_11_to_tile_1_11_1),
		.out_wire_1_2(vertical_tile_0_11_to_tile_1_11_2),
		.out_wire_1_3(vertical_tile_0_11_to_tile_1_11_3),
		.in_wire_1_0(vertical_tile_1_11_to_tile_0_11_0),
		.in_wire_1_1(vertical_tile_1_11_to_tile_0_11_1),
		.in_wire_1_2(vertical_tile_1_11_to_tile_0_11_2),
		.in_wire_1_3(vertical_tile_1_11_to_tile_0_11_3),
		.out_wire_2_0(horizontal_tile_0_11_to_tile_0_10_0),
		.out_wire_2_1(horizontal_tile_0_11_to_tile_0_10_1),
		.out_wire_2_2(horizontal_tile_0_11_to_tile_0_10_2),
		.out_wire_2_3(horizontal_tile_0_11_to_tile_0_10_3),
		.in_wire_2_0(horizontal_tile_0_10_to_tile_0_11_0),
		.in_wire_2_1(horizontal_tile_0_10_to_tile_0_11_1),
		.in_wire_2_2(horizontal_tile_0_10_to_tile_0_11_2),
		.in_wire_2_3(horizontal_tile_0_10_to_tile_0_11_3),
		.out_wire_0_0(horizontal_tile_0_11_to_tile_0_12_0),
		.out_wire_0_1(horizontal_tile_0_11_to_tile_0_12_1),
		.out_wire_0_2(horizontal_tile_0_11_to_tile_0_12_2),
		.out_wire_0_3(horizontal_tile_0_11_to_tile_0_12_3),
		.in_wire_0_0(horizontal_tile_0_12_to_tile_0_11_0),
		.in_wire_0_1(horizontal_tile_0_12_to_tile_0_11_1),
		.in_wire_0_2(horizontal_tile_0_12_to_tile_0_11_2),
		.in_wire_0_3(horizontal_tile_0_12_to_tile_0_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(12)
	);

	pe_tile_top pe_tile_0_12(
		.in_wire_3_0(input_to_grid_12),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_12_to_tile_1_12_0),
		.out_wire_1_1(vertical_tile_0_12_to_tile_1_12_1),
		.out_wire_1_2(vertical_tile_0_12_to_tile_1_12_2),
		.out_wire_1_3(vertical_tile_0_12_to_tile_1_12_3),
		.in_wire_1_0(vertical_tile_1_12_to_tile_0_12_0),
		.in_wire_1_1(vertical_tile_1_12_to_tile_0_12_1),
		.in_wire_1_2(vertical_tile_1_12_to_tile_0_12_2),
		.in_wire_1_3(vertical_tile_1_12_to_tile_0_12_3),
		.out_wire_2_0(horizontal_tile_0_12_to_tile_0_11_0),
		.out_wire_2_1(horizontal_tile_0_12_to_tile_0_11_1),
		.out_wire_2_2(horizontal_tile_0_12_to_tile_0_11_2),
		.out_wire_2_3(horizontal_tile_0_12_to_tile_0_11_3),
		.in_wire_2_0(horizontal_tile_0_11_to_tile_0_12_0),
		.in_wire_2_1(horizontal_tile_0_11_to_tile_0_12_1),
		.in_wire_2_2(horizontal_tile_0_11_to_tile_0_12_2),
		.in_wire_2_3(horizontal_tile_0_11_to_tile_0_12_3),
		.out_wire_0_0(horizontal_tile_0_12_to_tile_0_13_0),
		.out_wire_0_1(horizontal_tile_0_12_to_tile_0_13_1),
		.out_wire_0_2(horizontal_tile_0_12_to_tile_0_13_2),
		.out_wire_0_3(horizontal_tile_0_12_to_tile_0_13_3),
		.in_wire_0_0(horizontal_tile_0_13_to_tile_0_12_0),
		.in_wire_0_1(horizontal_tile_0_13_to_tile_0_12_1),
		.in_wire_0_2(horizontal_tile_0_13_to_tile_0_12_2),
		.in_wire_0_3(horizontal_tile_0_13_to_tile_0_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(13)
	);

	pe_tile_top pe_tile_0_13(
		.in_wire_3_0(input_to_grid_13),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_13_to_tile_1_13_0),
		.out_wire_1_1(vertical_tile_0_13_to_tile_1_13_1),
		.out_wire_1_2(vertical_tile_0_13_to_tile_1_13_2),
		.out_wire_1_3(vertical_tile_0_13_to_tile_1_13_3),
		.in_wire_1_0(vertical_tile_1_13_to_tile_0_13_0),
		.in_wire_1_1(vertical_tile_1_13_to_tile_0_13_1),
		.in_wire_1_2(vertical_tile_1_13_to_tile_0_13_2),
		.in_wire_1_3(vertical_tile_1_13_to_tile_0_13_3),
		.out_wire_2_0(horizontal_tile_0_13_to_tile_0_12_0),
		.out_wire_2_1(horizontal_tile_0_13_to_tile_0_12_1),
		.out_wire_2_2(horizontal_tile_0_13_to_tile_0_12_2),
		.out_wire_2_3(horizontal_tile_0_13_to_tile_0_12_3),
		.in_wire_2_0(horizontal_tile_0_12_to_tile_0_13_0),
		.in_wire_2_1(horizontal_tile_0_12_to_tile_0_13_1),
		.in_wire_2_2(horizontal_tile_0_12_to_tile_0_13_2),
		.in_wire_2_3(horizontal_tile_0_12_to_tile_0_13_3),
		.out_wire_0_0(horizontal_tile_0_13_to_tile_0_14_0),
		.out_wire_0_1(horizontal_tile_0_13_to_tile_0_14_1),
		.out_wire_0_2(horizontal_tile_0_13_to_tile_0_14_2),
		.out_wire_0_3(horizontal_tile_0_13_to_tile_0_14_3),
		.in_wire_0_0(horizontal_tile_0_14_to_tile_0_13_0),
		.in_wire_0_1(horizontal_tile_0_14_to_tile_0_13_1),
		.in_wire_0_2(horizontal_tile_0_14_to_tile_0_13_2),
		.in_wire_0_3(horizontal_tile_0_14_to_tile_0_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(14)
	);

	pe_tile_top pe_tile_0_14(
		.in_wire_3_0(input_to_grid_14),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_14_to_tile_1_14_0),
		.out_wire_1_1(vertical_tile_0_14_to_tile_1_14_1),
		.out_wire_1_2(vertical_tile_0_14_to_tile_1_14_2),
		.out_wire_1_3(vertical_tile_0_14_to_tile_1_14_3),
		.in_wire_1_0(vertical_tile_1_14_to_tile_0_14_0),
		.in_wire_1_1(vertical_tile_1_14_to_tile_0_14_1),
		.in_wire_1_2(vertical_tile_1_14_to_tile_0_14_2),
		.in_wire_1_3(vertical_tile_1_14_to_tile_0_14_3),
		.out_wire_2_0(horizontal_tile_0_14_to_tile_0_13_0),
		.out_wire_2_1(horizontal_tile_0_14_to_tile_0_13_1),
		.out_wire_2_2(horizontal_tile_0_14_to_tile_0_13_2),
		.out_wire_2_3(horizontal_tile_0_14_to_tile_0_13_3),
		.in_wire_2_0(horizontal_tile_0_13_to_tile_0_14_0),
		.in_wire_2_1(horizontal_tile_0_13_to_tile_0_14_1),
		.in_wire_2_2(horizontal_tile_0_13_to_tile_0_14_2),
		.in_wire_2_3(horizontal_tile_0_13_to_tile_0_14_3),
		.out_wire_0_0(horizontal_tile_0_14_to_tile_0_15_0),
		.out_wire_0_1(horizontal_tile_0_14_to_tile_0_15_1),
		.out_wire_0_2(horizontal_tile_0_14_to_tile_0_15_2),
		.out_wire_0_3(horizontal_tile_0_14_to_tile_0_15_3),
		.in_wire_0_0(horizontal_tile_0_15_to_tile_0_14_0),
		.in_wire_0_1(horizontal_tile_0_15_to_tile_0_14_1),
		.in_wire_0_2(horizontal_tile_0_15_to_tile_0_14_2),
		.in_wire_0_3(horizontal_tile_0_15_to_tile_0_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(15)
	);

	pe_tile_top pe_tile_0_15(
		.in_wire_3_0(input_to_grid_15),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_15_to_tile_1_15_0),
		.out_wire_1_1(vertical_tile_0_15_to_tile_1_15_1),
		.out_wire_1_2(vertical_tile_0_15_to_tile_1_15_2),
		.out_wire_1_3(vertical_tile_0_15_to_tile_1_15_3),
		.in_wire_1_0(vertical_tile_1_15_to_tile_0_15_0),
		.in_wire_1_1(vertical_tile_1_15_to_tile_0_15_1),
		.in_wire_1_2(vertical_tile_1_15_to_tile_0_15_2),
		.in_wire_1_3(vertical_tile_1_15_to_tile_0_15_3),
		.out_wire_2_0(horizontal_tile_0_15_to_tile_0_14_0),
		.out_wire_2_1(horizontal_tile_0_15_to_tile_0_14_1),
		.out_wire_2_2(horizontal_tile_0_15_to_tile_0_14_2),
		.out_wire_2_3(horizontal_tile_0_15_to_tile_0_14_3),
		.in_wire_2_0(horizontal_tile_0_14_to_tile_0_15_0),
		.in_wire_2_1(horizontal_tile_0_14_to_tile_0_15_1),
		.in_wire_2_2(horizontal_tile_0_14_to_tile_0_15_2),
		.in_wire_2_3(horizontal_tile_0_14_to_tile_0_15_3),
		.out_wire_0_0(horizontal_tile_0_15_to_tile_0_16_0),
		.out_wire_0_1(horizontal_tile_0_15_to_tile_0_16_1),
		.out_wire_0_2(horizontal_tile_0_15_to_tile_0_16_2),
		.out_wire_0_3(horizontal_tile_0_15_to_tile_0_16_3),
		.in_wire_0_0(horizontal_tile_0_16_to_tile_0_15_0),
		.in_wire_0_1(horizontal_tile_0_16_to_tile_0_15_1),
		.in_wire_0_2(horizontal_tile_0_16_to_tile_0_15_2),
		.in_wire_0_3(horizontal_tile_0_16_to_tile_0_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(16)
	);

	pe_tile_top pe_tile_0_16(
		.in_wire_3_0(input_to_grid_16),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_16_to_tile_1_16_0),
		.out_wire_1_1(vertical_tile_0_16_to_tile_1_16_1),
		.out_wire_1_2(vertical_tile_0_16_to_tile_1_16_2),
		.out_wire_1_3(vertical_tile_0_16_to_tile_1_16_3),
		.in_wire_1_0(vertical_tile_1_16_to_tile_0_16_0),
		.in_wire_1_1(vertical_tile_1_16_to_tile_0_16_1),
		.in_wire_1_2(vertical_tile_1_16_to_tile_0_16_2),
		.in_wire_1_3(vertical_tile_1_16_to_tile_0_16_3),
		.out_wire_2_0(horizontal_tile_0_16_to_tile_0_15_0),
		.out_wire_2_1(horizontal_tile_0_16_to_tile_0_15_1),
		.out_wire_2_2(horizontal_tile_0_16_to_tile_0_15_2),
		.out_wire_2_3(horizontal_tile_0_16_to_tile_0_15_3),
		.in_wire_2_0(horizontal_tile_0_15_to_tile_0_16_0),
		.in_wire_2_1(horizontal_tile_0_15_to_tile_0_16_1),
		.in_wire_2_2(horizontal_tile_0_15_to_tile_0_16_2),
		.in_wire_2_3(horizontal_tile_0_15_to_tile_0_16_3),
		.out_wire_0_0(horizontal_tile_0_16_to_tile_0_17_0),
		.out_wire_0_1(horizontal_tile_0_16_to_tile_0_17_1),
		.out_wire_0_2(horizontal_tile_0_16_to_tile_0_17_2),
		.out_wire_0_3(horizontal_tile_0_16_to_tile_0_17_3),
		.in_wire_0_0(horizontal_tile_0_17_to_tile_0_16_0),
		.in_wire_0_1(horizontal_tile_0_17_to_tile_0_16_1),
		.in_wire_0_2(horizontal_tile_0_17_to_tile_0_16_2),
		.in_wire_0_3(horizontal_tile_0_17_to_tile_0_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(17)
	);

	pe_tile_top pe_tile_0_17(
		.in_wire_3_0(input_to_grid_17),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_17_to_tile_1_17_0),
		.out_wire_1_1(vertical_tile_0_17_to_tile_1_17_1),
		.out_wire_1_2(vertical_tile_0_17_to_tile_1_17_2),
		.out_wire_1_3(vertical_tile_0_17_to_tile_1_17_3),
		.in_wire_1_0(vertical_tile_1_17_to_tile_0_17_0),
		.in_wire_1_1(vertical_tile_1_17_to_tile_0_17_1),
		.in_wire_1_2(vertical_tile_1_17_to_tile_0_17_2),
		.in_wire_1_3(vertical_tile_1_17_to_tile_0_17_3),
		.out_wire_2_0(horizontal_tile_0_17_to_tile_0_16_0),
		.out_wire_2_1(horizontal_tile_0_17_to_tile_0_16_1),
		.out_wire_2_2(horizontal_tile_0_17_to_tile_0_16_2),
		.out_wire_2_3(horizontal_tile_0_17_to_tile_0_16_3),
		.in_wire_2_0(horizontal_tile_0_16_to_tile_0_17_0),
		.in_wire_2_1(horizontal_tile_0_16_to_tile_0_17_1),
		.in_wire_2_2(horizontal_tile_0_16_to_tile_0_17_2),
		.in_wire_2_3(horizontal_tile_0_16_to_tile_0_17_3),
		.out_wire_0_0(horizontal_tile_0_17_to_tile_0_18_0),
		.out_wire_0_1(horizontal_tile_0_17_to_tile_0_18_1),
		.out_wire_0_2(horizontal_tile_0_17_to_tile_0_18_2),
		.out_wire_0_3(horizontal_tile_0_17_to_tile_0_18_3),
		.in_wire_0_0(horizontal_tile_0_18_to_tile_0_17_0),
		.in_wire_0_1(horizontal_tile_0_18_to_tile_0_17_1),
		.in_wire_0_2(horizontal_tile_0_18_to_tile_0_17_2),
		.in_wire_0_3(horizontal_tile_0_18_to_tile_0_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(18)
	);

	pe_tile_top pe_tile_0_18(
		.in_wire_3_0(input_to_grid_18),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_18_to_tile_1_18_0),
		.out_wire_1_1(vertical_tile_0_18_to_tile_1_18_1),
		.out_wire_1_2(vertical_tile_0_18_to_tile_1_18_2),
		.out_wire_1_3(vertical_tile_0_18_to_tile_1_18_3),
		.in_wire_1_0(vertical_tile_1_18_to_tile_0_18_0),
		.in_wire_1_1(vertical_tile_1_18_to_tile_0_18_1),
		.in_wire_1_2(vertical_tile_1_18_to_tile_0_18_2),
		.in_wire_1_3(vertical_tile_1_18_to_tile_0_18_3),
		.out_wire_2_0(horizontal_tile_0_18_to_tile_0_17_0),
		.out_wire_2_1(horizontal_tile_0_18_to_tile_0_17_1),
		.out_wire_2_2(horizontal_tile_0_18_to_tile_0_17_2),
		.out_wire_2_3(horizontal_tile_0_18_to_tile_0_17_3),
		.in_wire_2_0(horizontal_tile_0_17_to_tile_0_18_0),
		.in_wire_2_1(horizontal_tile_0_17_to_tile_0_18_1),
		.in_wire_2_2(horizontal_tile_0_17_to_tile_0_18_2),
		.in_wire_2_3(horizontal_tile_0_17_to_tile_0_18_3),
		.out_wire_0_0(horizontal_tile_0_18_to_tile_0_19_0),
		.out_wire_0_1(horizontal_tile_0_18_to_tile_0_19_1),
		.out_wire_0_2(horizontal_tile_0_18_to_tile_0_19_2),
		.out_wire_0_3(horizontal_tile_0_18_to_tile_0_19_3),
		.in_wire_0_0(horizontal_tile_0_19_to_tile_0_18_0),
		.in_wire_0_1(horizontal_tile_0_19_to_tile_0_18_1),
		.in_wire_0_2(horizontal_tile_0_19_to_tile_0_18_2),
		.in_wire_0_3(horizontal_tile_0_19_to_tile_0_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(19)
	);

	pe_tile_top pe_tile_0_19(
		.in_wire_3_0(input_to_grid_19),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_19_to_tile_1_19_0),
		.out_wire_1_1(vertical_tile_0_19_to_tile_1_19_1),
		.out_wire_1_2(vertical_tile_0_19_to_tile_1_19_2),
		.out_wire_1_3(vertical_tile_0_19_to_tile_1_19_3),
		.in_wire_1_0(vertical_tile_1_19_to_tile_0_19_0),
		.in_wire_1_1(vertical_tile_1_19_to_tile_0_19_1),
		.in_wire_1_2(vertical_tile_1_19_to_tile_0_19_2),
		.in_wire_1_3(vertical_tile_1_19_to_tile_0_19_3),
		.out_wire_2_0(horizontal_tile_0_19_to_tile_0_18_0),
		.out_wire_2_1(horizontal_tile_0_19_to_tile_0_18_1),
		.out_wire_2_2(horizontal_tile_0_19_to_tile_0_18_2),
		.out_wire_2_3(horizontal_tile_0_19_to_tile_0_18_3),
		.in_wire_2_0(horizontal_tile_0_18_to_tile_0_19_0),
		.in_wire_2_1(horizontal_tile_0_18_to_tile_0_19_1),
		.in_wire_2_2(horizontal_tile_0_18_to_tile_0_19_2),
		.in_wire_2_3(horizontal_tile_0_18_to_tile_0_19_3),
		.out_wire_0_0(horizontal_tile_0_19_to_tile_0_20_0),
		.out_wire_0_1(horizontal_tile_0_19_to_tile_0_20_1),
		.out_wire_0_2(horizontal_tile_0_19_to_tile_0_20_2),
		.out_wire_0_3(horizontal_tile_0_19_to_tile_0_20_3),
		.in_wire_0_0(horizontal_tile_0_20_to_tile_0_19_0),
		.in_wire_0_1(horizontal_tile_0_20_to_tile_0_19_1),
		.in_wire_0_2(horizontal_tile_0_20_to_tile_0_19_2),
		.in_wire_0_3(horizontal_tile_0_20_to_tile_0_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(20)
	);

	pe_tile_top pe_tile_0_20(
		.in_wire_3_0(input_to_grid_20),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_20_to_tile_1_20_0),
		.out_wire_1_1(vertical_tile_0_20_to_tile_1_20_1),
		.out_wire_1_2(vertical_tile_0_20_to_tile_1_20_2),
		.out_wire_1_3(vertical_tile_0_20_to_tile_1_20_3),
		.in_wire_1_0(vertical_tile_1_20_to_tile_0_20_0),
		.in_wire_1_1(vertical_tile_1_20_to_tile_0_20_1),
		.in_wire_1_2(vertical_tile_1_20_to_tile_0_20_2),
		.in_wire_1_3(vertical_tile_1_20_to_tile_0_20_3),
		.out_wire_2_0(horizontal_tile_0_20_to_tile_0_19_0),
		.out_wire_2_1(horizontal_tile_0_20_to_tile_0_19_1),
		.out_wire_2_2(horizontal_tile_0_20_to_tile_0_19_2),
		.out_wire_2_3(horizontal_tile_0_20_to_tile_0_19_3),
		.in_wire_2_0(horizontal_tile_0_19_to_tile_0_20_0),
		.in_wire_2_1(horizontal_tile_0_19_to_tile_0_20_1),
		.in_wire_2_2(horizontal_tile_0_19_to_tile_0_20_2),
		.in_wire_2_3(horizontal_tile_0_19_to_tile_0_20_3),
		.out_wire_0_0(horizontal_tile_0_20_to_tile_0_21_0),
		.out_wire_0_1(horizontal_tile_0_20_to_tile_0_21_1),
		.out_wire_0_2(horizontal_tile_0_20_to_tile_0_21_2),
		.out_wire_0_3(horizontal_tile_0_20_to_tile_0_21_3),
		.in_wire_0_0(horizontal_tile_0_21_to_tile_0_20_0),
		.in_wire_0_1(horizontal_tile_0_21_to_tile_0_20_1),
		.in_wire_0_2(horizontal_tile_0_21_to_tile_0_20_2),
		.in_wire_0_3(horizontal_tile_0_21_to_tile_0_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(21)
	);

	pe_tile_top pe_tile_0_21(
		.in_wire_3_0(input_to_grid_21),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_21_to_tile_1_21_0),
		.out_wire_1_1(vertical_tile_0_21_to_tile_1_21_1),
		.out_wire_1_2(vertical_tile_0_21_to_tile_1_21_2),
		.out_wire_1_3(vertical_tile_0_21_to_tile_1_21_3),
		.in_wire_1_0(vertical_tile_1_21_to_tile_0_21_0),
		.in_wire_1_1(vertical_tile_1_21_to_tile_0_21_1),
		.in_wire_1_2(vertical_tile_1_21_to_tile_0_21_2),
		.in_wire_1_3(vertical_tile_1_21_to_tile_0_21_3),
		.out_wire_2_0(horizontal_tile_0_21_to_tile_0_20_0),
		.out_wire_2_1(horizontal_tile_0_21_to_tile_0_20_1),
		.out_wire_2_2(horizontal_tile_0_21_to_tile_0_20_2),
		.out_wire_2_3(horizontal_tile_0_21_to_tile_0_20_3),
		.in_wire_2_0(horizontal_tile_0_20_to_tile_0_21_0),
		.in_wire_2_1(horizontal_tile_0_20_to_tile_0_21_1),
		.in_wire_2_2(horizontal_tile_0_20_to_tile_0_21_2),
		.in_wire_2_3(horizontal_tile_0_20_to_tile_0_21_3),
		.out_wire_0_0(horizontal_tile_0_21_to_tile_0_22_0),
		.out_wire_0_1(horizontal_tile_0_21_to_tile_0_22_1),
		.out_wire_0_2(horizontal_tile_0_21_to_tile_0_22_2),
		.out_wire_0_3(horizontal_tile_0_21_to_tile_0_22_3),
		.in_wire_0_0(horizontal_tile_0_22_to_tile_0_21_0),
		.in_wire_0_1(horizontal_tile_0_22_to_tile_0_21_1),
		.in_wire_0_2(horizontal_tile_0_22_to_tile_0_21_2),
		.in_wire_0_3(horizontal_tile_0_22_to_tile_0_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(22)
	);

	pe_tile_top pe_tile_0_22(
		.in_wire_3_0(input_to_grid_22),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_22_to_tile_1_22_0),
		.out_wire_1_1(vertical_tile_0_22_to_tile_1_22_1),
		.out_wire_1_2(vertical_tile_0_22_to_tile_1_22_2),
		.out_wire_1_3(vertical_tile_0_22_to_tile_1_22_3),
		.in_wire_1_0(vertical_tile_1_22_to_tile_0_22_0),
		.in_wire_1_1(vertical_tile_1_22_to_tile_0_22_1),
		.in_wire_1_2(vertical_tile_1_22_to_tile_0_22_2),
		.in_wire_1_3(vertical_tile_1_22_to_tile_0_22_3),
		.out_wire_2_0(horizontal_tile_0_22_to_tile_0_21_0),
		.out_wire_2_1(horizontal_tile_0_22_to_tile_0_21_1),
		.out_wire_2_2(horizontal_tile_0_22_to_tile_0_21_2),
		.out_wire_2_3(horizontal_tile_0_22_to_tile_0_21_3),
		.in_wire_2_0(horizontal_tile_0_21_to_tile_0_22_0),
		.in_wire_2_1(horizontal_tile_0_21_to_tile_0_22_1),
		.in_wire_2_2(horizontal_tile_0_21_to_tile_0_22_2),
		.in_wire_2_3(horizontal_tile_0_21_to_tile_0_22_3),
		.out_wire_0_0(horizontal_tile_0_22_to_tile_0_23_0),
		.out_wire_0_1(horizontal_tile_0_22_to_tile_0_23_1),
		.out_wire_0_2(horizontal_tile_0_22_to_tile_0_23_2),
		.out_wire_0_3(horizontal_tile_0_22_to_tile_0_23_3),
		.in_wire_0_0(horizontal_tile_0_23_to_tile_0_22_0),
		.in_wire_0_1(horizontal_tile_0_23_to_tile_0_22_1),
		.in_wire_0_2(horizontal_tile_0_23_to_tile_0_22_2),
		.in_wire_0_3(horizontal_tile_0_23_to_tile_0_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(23)
	);

	pe_tile_top pe_tile_0_23(
		.in_wire_3_0(input_to_grid_23),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_23_to_tile_1_23_0),
		.out_wire_1_1(vertical_tile_0_23_to_tile_1_23_1),
		.out_wire_1_2(vertical_tile_0_23_to_tile_1_23_2),
		.out_wire_1_3(vertical_tile_0_23_to_tile_1_23_3),
		.in_wire_1_0(vertical_tile_1_23_to_tile_0_23_0),
		.in_wire_1_1(vertical_tile_1_23_to_tile_0_23_1),
		.in_wire_1_2(vertical_tile_1_23_to_tile_0_23_2),
		.in_wire_1_3(vertical_tile_1_23_to_tile_0_23_3),
		.out_wire_2_0(horizontal_tile_0_23_to_tile_0_22_0),
		.out_wire_2_1(horizontal_tile_0_23_to_tile_0_22_1),
		.out_wire_2_2(horizontal_tile_0_23_to_tile_0_22_2),
		.out_wire_2_3(horizontal_tile_0_23_to_tile_0_22_3),
		.in_wire_2_0(horizontal_tile_0_22_to_tile_0_23_0),
		.in_wire_2_1(horizontal_tile_0_22_to_tile_0_23_1),
		.in_wire_2_2(horizontal_tile_0_22_to_tile_0_23_2),
		.in_wire_2_3(horizontal_tile_0_22_to_tile_0_23_3),
		.out_wire_0_0(horizontal_tile_0_23_to_tile_0_24_0),
		.out_wire_0_1(horizontal_tile_0_23_to_tile_0_24_1),
		.out_wire_0_2(horizontal_tile_0_23_to_tile_0_24_2),
		.out_wire_0_3(horizontal_tile_0_23_to_tile_0_24_3),
		.in_wire_0_0(horizontal_tile_0_24_to_tile_0_23_0),
		.in_wire_0_1(horizontal_tile_0_24_to_tile_0_23_1),
		.in_wire_0_2(horizontal_tile_0_24_to_tile_0_23_2),
		.in_wire_0_3(horizontal_tile_0_24_to_tile_0_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(24)
	);

	pe_tile_top pe_tile_0_24(
		.in_wire_3_0(input_to_grid_24),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_24_to_tile_1_24_0),
		.out_wire_1_1(vertical_tile_0_24_to_tile_1_24_1),
		.out_wire_1_2(vertical_tile_0_24_to_tile_1_24_2),
		.out_wire_1_3(vertical_tile_0_24_to_tile_1_24_3),
		.in_wire_1_0(vertical_tile_1_24_to_tile_0_24_0),
		.in_wire_1_1(vertical_tile_1_24_to_tile_0_24_1),
		.in_wire_1_2(vertical_tile_1_24_to_tile_0_24_2),
		.in_wire_1_3(vertical_tile_1_24_to_tile_0_24_3),
		.out_wire_2_0(horizontal_tile_0_24_to_tile_0_23_0),
		.out_wire_2_1(horizontal_tile_0_24_to_tile_0_23_1),
		.out_wire_2_2(horizontal_tile_0_24_to_tile_0_23_2),
		.out_wire_2_3(horizontal_tile_0_24_to_tile_0_23_3),
		.in_wire_2_0(horizontal_tile_0_23_to_tile_0_24_0),
		.in_wire_2_1(horizontal_tile_0_23_to_tile_0_24_1),
		.in_wire_2_2(horizontal_tile_0_23_to_tile_0_24_2),
		.in_wire_2_3(horizontal_tile_0_23_to_tile_0_24_3),
		.out_wire_0_0(horizontal_tile_0_24_to_tile_0_25_0),
		.out_wire_0_1(horizontal_tile_0_24_to_tile_0_25_1),
		.out_wire_0_2(horizontal_tile_0_24_to_tile_0_25_2),
		.out_wire_0_3(horizontal_tile_0_24_to_tile_0_25_3),
		.in_wire_0_0(horizontal_tile_0_25_to_tile_0_24_0),
		.in_wire_0_1(horizontal_tile_0_25_to_tile_0_24_1),
		.in_wire_0_2(horizontal_tile_0_25_to_tile_0_24_2),
		.in_wire_0_3(horizontal_tile_0_25_to_tile_0_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(25)
	);

	pe_tile_top pe_tile_0_25(
		.in_wire_3_0(input_to_grid_25),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_25_to_tile_1_25_0),
		.out_wire_1_1(vertical_tile_0_25_to_tile_1_25_1),
		.out_wire_1_2(vertical_tile_0_25_to_tile_1_25_2),
		.out_wire_1_3(vertical_tile_0_25_to_tile_1_25_3),
		.in_wire_1_0(vertical_tile_1_25_to_tile_0_25_0),
		.in_wire_1_1(vertical_tile_1_25_to_tile_0_25_1),
		.in_wire_1_2(vertical_tile_1_25_to_tile_0_25_2),
		.in_wire_1_3(vertical_tile_1_25_to_tile_0_25_3),
		.out_wire_2_0(horizontal_tile_0_25_to_tile_0_24_0),
		.out_wire_2_1(horizontal_tile_0_25_to_tile_0_24_1),
		.out_wire_2_2(horizontal_tile_0_25_to_tile_0_24_2),
		.out_wire_2_3(horizontal_tile_0_25_to_tile_0_24_3),
		.in_wire_2_0(horizontal_tile_0_24_to_tile_0_25_0),
		.in_wire_2_1(horizontal_tile_0_24_to_tile_0_25_1),
		.in_wire_2_2(horizontal_tile_0_24_to_tile_0_25_2),
		.in_wire_2_3(horizontal_tile_0_24_to_tile_0_25_3),
		.out_wire_0_0(horizontal_tile_0_25_to_tile_0_26_0),
		.out_wire_0_1(horizontal_tile_0_25_to_tile_0_26_1),
		.out_wire_0_2(horizontal_tile_0_25_to_tile_0_26_2),
		.out_wire_0_3(horizontal_tile_0_25_to_tile_0_26_3),
		.in_wire_0_0(horizontal_tile_0_26_to_tile_0_25_0),
		.in_wire_0_1(horizontal_tile_0_26_to_tile_0_25_1),
		.in_wire_0_2(horizontal_tile_0_26_to_tile_0_25_2),
		.in_wire_0_3(horizontal_tile_0_26_to_tile_0_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(26)
	);

	pe_tile_top pe_tile_0_26(
		.in_wire_3_0(input_to_grid_26),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_26_to_tile_1_26_0),
		.out_wire_1_1(vertical_tile_0_26_to_tile_1_26_1),
		.out_wire_1_2(vertical_tile_0_26_to_tile_1_26_2),
		.out_wire_1_3(vertical_tile_0_26_to_tile_1_26_3),
		.in_wire_1_0(vertical_tile_1_26_to_tile_0_26_0),
		.in_wire_1_1(vertical_tile_1_26_to_tile_0_26_1),
		.in_wire_1_2(vertical_tile_1_26_to_tile_0_26_2),
		.in_wire_1_3(vertical_tile_1_26_to_tile_0_26_3),
		.out_wire_2_0(horizontal_tile_0_26_to_tile_0_25_0),
		.out_wire_2_1(horizontal_tile_0_26_to_tile_0_25_1),
		.out_wire_2_2(horizontal_tile_0_26_to_tile_0_25_2),
		.out_wire_2_3(horizontal_tile_0_26_to_tile_0_25_3),
		.in_wire_2_0(horizontal_tile_0_25_to_tile_0_26_0),
		.in_wire_2_1(horizontal_tile_0_25_to_tile_0_26_1),
		.in_wire_2_2(horizontal_tile_0_25_to_tile_0_26_2),
		.in_wire_2_3(horizontal_tile_0_25_to_tile_0_26_3),
		.out_wire_0_0(horizontal_tile_0_26_to_tile_0_27_0),
		.out_wire_0_1(horizontal_tile_0_26_to_tile_0_27_1),
		.out_wire_0_2(horizontal_tile_0_26_to_tile_0_27_2),
		.out_wire_0_3(horizontal_tile_0_26_to_tile_0_27_3),
		.in_wire_0_0(horizontal_tile_0_27_to_tile_0_26_0),
		.in_wire_0_1(horizontal_tile_0_27_to_tile_0_26_1),
		.in_wire_0_2(horizontal_tile_0_27_to_tile_0_26_2),
		.in_wire_0_3(horizontal_tile_0_27_to_tile_0_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(27)
	);

	pe_tile_top pe_tile_0_27(
		.in_wire_3_0(input_to_grid_27),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_27_to_tile_1_27_0),
		.out_wire_1_1(vertical_tile_0_27_to_tile_1_27_1),
		.out_wire_1_2(vertical_tile_0_27_to_tile_1_27_2),
		.out_wire_1_3(vertical_tile_0_27_to_tile_1_27_3),
		.in_wire_1_0(vertical_tile_1_27_to_tile_0_27_0),
		.in_wire_1_1(vertical_tile_1_27_to_tile_0_27_1),
		.in_wire_1_2(vertical_tile_1_27_to_tile_0_27_2),
		.in_wire_1_3(vertical_tile_1_27_to_tile_0_27_3),
		.out_wire_2_0(horizontal_tile_0_27_to_tile_0_26_0),
		.out_wire_2_1(horizontal_tile_0_27_to_tile_0_26_1),
		.out_wire_2_2(horizontal_tile_0_27_to_tile_0_26_2),
		.out_wire_2_3(horizontal_tile_0_27_to_tile_0_26_3),
		.in_wire_2_0(horizontal_tile_0_26_to_tile_0_27_0),
		.in_wire_2_1(horizontal_tile_0_26_to_tile_0_27_1),
		.in_wire_2_2(horizontal_tile_0_26_to_tile_0_27_2),
		.in_wire_2_3(horizontal_tile_0_26_to_tile_0_27_3),
		.out_wire_0_0(horizontal_tile_0_27_to_tile_0_28_0),
		.out_wire_0_1(horizontal_tile_0_27_to_tile_0_28_1),
		.out_wire_0_2(horizontal_tile_0_27_to_tile_0_28_2),
		.out_wire_0_3(horizontal_tile_0_27_to_tile_0_28_3),
		.in_wire_0_0(horizontal_tile_0_28_to_tile_0_27_0),
		.in_wire_0_1(horizontal_tile_0_28_to_tile_0_27_1),
		.in_wire_0_2(horizontal_tile_0_28_to_tile_0_27_2),
		.in_wire_0_3(horizontal_tile_0_28_to_tile_0_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(28)
	);

	pe_tile_top pe_tile_0_28(
		.in_wire_3_0(input_to_grid_28),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_28_to_tile_1_28_0),
		.out_wire_1_1(vertical_tile_0_28_to_tile_1_28_1),
		.out_wire_1_2(vertical_tile_0_28_to_tile_1_28_2),
		.out_wire_1_3(vertical_tile_0_28_to_tile_1_28_3),
		.in_wire_1_0(vertical_tile_1_28_to_tile_0_28_0),
		.in_wire_1_1(vertical_tile_1_28_to_tile_0_28_1),
		.in_wire_1_2(vertical_tile_1_28_to_tile_0_28_2),
		.in_wire_1_3(vertical_tile_1_28_to_tile_0_28_3),
		.out_wire_2_0(horizontal_tile_0_28_to_tile_0_27_0),
		.out_wire_2_1(horizontal_tile_0_28_to_tile_0_27_1),
		.out_wire_2_2(horizontal_tile_0_28_to_tile_0_27_2),
		.out_wire_2_3(horizontal_tile_0_28_to_tile_0_27_3),
		.in_wire_2_0(horizontal_tile_0_27_to_tile_0_28_0),
		.in_wire_2_1(horizontal_tile_0_27_to_tile_0_28_1),
		.in_wire_2_2(horizontal_tile_0_27_to_tile_0_28_2),
		.in_wire_2_3(horizontal_tile_0_27_to_tile_0_28_3),
		.out_wire_0_0(horizontal_tile_0_28_to_tile_0_29_0),
		.out_wire_0_1(horizontal_tile_0_28_to_tile_0_29_1),
		.out_wire_0_2(horizontal_tile_0_28_to_tile_0_29_2),
		.out_wire_0_3(horizontal_tile_0_28_to_tile_0_29_3),
		.in_wire_0_0(horizontal_tile_0_29_to_tile_0_28_0),
		.in_wire_0_1(horizontal_tile_0_29_to_tile_0_28_1),
		.in_wire_0_2(horizontal_tile_0_29_to_tile_0_28_2),
		.in_wire_0_3(horizontal_tile_0_29_to_tile_0_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(29)
	);

	pe_tile_top pe_tile_0_29(
		.in_wire_3_0(input_to_grid_29),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_29_to_tile_1_29_0),
		.out_wire_1_1(vertical_tile_0_29_to_tile_1_29_1),
		.out_wire_1_2(vertical_tile_0_29_to_tile_1_29_2),
		.out_wire_1_3(vertical_tile_0_29_to_tile_1_29_3),
		.in_wire_1_0(vertical_tile_1_29_to_tile_0_29_0),
		.in_wire_1_1(vertical_tile_1_29_to_tile_0_29_1),
		.in_wire_1_2(vertical_tile_1_29_to_tile_0_29_2),
		.in_wire_1_3(vertical_tile_1_29_to_tile_0_29_3),
		.out_wire_2_0(horizontal_tile_0_29_to_tile_0_28_0),
		.out_wire_2_1(horizontal_tile_0_29_to_tile_0_28_1),
		.out_wire_2_2(horizontal_tile_0_29_to_tile_0_28_2),
		.out_wire_2_3(horizontal_tile_0_29_to_tile_0_28_3),
		.in_wire_2_0(horizontal_tile_0_28_to_tile_0_29_0),
		.in_wire_2_1(horizontal_tile_0_28_to_tile_0_29_1),
		.in_wire_2_2(horizontal_tile_0_28_to_tile_0_29_2),
		.in_wire_2_3(horizontal_tile_0_28_to_tile_0_29_3),
		.out_wire_0_0(horizontal_tile_0_29_to_tile_0_30_0),
		.out_wire_0_1(horizontal_tile_0_29_to_tile_0_30_1),
		.out_wire_0_2(horizontal_tile_0_29_to_tile_0_30_2),
		.out_wire_0_3(horizontal_tile_0_29_to_tile_0_30_3),
		.in_wire_0_0(horizontal_tile_0_30_to_tile_0_29_0),
		.in_wire_0_1(horizontal_tile_0_30_to_tile_0_29_1),
		.in_wire_0_2(horizontal_tile_0_30_to_tile_0_29_2),
		.in_wire_0_3(horizontal_tile_0_30_to_tile_0_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(30)
	);

	pe_tile_top pe_tile_0_30(
		.in_wire_3_0(input_to_grid_30),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_30_to_tile_1_30_0),
		.out_wire_1_1(vertical_tile_0_30_to_tile_1_30_1),
		.out_wire_1_2(vertical_tile_0_30_to_tile_1_30_2),
		.out_wire_1_3(vertical_tile_0_30_to_tile_1_30_3),
		.in_wire_1_0(vertical_tile_1_30_to_tile_0_30_0),
		.in_wire_1_1(vertical_tile_1_30_to_tile_0_30_1),
		.in_wire_1_2(vertical_tile_1_30_to_tile_0_30_2),
		.in_wire_1_3(vertical_tile_1_30_to_tile_0_30_3),
		.out_wire_2_0(horizontal_tile_0_30_to_tile_0_29_0),
		.out_wire_2_1(horizontal_tile_0_30_to_tile_0_29_1),
		.out_wire_2_2(horizontal_tile_0_30_to_tile_0_29_2),
		.out_wire_2_3(horizontal_tile_0_30_to_tile_0_29_3),
		.in_wire_2_0(horizontal_tile_0_29_to_tile_0_30_0),
		.in_wire_2_1(horizontal_tile_0_29_to_tile_0_30_1),
		.in_wire_2_2(horizontal_tile_0_29_to_tile_0_30_2),
		.in_wire_2_3(horizontal_tile_0_29_to_tile_0_30_3),
		.out_wire_0_0(horizontal_tile_0_30_to_tile_0_31_0),
		.out_wire_0_1(horizontal_tile_0_30_to_tile_0_31_1),
		.out_wire_0_2(horizontal_tile_0_30_to_tile_0_31_2),
		.out_wire_0_3(horizontal_tile_0_30_to_tile_0_31_3),
		.in_wire_0_0(horizontal_tile_0_31_to_tile_0_30_0),
		.in_wire_0_1(horizontal_tile_0_31_to_tile_0_30_1),
		.in_wire_0_2(horizontal_tile_0_31_to_tile_0_30_2),
		.in_wire_0_3(horizontal_tile_0_31_to_tile_0_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(31)
	);

	pe_tile_top_right pe_tile_0_31(
		.in_wire_3_0(input_to_grid_31),
		.in_wire_3_1(1'b0),
		.in_wire_3_2(1'b0),
		.in_wire_3_3(1'b0),
		.out_wire_1_0(vertical_tile_0_31_to_tile_1_31_0),
		.out_wire_1_1(vertical_tile_0_31_to_tile_1_31_1),
		.out_wire_1_2(vertical_tile_0_31_to_tile_1_31_2),
		.out_wire_1_3(vertical_tile_0_31_to_tile_1_31_3),
		.in_wire_1_0(vertical_tile_1_31_to_tile_0_31_0),
		.in_wire_1_1(vertical_tile_1_31_to_tile_0_31_1),
		.in_wire_1_2(vertical_tile_1_31_to_tile_0_31_2),
		.in_wire_1_3(vertical_tile_1_31_to_tile_0_31_3),
		.out_wire_2_0(horizontal_tile_0_31_to_tile_0_30_0),
		.out_wire_2_1(horizontal_tile_0_31_to_tile_0_30_1),
		.out_wire_2_2(horizontal_tile_0_31_to_tile_0_30_2),
		.out_wire_2_3(horizontal_tile_0_31_to_tile_0_30_3),
		.in_wire_2_0(horizontal_tile_0_30_to_tile_0_31_0),
		.in_wire_2_1(horizontal_tile_0_30_to_tile_0_31_1),
		.in_wire_2_2(horizontal_tile_0_30_to_tile_0_31_2),
		.in_wire_2_3(horizontal_tile_0_30_to_tile_0_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(32)
	);

	pe_tile_left pe_tile_1_0(
		.out_wire_3_0(vertical_tile_1_0_to_tile_0_0_0),
		.out_wire_3_1(vertical_tile_1_0_to_tile_0_0_1),
		.out_wire_3_2(vertical_tile_1_0_to_tile_0_0_2),
		.out_wire_3_3(vertical_tile_1_0_to_tile_0_0_3),
		.in_wire_3_0(vertical_tile_0_0_to_tile_1_0_0),
		.in_wire_3_1(vertical_tile_0_0_to_tile_1_0_1),
		.in_wire_3_2(vertical_tile_0_0_to_tile_1_0_2),
		.in_wire_3_3(vertical_tile_0_0_to_tile_1_0_3),
		.out_wire_1_0(vertical_tile_1_0_to_tile_2_0_0),
		.out_wire_1_1(vertical_tile_1_0_to_tile_2_0_1),
		.out_wire_1_2(vertical_tile_1_0_to_tile_2_0_2),
		.out_wire_1_3(vertical_tile_1_0_to_tile_2_0_3),
		.in_wire_1_0(vertical_tile_2_0_to_tile_1_0_0),
		.in_wire_1_1(vertical_tile_2_0_to_tile_1_0_1),
		.in_wire_1_2(vertical_tile_2_0_to_tile_1_0_2),
		.in_wire_1_3(vertical_tile_2_0_to_tile_1_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_1_0_to_tile_1_1_0),
		.out_wire_0_1(horizontal_tile_1_0_to_tile_1_1_1),
		.out_wire_0_2(horizontal_tile_1_0_to_tile_1_1_2),
		.out_wire_0_3(horizontal_tile_1_0_to_tile_1_1_3),
		.in_wire_0_0(horizontal_tile_1_1_to_tile_1_0_0),
		.in_wire_0_1(horizontal_tile_1_1_to_tile_1_0_1),
		.in_wire_0_2(horizontal_tile_1_1_to_tile_1_0_2),
		.in_wire_0_3(horizontal_tile_1_1_to_tile_1_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(33)
	);

	pe_tile pe_tile_1_1(
		.out_wire_3_0(vertical_tile_1_1_to_tile_0_1_0),
		.out_wire_3_1(vertical_tile_1_1_to_tile_0_1_1),
		.out_wire_3_2(vertical_tile_1_1_to_tile_0_1_2),
		.out_wire_3_3(vertical_tile_1_1_to_tile_0_1_3),
		.in_wire_3_0(vertical_tile_0_1_to_tile_1_1_0),
		.in_wire_3_1(vertical_tile_0_1_to_tile_1_1_1),
		.in_wire_3_2(vertical_tile_0_1_to_tile_1_1_2),
		.in_wire_3_3(vertical_tile_0_1_to_tile_1_1_3),
		.out_wire_1_0(vertical_tile_1_1_to_tile_2_1_0),
		.out_wire_1_1(vertical_tile_1_1_to_tile_2_1_1),
		.out_wire_1_2(vertical_tile_1_1_to_tile_2_1_2),
		.out_wire_1_3(vertical_tile_1_1_to_tile_2_1_3),
		.in_wire_1_0(vertical_tile_2_1_to_tile_1_1_0),
		.in_wire_1_1(vertical_tile_2_1_to_tile_1_1_1),
		.in_wire_1_2(vertical_tile_2_1_to_tile_1_1_2),
		.in_wire_1_3(vertical_tile_2_1_to_tile_1_1_3),
		.out_wire_2_0(horizontal_tile_1_1_to_tile_1_0_0),
		.out_wire_2_1(horizontal_tile_1_1_to_tile_1_0_1),
		.out_wire_2_2(horizontal_tile_1_1_to_tile_1_0_2),
		.out_wire_2_3(horizontal_tile_1_1_to_tile_1_0_3),
		.in_wire_2_0(horizontal_tile_1_0_to_tile_1_1_0),
		.in_wire_2_1(horizontal_tile_1_0_to_tile_1_1_1),
		.in_wire_2_2(horizontal_tile_1_0_to_tile_1_1_2),
		.in_wire_2_3(horizontal_tile_1_0_to_tile_1_1_3),
		.out_wire_0_0(horizontal_tile_1_1_to_tile_1_2_0),
		.out_wire_0_1(horizontal_tile_1_1_to_tile_1_2_1),
		.out_wire_0_2(horizontal_tile_1_1_to_tile_1_2_2),
		.out_wire_0_3(horizontal_tile_1_1_to_tile_1_2_3),
		.in_wire_0_0(horizontal_tile_1_2_to_tile_1_1_0),
		.in_wire_0_1(horizontal_tile_1_2_to_tile_1_1_1),
		.in_wire_0_2(horizontal_tile_1_2_to_tile_1_1_2),
		.in_wire_0_3(horizontal_tile_1_2_to_tile_1_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(34)
	);

	pe_tile pe_tile_1_2(
		.out_wire_3_0(vertical_tile_1_2_to_tile_0_2_0),
		.out_wire_3_1(vertical_tile_1_2_to_tile_0_2_1),
		.out_wire_3_2(vertical_tile_1_2_to_tile_0_2_2),
		.out_wire_3_3(vertical_tile_1_2_to_tile_0_2_3),
		.in_wire_3_0(vertical_tile_0_2_to_tile_1_2_0),
		.in_wire_3_1(vertical_tile_0_2_to_tile_1_2_1),
		.in_wire_3_2(vertical_tile_0_2_to_tile_1_2_2),
		.in_wire_3_3(vertical_tile_0_2_to_tile_1_2_3),
		.out_wire_1_0(vertical_tile_1_2_to_tile_2_2_0),
		.out_wire_1_1(vertical_tile_1_2_to_tile_2_2_1),
		.out_wire_1_2(vertical_tile_1_2_to_tile_2_2_2),
		.out_wire_1_3(vertical_tile_1_2_to_tile_2_2_3),
		.in_wire_1_0(vertical_tile_2_2_to_tile_1_2_0),
		.in_wire_1_1(vertical_tile_2_2_to_tile_1_2_1),
		.in_wire_1_2(vertical_tile_2_2_to_tile_1_2_2),
		.in_wire_1_3(vertical_tile_2_2_to_tile_1_2_3),
		.out_wire_2_0(horizontal_tile_1_2_to_tile_1_1_0),
		.out_wire_2_1(horizontal_tile_1_2_to_tile_1_1_1),
		.out_wire_2_2(horizontal_tile_1_2_to_tile_1_1_2),
		.out_wire_2_3(horizontal_tile_1_2_to_tile_1_1_3),
		.in_wire_2_0(horizontal_tile_1_1_to_tile_1_2_0),
		.in_wire_2_1(horizontal_tile_1_1_to_tile_1_2_1),
		.in_wire_2_2(horizontal_tile_1_1_to_tile_1_2_2),
		.in_wire_2_3(horizontal_tile_1_1_to_tile_1_2_3),
		.out_wire_0_0(horizontal_tile_1_2_to_tile_1_3_0),
		.out_wire_0_1(horizontal_tile_1_2_to_tile_1_3_1),
		.out_wire_0_2(horizontal_tile_1_2_to_tile_1_3_2),
		.out_wire_0_3(horizontal_tile_1_2_to_tile_1_3_3),
		.in_wire_0_0(horizontal_tile_1_3_to_tile_1_2_0),
		.in_wire_0_1(horizontal_tile_1_3_to_tile_1_2_1),
		.in_wire_0_2(horizontal_tile_1_3_to_tile_1_2_2),
		.in_wire_0_3(horizontal_tile_1_3_to_tile_1_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(35)
	);

	pe_tile pe_tile_1_3(
		.out_wire_3_0(vertical_tile_1_3_to_tile_0_3_0),
		.out_wire_3_1(vertical_tile_1_3_to_tile_0_3_1),
		.out_wire_3_2(vertical_tile_1_3_to_tile_0_3_2),
		.out_wire_3_3(vertical_tile_1_3_to_tile_0_3_3),
		.in_wire_3_0(vertical_tile_0_3_to_tile_1_3_0),
		.in_wire_3_1(vertical_tile_0_3_to_tile_1_3_1),
		.in_wire_3_2(vertical_tile_0_3_to_tile_1_3_2),
		.in_wire_3_3(vertical_tile_0_3_to_tile_1_3_3),
		.out_wire_1_0(vertical_tile_1_3_to_tile_2_3_0),
		.out_wire_1_1(vertical_tile_1_3_to_tile_2_3_1),
		.out_wire_1_2(vertical_tile_1_3_to_tile_2_3_2),
		.out_wire_1_3(vertical_tile_1_3_to_tile_2_3_3),
		.in_wire_1_0(vertical_tile_2_3_to_tile_1_3_0),
		.in_wire_1_1(vertical_tile_2_3_to_tile_1_3_1),
		.in_wire_1_2(vertical_tile_2_3_to_tile_1_3_2),
		.in_wire_1_3(vertical_tile_2_3_to_tile_1_3_3),
		.out_wire_2_0(horizontal_tile_1_3_to_tile_1_2_0),
		.out_wire_2_1(horizontal_tile_1_3_to_tile_1_2_1),
		.out_wire_2_2(horizontal_tile_1_3_to_tile_1_2_2),
		.out_wire_2_3(horizontal_tile_1_3_to_tile_1_2_3),
		.in_wire_2_0(horizontal_tile_1_2_to_tile_1_3_0),
		.in_wire_2_1(horizontal_tile_1_2_to_tile_1_3_1),
		.in_wire_2_2(horizontal_tile_1_2_to_tile_1_3_2),
		.in_wire_2_3(horizontal_tile_1_2_to_tile_1_3_3),
		.out_wire_0_0(horizontal_tile_1_3_to_tile_1_4_0),
		.out_wire_0_1(horizontal_tile_1_3_to_tile_1_4_1),
		.out_wire_0_2(horizontal_tile_1_3_to_tile_1_4_2),
		.out_wire_0_3(horizontal_tile_1_3_to_tile_1_4_3),
		.in_wire_0_0(horizontal_tile_1_4_to_tile_1_3_0),
		.in_wire_0_1(horizontal_tile_1_4_to_tile_1_3_1),
		.in_wire_0_2(horizontal_tile_1_4_to_tile_1_3_2),
		.in_wire_0_3(horizontal_tile_1_4_to_tile_1_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(36)
	);

	pe_tile pe_tile_1_4(
		.out_wire_3_0(vertical_tile_1_4_to_tile_0_4_0),
		.out_wire_3_1(vertical_tile_1_4_to_tile_0_4_1),
		.out_wire_3_2(vertical_tile_1_4_to_tile_0_4_2),
		.out_wire_3_3(vertical_tile_1_4_to_tile_0_4_3),
		.in_wire_3_0(vertical_tile_0_4_to_tile_1_4_0),
		.in_wire_3_1(vertical_tile_0_4_to_tile_1_4_1),
		.in_wire_3_2(vertical_tile_0_4_to_tile_1_4_2),
		.in_wire_3_3(vertical_tile_0_4_to_tile_1_4_3),
		.out_wire_1_0(vertical_tile_1_4_to_tile_2_4_0),
		.out_wire_1_1(vertical_tile_1_4_to_tile_2_4_1),
		.out_wire_1_2(vertical_tile_1_4_to_tile_2_4_2),
		.out_wire_1_3(vertical_tile_1_4_to_tile_2_4_3),
		.in_wire_1_0(vertical_tile_2_4_to_tile_1_4_0),
		.in_wire_1_1(vertical_tile_2_4_to_tile_1_4_1),
		.in_wire_1_2(vertical_tile_2_4_to_tile_1_4_2),
		.in_wire_1_3(vertical_tile_2_4_to_tile_1_4_3),
		.out_wire_2_0(horizontal_tile_1_4_to_tile_1_3_0),
		.out_wire_2_1(horizontal_tile_1_4_to_tile_1_3_1),
		.out_wire_2_2(horizontal_tile_1_4_to_tile_1_3_2),
		.out_wire_2_3(horizontal_tile_1_4_to_tile_1_3_3),
		.in_wire_2_0(horizontal_tile_1_3_to_tile_1_4_0),
		.in_wire_2_1(horizontal_tile_1_3_to_tile_1_4_1),
		.in_wire_2_2(horizontal_tile_1_3_to_tile_1_4_2),
		.in_wire_2_3(horizontal_tile_1_3_to_tile_1_4_3),
		.out_wire_0_0(horizontal_tile_1_4_to_tile_1_5_0),
		.out_wire_0_1(horizontal_tile_1_4_to_tile_1_5_1),
		.out_wire_0_2(horizontal_tile_1_4_to_tile_1_5_2),
		.out_wire_0_3(horizontal_tile_1_4_to_tile_1_5_3),
		.in_wire_0_0(horizontal_tile_1_5_to_tile_1_4_0),
		.in_wire_0_1(horizontal_tile_1_5_to_tile_1_4_1),
		.in_wire_0_2(horizontal_tile_1_5_to_tile_1_4_2),
		.in_wire_0_3(horizontal_tile_1_5_to_tile_1_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(37)
	);

	pe_tile pe_tile_1_5(
		.out_wire_3_0(vertical_tile_1_5_to_tile_0_5_0),
		.out_wire_3_1(vertical_tile_1_5_to_tile_0_5_1),
		.out_wire_3_2(vertical_tile_1_5_to_tile_0_5_2),
		.out_wire_3_3(vertical_tile_1_5_to_tile_0_5_3),
		.in_wire_3_0(vertical_tile_0_5_to_tile_1_5_0),
		.in_wire_3_1(vertical_tile_0_5_to_tile_1_5_1),
		.in_wire_3_2(vertical_tile_0_5_to_tile_1_5_2),
		.in_wire_3_3(vertical_tile_0_5_to_tile_1_5_3),
		.out_wire_1_0(vertical_tile_1_5_to_tile_2_5_0),
		.out_wire_1_1(vertical_tile_1_5_to_tile_2_5_1),
		.out_wire_1_2(vertical_tile_1_5_to_tile_2_5_2),
		.out_wire_1_3(vertical_tile_1_5_to_tile_2_5_3),
		.in_wire_1_0(vertical_tile_2_5_to_tile_1_5_0),
		.in_wire_1_1(vertical_tile_2_5_to_tile_1_5_1),
		.in_wire_1_2(vertical_tile_2_5_to_tile_1_5_2),
		.in_wire_1_3(vertical_tile_2_5_to_tile_1_5_3),
		.out_wire_2_0(horizontal_tile_1_5_to_tile_1_4_0),
		.out_wire_2_1(horizontal_tile_1_5_to_tile_1_4_1),
		.out_wire_2_2(horizontal_tile_1_5_to_tile_1_4_2),
		.out_wire_2_3(horizontal_tile_1_5_to_tile_1_4_3),
		.in_wire_2_0(horizontal_tile_1_4_to_tile_1_5_0),
		.in_wire_2_1(horizontal_tile_1_4_to_tile_1_5_1),
		.in_wire_2_2(horizontal_tile_1_4_to_tile_1_5_2),
		.in_wire_2_3(horizontal_tile_1_4_to_tile_1_5_3),
		.out_wire_0_0(horizontal_tile_1_5_to_tile_1_6_0),
		.out_wire_0_1(horizontal_tile_1_5_to_tile_1_6_1),
		.out_wire_0_2(horizontal_tile_1_5_to_tile_1_6_2),
		.out_wire_0_3(horizontal_tile_1_5_to_tile_1_6_3),
		.in_wire_0_0(horizontal_tile_1_6_to_tile_1_5_0),
		.in_wire_0_1(horizontal_tile_1_6_to_tile_1_5_1),
		.in_wire_0_2(horizontal_tile_1_6_to_tile_1_5_2),
		.in_wire_0_3(horizontal_tile_1_6_to_tile_1_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(38)
	);

	pe_tile pe_tile_1_6(
		.out_wire_3_0(vertical_tile_1_6_to_tile_0_6_0),
		.out_wire_3_1(vertical_tile_1_6_to_tile_0_6_1),
		.out_wire_3_2(vertical_tile_1_6_to_tile_0_6_2),
		.out_wire_3_3(vertical_tile_1_6_to_tile_0_6_3),
		.in_wire_3_0(vertical_tile_0_6_to_tile_1_6_0),
		.in_wire_3_1(vertical_tile_0_6_to_tile_1_6_1),
		.in_wire_3_2(vertical_tile_0_6_to_tile_1_6_2),
		.in_wire_3_3(vertical_tile_0_6_to_tile_1_6_3),
		.out_wire_1_0(vertical_tile_1_6_to_tile_2_6_0),
		.out_wire_1_1(vertical_tile_1_6_to_tile_2_6_1),
		.out_wire_1_2(vertical_tile_1_6_to_tile_2_6_2),
		.out_wire_1_3(vertical_tile_1_6_to_tile_2_6_3),
		.in_wire_1_0(vertical_tile_2_6_to_tile_1_6_0),
		.in_wire_1_1(vertical_tile_2_6_to_tile_1_6_1),
		.in_wire_1_2(vertical_tile_2_6_to_tile_1_6_2),
		.in_wire_1_3(vertical_tile_2_6_to_tile_1_6_3),
		.out_wire_2_0(horizontal_tile_1_6_to_tile_1_5_0),
		.out_wire_2_1(horizontal_tile_1_6_to_tile_1_5_1),
		.out_wire_2_2(horizontal_tile_1_6_to_tile_1_5_2),
		.out_wire_2_3(horizontal_tile_1_6_to_tile_1_5_3),
		.in_wire_2_0(horizontal_tile_1_5_to_tile_1_6_0),
		.in_wire_2_1(horizontal_tile_1_5_to_tile_1_6_1),
		.in_wire_2_2(horizontal_tile_1_5_to_tile_1_6_2),
		.in_wire_2_3(horizontal_tile_1_5_to_tile_1_6_3),
		.out_wire_0_0(horizontal_tile_1_6_to_tile_1_7_0),
		.out_wire_0_1(horizontal_tile_1_6_to_tile_1_7_1),
		.out_wire_0_2(horizontal_tile_1_6_to_tile_1_7_2),
		.out_wire_0_3(horizontal_tile_1_6_to_tile_1_7_3),
		.in_wire_0_0(horizontal_tile_1_7_to_tile_1_6_0),
		.in_wire_0_1(horizontal_tile_1_7_to_tile_1_6_1),
		.in_wire_0_2(horizontal_tile_1_7_to_tile_1_6_2),
		.in_wire_0_3(horizontal_tile_1_7_to_tile_1_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(39)
	);

	pe_tile pe_tile_1_7(
		.out_wire_3_0(vertical_tile_1_7_to_tile_0_7_0),
		.out_wire_3_1(vertical_tile_1_7_to_tile_0_7_1),
		.out_wire_3_2(vertical_tile_1_7_to_tile_0_7_2),
		.out_wire_3_3(vertical_tile_1_7_to_tile_0_7_3),
		.in_wire_3_0(vertical_tile_0_7_to_tile_1_7_0),
		.in_wire_3_1(vertical_tile_0_7_to_tile_1_7_1),
		.in_wire_3_2(vertical_tile_0_7_to_tile_1_7_2),
		.in_wire_3_3(vertical_tile_0_7_to_tile_1_7_3),
		.out_wire_1_0(vertical_tile_1_7_to_tile_2_7_0),
		.out_wire_1_1(vertical_tile_1_7_to_tile_2_7_1),
		.out_wire_1_2(vertical_tile_1_7_to_tile_2_7_2),
		.out_wire_1_3(vertical_tile_1_7_to_tile_2_7_3),
		.in_wire_1_0(vertical_tile_2_7_to_tile_1_7_0),
		.in_wire_1_1(vertical_tile_2_7_to_tile_1_7_1),
		.in_wire_1_2(vertical_tile_2_7_to_tile_1_7_2),
		.in_wire_1_3(vertical_tile_2_7_to_tile_1_7_3),
		.out_wire_2_0(horizontal_tile_1_7_to_tile_1_6_0),
		.out_wire_2_1(horizontal_tile_1_7_to_tile_1_6_1),
		.out_wire_2_2(horizontal_tile_1_7_to_tile_1_6_2),
		.out_wire_2_3(horizontal_tile_1_7_to_tile_1_6_3),
		.in_wire_2_0(horizontal_tile_1_6_to_tile_1_7_0),
		.in_wire_2_1(horizontal_tile_1_6_to_tile_1_7_1),
		.in_wire_2_2(horizontal_tile_1_6_to_tile_1_7_2),
		.in_wire_2_3(horizontal_tile_1_6_to_tile_1_7_3),
		.out_wire_0_0(horizontal_tile_1_7_to_tile_1_8_0),
		.out_wire_0_1(horizontal_tile_1_7_to_tile_1_8_1),
		.out_wire_0_2(horizontal_tile_1_7_to_tile_1_8_2),
		.out_wire_0_3(horizontal_tile_1_7_to_tile_1_8_3),
		.in_wire_0_0(horizontal_tile_1_8_to_tile_1_7_0),
		.in_wire_0_1(horizontal_tile_1_8_to_tile_1_7_1),
		.in_wire_0_2(horizontal_tile_1_8_to_tile_1_7_2),
		.in_wire_0_3(horizontal_tile_1_8_to_tile_1_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(40)
	);

	pe_tile pe_tile_1_8(
		.out_wire_3_0(vertical_tile_1_8_to_tile_0_8_0),
		.out_wire_3_1(vertical_tile_1_8_to_tile_0_8_1),
		.out_wire_3_2(vertical_tile_1_8_to_tile_0_8_2),
		.out_wire_3_3(vertical_tile_1_8_to_tile_0_8_3),
		.in_wire_3_0(vertical_tile_0_8_to_tile_1_8_0),
		.in_wire_3_1(vertical_tile_0_8_to_tile_1_8_1),
		.in_wire_3_2(vertical_tile_0_8_to_tile_1_8_2),
		.in_wire_3_3(vertical_tile_0_8_to_tile_1_8_3),
		.out_wire_1_0(vertical_tile_1_8_to_tile_2_8_0),
		.out_wire_1_1(vertical_tile_1_8_to_tile_2_8_1),
		.out_wire_1_2(vertical_tile_1_8_to_tile_2_8_2),
		.out_wire_1_3(vertical_tile_1_8_to_tile_2_8_3),
		.in_wire_1_0(vertical_tile_2_8_to_tile_1_8_0),
		.in_wire_1_1(vertical_tile_2_8_to_tile_1_8_1),
		.in_wire_1_2(vertical_tile_2_8_to_tile_1_8_2),
		.in_wire_1_3(vertical_tile_2_8_to_tile_1_8_3),
		.out_wire_2_0(horizontal_tile_1_8_to_tile_1_7_0),
		.out_wire_2_1(horizontal_tile_1_8_to_tile_1_7_1),
		.out_wire_2_2(horizontal_tile_1_8_to_tile_1_7_2),
		.out_wire_2_3(horizontal_tile_1_8_to_tile_1_7_3),
		.in_wire_2_0(horizontal_tile_1_7_to_tile_1_8_0),
		.in_wire_2_1(horizontal_tile_1_7_to_tile_1_8_1),
		.in_wire_2_2(horizontal_tile_1_7_to_tile_1_8_2),
		.in_wire_2_3(horizontal_tile_1_7_to_tile_1_8_3),
		.out_wire_0_0(horizontal_tile_1_8_to_tile_1_9_0),
		.out_wire_0_1(horizontal_tile_1_8_to_tile_1_9_1),
		.out_wire_0_2(horizontal_tile_1_8_to_tile_1_9_2),
		.out_wire_0_3(horizontal_tile_1_8_to_tile_1_9_3),
		.in_wire_0_0(horizontal_tile_1_9_to_tile_1_8_0),
		.in_wire_0_1(horizontal_tile_1_9_to_tile_1_8_1),
		.in_wire_0_2(horizontal_tile_1_9_to_tile_1_8_2),
		.in_wire_0_3(horizontal_tile_1_9_to_tile_1_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(41)
	);

	pe_tile pe_tile_1_9(
		.out_wire_3_0(vertical_tile_1_9_to_tile_0_9_0),
		.out_wire_3_1(vertical_tile_1_9_to_tile_0_9_1),
		.out_wire_3_2(vertical_tile_1_9_to_tile_0_9_2),
		.out_wire_3_3(vertical_tile_1_9_to_tile_0_9_3),
		.in_wire_3_0(vertical_tile_0_9_to_tile_1_9_0),
		.in_wire_3_1(vertical_tile_0_9_to_tile_1_9_1),
		.in_wire_3_2(vertical_tile_0_9_to_tile_1_9_2),
		.in_wire_3_3(vertical_tile_0_9_to_tile_1_9_3),
		.out_wire_1_0(vertical_tile_1_9_to_tile_2_9_0),
		.out_wire_1_1(vertical_tile_1_9_to_tile_2_9_1),
		.out_wire_1_2(vertical_tile_1_9_to_tile_2_9_2),
		.out_wire_1_3(vertical_tile_1_9_to_tile_2_9_3),
		.in_wire_1_0(vertical_tile_2_9_to_tile_1_9_0),
		.in_wire_1_1(vertical_tile_2_9_to_tile_1_9_1),
		.in_wire_1_2(vertical_tile_2_9_to_tile_1_9_2),
		.in_wire_1_3(vertical_tile_2_9_to_tile_1_9_3),
		.out_wire_2_0(horizontal_tile_1_9_to_tile_1_8_0),
		.out_wire_2_1(horizontal_tile_1_9_to_tile_1_8_1),
		.out_wire_2_2(horizontal_tile_1_9_to_tile_1_8_2),
		.out_wire_2_3(horizontal_tile_1_9_to_tile_1_8_3),
		.in_wire_2_0(horizontal_tile_1_8_to_tile_1_9_0),
		.in_wire_2_1(horizontal_tile_1_8_to_tile_1_9_1),
		.in_wire_2_2(horizontal_tile_1_8_to_tile_1_9_2),
		.in_wire_2_3(horizontal_tile_1_8_to_tile_1_9_3),
		.out_wire_0_0(horizontal_tile_1_9_to_tile_1_10_0),
		.out_wire_0_1(horizontal_tile_1_9_to_tile_1_10_1),
		.out_wire_0_2(horizontal_tile_1_9_to_tile_1_10_2),
		.out_wire_0_3(horizontal_tile_1_9_to_tile_1_10_3),
		.in_wire_0_0(horizontal_tile_1_10_to_tile_1_9_0),
		.in_wire_0_1(horizontal_tile_1_10_to_tile_1_9_1),
		.in_wire_0_2(horizontal_tile_1_10_to_tile_1_9_2),
		.in_wire_0_3(horizontal_tile_1_10_to_tile_1_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(42)
	);

	pe_tile pe_tile_1_10(
		.out_wire_3_0(vertical_tile_1_10_to_tile_0_10_0),
		.out_wire_3_1(vertical_tile_1_10_to_tile_0_10_1),
		.out_wire_3_2(vertical_tile_1_10_to_tile_0_10_2),
		.out_wire_3_3(vertical_tile_1_10_to_tile_0_10_3),
		.in_wire_3_0(vertical_tile_0_10_to_tile_1_10_0),
		.in_wire_3_1(vertical_tile_0_10_to_tile_1_10_1),
		.in_wire_3_2(vertical_tile_0_10_to_tile_1_10_2),
		.in_wire_3_3(vertical_tile_0_10_to_tile_1_10_3),
		.out_wire_1_0(vertical_tile_1_10_to_tile_2_10_0),
		.out_wire_1_1(vertical_tile_1_10_to_tile_2_10_1),
		.out_wire_1_2(vertical_tile_1_10_to_tile_2_10_2),
		.out_wire_1_3(vertical_tile_1_10_to_tile_2_10_3),
		.in_wire_1_0(vertical_tile_2_10_to_tile_1_10_0),
		.in_wire_1_1(vertical_tile_2_10_to_tile_1_10_1),
		.in_wire_1_2(vertical_tile_2_10_to_tile_1_10_2),
		.in_wire_1_3(vertical_tile_2_10_to_tile_1_10_3),
		.out_wire_2_0(horizontal_tile_1_10_to_tile_1_9_0),
		.out_wire_2_1(horizontal_tile_1_10_to_tile_1_9_1),
		.out_wire_2_2(horizontal_tile_1_10_to_tile_1_9_2),
		.out_wire_2_3(horizontal_tile_1_10_to_tile_1_9_3),
		.in_wire_2_0(horizontal_tile_1_9_to_tile_1_10_0),
		.in_wire_2_1(horizontal_tile_1_9_to_tile_1_10_1),
		.in_wire_2_2(horizontal_tile_1_9_to_tile_1_10_2),
		.in_wire_2_3(horizontal_tile_1_9_to_tile_1_10_3),
		.out_wire_0_0(horizontal_tile_1_10_to_tile_1_11_0),
		.out_wire_0_1(horizontal_tile_1_10_to_tile_1_11_1),
		.out_wire_0_2(horizontal_tile_1_10_to_tile_1_11_2),
		.out_wire_0_3(horizontal_tile_1_10_to_tile_1_11_3),
		.in_wire_0_0(horizontal_tile_1_11_to_tile_1_10_0),
		.in_wire_0_1(horizontal_tile_1_11_to_tile_1_10_1),
		.in_wire_0_2(horizontal_tile_1_11_to_tile_1_10_2),
		.in_wire_0_3(horizontal_tile_1_11_to_tile_1_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(43)
	);

	pe_tile pe_tile_1_11(
		.out_wire_3_0(vertical_tile_1_11_to_tile_0_11_0),
		.out_wire_3_1(vertical_tile_1_11_to_tile_0_11_1),
		.out_wire_3_2(vertical_tile_1_11_to_tile_0_11_2),
		.out_wire_3_3(vertical_tile_1_11_to_tile_0_11_3),
		.in_wire_3_0(vertical_tile_0_11_to_tile_1_11_0),
		.in_wire_3_1(vertical_tile_0_11_to_tile_1_11_1),
		.in_wire_3_2(vertical_tile_0_11_to_tile_1_11_2),
		.in_wire_3_3(vertical_tile_0_11_to_tile_1_11_3),
		.out_wire_1_0(vertical_tile_1_11_to_tile_2_11_0),
		.out_wire_1_1(vertical_tile_1_11_to_tile_2_11_1),
		.out_wire_1_2(vertical_tile_1_11_to_tile_2_11_2),
		.out_wire_1_3(vertical_tile_1_11_to_tile_2_11_3),
		.in_wire_1_0(vertical_tile_2_11_to_tile_1_11_0),
		.in_wire_1_1(vertical_tile_2_11_to_tile_1_11_1),
		.in_wire_1_2(vertical_tile_2_11_to_tile_1_11_2),
		.in_wire_1_3(vertical_tile_2_11_to_tile_1_11_3),
		.out_wire_2_0(horizontal_tile_1_11_to_tile_1_10_0),
		.out_wire_2_1(horizontal_tile_1_11_to_tile_1_10_1),
		.out_wire_2_2(horizontal_tile_1_11_to_tile_1_10_2),
		.out_wire_2_3(horizontal_tile_1_11_to_tile_1_10_3),
		.in_wire_2_0(horizontal_tile_1_10_to_tile_1_11_0),
		.in_wire_2_1(horizontal_tile_1_10_to_tile_1_11_1),
		.in_wire_2_2(horizontal_tile_1_10_to_tile_1_11_2),
		.in_wire_2_3(horizontal_tile_1_10_to_tile_1_11_3),
		.out_wire_0_0(horizontal_tile_1_11_to_tile_1_12_0),
		.out_wire_0_1(horizontal_tile_1_11_to_tile_1_12_1),
		.out_wire_0_2(horizontal_tile_1_11_to_tile_1_12_2),
		.out_wire_0_3(horizontal_tile_1_11_to_tile_1_12_3),
		.in_wire_0_0(horizontal_tile_1_12_to_tile_1_11_0),
		.in_wire_0_1(horizontal_tile_1_12_to_tile_1_11_1),
		.in_wire_0_2(horizontal_tile_1_12_to_tile_1_11_2),
		.in_wire_0_3(horizontal_tile_1_12_to_tile_1_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(44)
	);

	pe_tile pe_tile_1_12(
		.out_wire_3_0(vertical_tile_1_12_to_tile_0_12_0),
		.out_wire_3_1(vertical_tile_1_12_to_tile_0_12_1),
		.out_wire_3_2(vertical_tile_1_12_to_tile_0_12_2),
		.out_wire_3_3(vertical_tile_1_12_to_tile_0_12_3),
		.in_wire_3_0(vertical_tile_0_12_to_tile_1_12_0),
		.in_wire_3_1(vertical_tile_0_12_to_tile_1_12_1),
		.in_wire_3_2(vertical_tile_0_12_to_tile_1_12_2),
		.in_wire_3_3(vertical_tile_0_12_to_tile_1_12_3),
		.out_wire_1_0(vertical_tile_1_12_to_tile_2_12_0),
		.out_wire_1_1(vertical_tile_1_12_to_tile_2_12_1),
		.out_wire_1_2(vertical_tile_1_12_to_tile_2_12_2),
		.out_wire_1_3(vertical_tile_1_12_to_tile_2_12_3),
		.in_wire_1_0(vertical_tile_2_12_to_tile_1_12_0),
		.in_wire_1_1(vertical_tile_2_12_to_tile_1_12_1),
		.in_wire_1_2(vertical_tile_2_12_to_tile_1_12_2),
		.in_wire_1_3(vertical_tile_2_12_to_tile_1_12_3),
		.out_wire_2_0(horizontal_tile_1_12_to_tile_1_11_0),
		.out_wire_2_1(horizontal_tile_1_12_to_tile_1_11_1),
		.out_wire_2_2(horizontal_tile_1_12_to_tile_1_11_2),
		.out_wire_2_3(horizontal_tile_1_12_to_tile_1_11_3),
		.in_wire_2_0(horizontal_tile_1_11_to_tile_1_12_0),
		.in_wire_2_1(horizontal_tile_1_11_to_tile_1_12_1),
		.in_wire_2_2(horizontal_tile_1_11_to_tile_1_12_2),
		.in_wire_2_3(horizontal_tile_1_11_to_tile_1_12_3),
		.out_wire_0_0(horizontal_tile_1_12_to_tile_1_13_0),
		.out_wire_0_1(horizontal_tile_1_12_to_tile_1_13_1),
		.out_wire_0_2(horizontal_tile_1_12_to_tile_1_13_2),
		.out_wire_0_3(horizontal_tile_1_12_to_tile_1_13_3),
		.in_wire_0_0(horizontal_tile_1_13_to_tile_1_12_0),
		.in_wire_0_1(horizontal_tile_1_13_to_tile_1_12_1),
		.in_wire_0_2(horizontal_tile_1_13_to_tile_1_12_2),
		.in_wire_0_3(horizontal_tile_1_13_to_tile_1_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(45)
	);

	pe_tile pe_tile_1_13(
		.out_wire_3_0(vertical_tile_1_13_to_tile_0_13_0),
		.out_wire_3_1(vertical_tile_1_13_to_tile_0_13_1),
		.out_wire_3_2(vertical_tile_1_13_to_tile_0_13_2),
		.out_wire_3_3(vertical_tile_1_13_to_tile_0_13_3),
		.in_wire_3_0(vertical_tile_0_13_to_tile_1_13_0),
		.in_wire_3_1(vertical_tile_0_13_to_tile_1_13_1),
		.in_wire_3_2(vertical_tile_0_13_to_tile_1_13_2),
		.in_wire_3_3(vertical_tile_0_13_to_tile_1_13_3),
		.out_wire_1_0(vertical_tile_1_13_to_tile_2_13_0),
		.out_wire_1_1(vertical_tile_1_13_to_tile_2_13_1),
		.out_wire_1_2(vertical_tile_1_13_to_tile_2_13_2),
		.out_wire_1_3(vertical_tile_1_13_to_tile_2_13_3),
		.in_wire_1_0(vertical_tile_2_13_to_tile_1_13_0),
		.in_wire_1_1(vertical_tile_2_13_to_tile_1_13_1),
		.in_wire_1_2(vertical_tile_2_13_to_tile_1_13_2),
		.in_wire_1_3(vertical_tile_2_13_to_tile_1_13_3),
		.out_wire_2_0(horizontal_tile_1_13_to_tile_1_12_0),
		.out_wire_2_1(horizontal_tile_1_13_to_tile_1_12_1),
		.out_wire_2_2(horizontal_tile_1_13_to_tile_1_12_2),
		.out_wire_2_3(horizontal_tile_1_13_to_tile_1_12_3),
		.in_wire_2_0(horizontal_tile_1_12_to_tile_1_13_0),
		.in_wire_2_1(horizontal_tile_1_12_to_tile_1_13_1),
		.in_wire_2_2(horizontal_tile_1_12_to_tile_1_13_2),
		.in_wire_2_3(horizontal_tile_1_12_to_tile_1_13_3),
		.out_wire_0_0(horizontal_tile_1_13_to_tile_1_14_0),
		.out_wire_0_1(horizontal_tile_1_13_to_tile_1_14_1),
		.out_wire_0_2(horizontal_tile_1_13_to_tile_1_14_2),
		.out_wire_0_3(horizontal_tile_1_13_to_tile_1_14_3),
		.in_wire_0_0(horizontal_tile_1_14_to_tile_1_13_0),
		.in_wire_0_1(horizontal_tile_1_14_to_tile_1_13_1),
		.in_wire_0_2(horizontal_tile_1_14_to_tile_1_13_2),
		.in_wire_0_3(horizontal_tile_1_14_to_tile_1_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(46)
	);

	pe_tile pe_tile_1_14(
		.out_wire_3_0(vertical_tile_1_14_to_tile_0_14_0),
		.out_wire_3_1(vertical_tile_1_14_to_tile_0_14_1),
		.out_wire_3_2(vertical_tile_1_14_to_tile_0_14_2),
		.out_wire_3_3(vertical_tile_1_14_to_tile_0_14_3),
		.in_wire_3_0(vertical_tile_0_14_to_tile_1_14_0),
		.in_wire_3_1(vertical_tile_0_14_to_tile_1_14_1),
		.in_wire_3_2(vertical_tile_0_14_to_tile_1_14_2),
		.in_wire_3_3(vertical_tile_0_14_to_tile_1_14_3),
		.out_wire_1_0(vertical_tile_1_14_to_tile_2_14_0),
		.out_wire_1_1(vertical_tile_1_14_to_tile_2_14_1),
		.out_wire_1_2(vertical_tile_1_14_to_tile_2_14_2),
		.out_wire_1_3(vertical_tile_1_14_to_tile_2_14_3),
		.in_wire_1_0(vertical_tile_2_14_to_tile_1_14_0),
		.in_wire_1_1(vertical_tile_2_14_to_tile_1_14_1),
		.in_wire_1_2(vertical_tile_2_14_to_tile_1_14_2),
		.in_wire_1_3(vertical_tile_2_14_to_tile_1_14_3),
		.out_wire_2_0(horizontal_tile_1_14_to_tile_1_13_0),
		.out_wire_2_1(horizontal_tile_1_14_to_tile_1_13_1),
		.out_wire_2_2(horizontal_tile_1_14_to_tile_1_13_2),
		.out_wire_2_3(horizontal_tile_1_14_to_tile_1_13_3),
		.in_wire_2_0(horizontal_tile_1_13_to_tile_1_14_0),
		.in_wire_2_1(horizontal_tile_1_13_to_tile_1_14_1),
		.in_wire_2_2(horizontal_tile_1_13_to_tile_1_14_2),
		.in_wire_2_3(horizontal_tile_1_13_to_tile_1_14_3),
		.out_wire_0_0(horizontal_tile_1_14_to_tile_1_15_0),
		.out_wire_0_1(horizontal_tile_1_14_to_tile_1_15_1),
		.out_wire_0_2(horizontal_tile_1_14_to_tile_1_15_2),
		.out_wire_0_3(horizontal_tile_1_14_to_tile_1_15_3),
		.in_wire_0_0(horizontal_tile_1_15_to_tile_1_14_0),
		.in_wire_0_1(horizontal_tile_1_15_to_tile_1_14_1),
		.in_wire_0_2(horizontal_tile_1_15_to_tile_1_14_2),
		.in_wire_0_3(horizontal_tile_1_15_to_tile_1_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(47)
	);

	pe_tile pe_tile_1_15(
		.out_wire_3_0(vertical_tile_1_15_to_tile_0_15_0),
		.out_wire_3_1(vertical_tile_1_15_to_tile_0_15_1),
		.out_wire_3_2(vertical_tile_1_15_to_tile_0_15_2),
		.out_wire_3_3(vertical_tile_1_15_to_tile_0_15_3),
		.in_wire_3_0(vertical_tile_0_15_to_tile_1_15_0),
		.in_wire_3_1(vertical_tile_0_15_to_tile_1_15_1),
		.in_wire_3_2(vertical_tile_0_15_to_tile_1_15_2),
		.in_wire_3_3(vertical_tile_0_15_to_tile_1_15_3),
		.out_wire_1_0(vertical_tile_1_15_to_tile_2_15_0),
		.out_wire_1_1(vertical_tile_1_15_to_tile_2_15_1),
		.out_wire_1_2(vertical_tile_1_15_to_tile_2_15_2),
		.out_wire_1_3(vertical_tile_1_15_to_tile_2_15_3),
		.in_wire_1_0(vertical_tile_2_15_to_tile_1_15_0),
		.in_wire_1_1(vertical_tile_2_15_to_tile_1_15_1),
		.in_wire_1_2(vertical_tile_2_15_to_tile_1_15_2),
		.in_wire_1_3(vertical_tile_2_15_to_tile_1_15_3),
		.out_wire_2_0(horizontal_tile_1_15_to_tile_1_14_0),
		.out_wire_2_1(horizontal_tile_1_15_to_tile_1_14_1),
		.out_wire_2_2(horizontal_tile_1_15_to_tile_1_14_2),
		.out_wire_2_3(horizontal_tile_1_15_to_tile_1_14_3),
		.in_wire_2_0(horizontal_tile_1_14_to_tile_1_15_0),
		.in_wire_2_1(horizontal_tile_1_14_to_tile_1_15_1),
		.in_wire_2_2(horizontal_tile_1_14_to_tile_1_15_2),
		.in_wire_2_3(horizontal_tile_1_14_to_tile_1_15_3),
		.out_wire_0_0(horizontal_tile_1_15_to_tile_1_16_0),
		.out_wire_0_1(horizontal_tile_1_15_to_tile_1_16_1),
		.out_wire_0_2(horizontal_tile_1_15_to_tile_1_16_2),
		.out_wire_0_3(horizontal_tile_1_15_to_tile_1_16_3),
		.in_wire_0_0(horizontal_tile_1_16_to_tile_1_15_0),
		.in_wire_0_1(horizontal_tile_1_16_to_tile_1_15_1),
		.in_wire_0_2(horizontal_tile_1_16_to_tile_1_15_2),
		.in_wire_0_3(horizontal_tile_1_16_to_tile_1_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(48)
	);

	pe_tile pe_tile_1_16(
		.out_wire_3_0(vertical_tile_1_16_to_tile_0_16_0),
		.out_wire_3_1(vertical_tile_1_16_to_tile_0_16_1),
		.out_wire_3_2(vertical_tile_1_16_to_tile_0_16_2),
		.out_wire_3_3(vertical_tile_1_16_to_tile_0_16_3),
		.in_wire_3_0(vertical_tile_0_16_to_tile_1_16_0),
		.in_wire_3_1(vertical_tile_0_16_to_tile_1_16_1),
		.in_wire_3_2(vertical_tile_0_16_to_tile_1_16_2),
		.in_wire_3_3(vertical_tile_0_16_to_tile_1_16_3),
		.out_wire_1_0(vertical_tile_1_16_to_tile_2_16_0),
		.out_wire_1_1(vertical_tile_1_16_to_tile_2_16_1),
		.out_wire_1_2(vertical_tile_1_16_to_tile_2_16_2),
		.out_wire_1_3(vertical_tile_1_16_to_tile_2_16_3),
		.in_wire_1_0(vertical_tile_2_16_to_tile_1_16_0),
		.in_wire_1_1(vertical_tile_2_16_to_tile_1_16_1),
		.in_wire_1_2(vertical_tile_2_16_to_tile_1_16_2),
		.in_wire_1_3(vertical_tile_2_16_to_tile_1_16_3),
		.out_wire_2_0(horizontal_tile_1_16_to_tile_1_15_0),
		.out_wire_2_1(horizontal_tile_1_16_to_tile_1_15_1),
		.out_wire_2_2(horizontal_tile_1_16_to_tile_1_15_2),
		.out_wire_2_3(horizontal_tile_1_16_to_tile_1_15_3),
		.in_wire_2_0(horizontal_tile_1_15_to_tile_1_16_0),
		.in_wire_2_1(horizontal_tile_1_15_to_tile_1_16_1),
		.in_wire_2_2(horizontal_tile_1_15_to_tile_1_16_2),
		.in_wire_2_3(horizontal_tile_1_15_to_tile_1_16_3),
		.out_wire_0_0(horizontal_tile_1_16_to_tile_1_17_0),
		.out_wire_0_1(horizontal_tile_1_16_to_tile_1_17_1),
		.out_wire_0_2(horizontal_tile_1_16_to_tile_1_17_2),
		.out_wire_0_3(horizontal_tile_1_16_to_tile_1_17_3),
		.in_wire_0_0(horizontal_tile_1_17_to_tile_1_16_0),
		.in_wire_0_1(horizontal_tile_1_17_to_tile_1_16_1),
		.in_wire_0_2(horizontal_tile_1_17_to_tile_1_16_2),
		.in_wire_0_3(horizontal_tile_1_17_to_tile_1_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(49)
	);

	pe_tile pe_tile_1_17(
		.out_wire_3_0(vertical_tile_1_17_to_tile_0_17_0),
		.out_wire_3_1(vertical_tile_1_17_to_tile_0_17_1),
		.out_wire_3_2(vertical_tile_1_17_to_tile_0_17_2),
		.out_wire_3_3(vertical_tile_1_17_to_tile_0_17_3),
		.in_wire_3_0(vertical_tile_0_17_to_tile_1_17_0),
		.in_wire_3_1(vertical_tile_0_17_to_tile_1_17_1),
		.in_wire_3_2(vertical_tile_0_17_to_tile_1_17_2),
		.in_wire_3_3(vertical_tile_0_17_to_tile_1_17_3),
		.out_wire_1_0(vertical_tile_1_17_to_tile_2_17_0),
		.out_wire_1_1(vertical_tile_1_17_to_tile_2_17_1),
		.out_wire_1_2(vertical_tile_1_17_to_tile_2_17_2),
		.out_wire_1_3(vertical_tile_1_17_to_tile_2_17_3),
		.in_wire_1_0(vertical_tile_2_17_to_tile_1_17_0),
		.in_wire_1_1(vertical_tile_2_17_to_tile_1_17_1),
		.in_wire_1_2(vertical_tile_2_17_to_tile_1_17_2),
		.in_wire_1_3(vertical_tile_2_17_to_tile_1_17_3),
		.out_wire_2_0(horizontal_tile_1_17_to_tile_1_16_0),
		.out_wire_2_1(horizontal_tile_1_17_to_tile_1_16_1),
		.out_wire_2_2(horizontal_tile_1_17_to_tile_1_16_2),
		.out_wire_2_3(horizontal_tile_1_17_to_tile_1_16_3),
		.in_wire_2_0(horizontal_tile_1_16_to_tile_1_17_0),
		.in_wire_2_1(horizontal_tile_1_16_to_tile_1_17_1),
		.in_wire_2_2(horizontal_tile_1_16_to_tile_1_17_2),
		.in_wire_2_3(horizontal_tile_1_16_to_tile_1_17_3),
		.out_wire_0_0(horizontal_tile_1_17_to_tile_1_18_0),
		.out_wire_0_1(horizontal_tile_1_17_to_tile_1_18_1),
		.out_wire_0_2(horizontal_tile_1_17_to_tile_1_18_2),
		.out_wire_0_3(horizontal_tile_1_17_to_tile_1_18_3),
		.in_wire_0_0(horizontal_tile_1_18_to_tile_1_17_0),
		.in_wire_0_1(horizontal_tile_1_18_to_tile_1_17_1),
		.in_wire_0_2(horizontal_tile_1_18_to_tile_1_17_2),
		.in_wire_0_3(horizontal_tile_1_18_to_tile_1_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(50)
	);

	pe_tile pe_tile_1_18(
		.out_wire_3_0(vertical_tile_1_18_to_tile_0_18_0),
		.out_wire_3_1(vertical_tile_1_18_to_tile_0_18_1),
		.out_wire_3_2(vertical_tile_1_18_to_tile_0_18_2),
		.out_wire_3_3(vertical_tile_1_18_to_tile_0_18_3),
		.in_wire_3_0(vertical_tile_0_18_to_tile_1_18_0),
		.in_wire_3_1(vertical_tile_0_18_to_tile_1_18_1),
		.in_wire_3_2(vertical_tile_0_18_to_tile_1_18_2),
		.in_wire_3_3(vertical_tile_0_18_to_tile_1_18_3),
		.out_wire_1_0(vertical_tile_1_18_to_tile_2_18_0),
		.out_wire_1_1(vertical_tile_1_18_to_tile_2_18_1),
		.out_wire_1_2(vertical_tile_1_18_to_tile_2_18_2),
		.out_wire_1_3(vertical_tile_1_18_to_tile_2_18_3),
		.in_wire_1_0(vertical_tile_2_18_to_tile_1_18_0),
		.in_wire_1_1(vertical_tile_2_18_to_tile_1_18_1),
		.in_wire_1_2(vertical_tile_2_18_to_tile_1_18_2),
		.in_wire_1_3(vertical_tile_2_18_to_tile_1_18_3),
		.out_wire_2_0(horizontal_tile_1_18_to_tile_1_17_0),
		.out_wire_2_1(horizontal_tile_1_18_to_tile_1_17_1),
		.out_wire_2_2(horizontal_tile_1_18_to_tile_1_17_2),
		.out_wire_2_3(horizontal_tile_1_18_to_tile_1_17_3),
		.in_wire_2_0(horizontal_tile_1_17_to_tile_1_18_0),
		.in_wire_2_1(horizontal_tile_1_17_to_tile_1_18_1),
		.in_wire_2_2(horizontal_tile_1_17_to_tile_1_18_2),
		.in_wire_2_3(horizontal_tile_1_17_to_tile_1_18_3),
		.out_wire_0_0(horizontal_tile_1_18_to_tile_1_19_0),
		.out_wire_0_1(horizontal_tile_1_18_to_tile_1_19_1),
		.out_wire_0_2(horizontal_tile_1_18_to_tile_1_19_2),
		.out_wire_0_3(horizontal_tile_1_18_to_tile_1_19_3),
		.in_wire_0_0(horizontal_tile_1_19_to_tile_1_18_0),
		.in_wire_0_1(horizontal_tile_1_19_to_tile_1_18_1),
		.in_wire_0_2(horizontal_tile_1_19_to_tile_1_18_2),
		.in_wire_0_3(horizontal_tile_1_19_to_tile_1_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(51)
	);

	pe_tile pe_tile_1_19(
		.out_wire_3_0(vertical_tile_1_19_to_tile_0_19_0),
		.out_wire_3_1(vertical_tile_1_19_to_tile_0_19_1),
		.out_wire_3_2(vertical_tile_1_19_to_tile_0_19_2),
		.out_wire_3_3(vertical_tile_1_19_to_tile_0_19_3),
		.in_wire_3_0(vertical_tile_0_19_to_tile_1_19_0),
		.in_wire_3_1(vertical_tile_0_19_to_tile_1_19_1),
		.in_wire_3_2(vertical_tile_0_19_to_tile_1_19_2),
		.in_wire_3_3(vertical_tile_0_19_to_tile_1_19_3),
		.out_wire_1_0(vertical_tile_1_19_to_tile_2_19_0),
		.out_wire_1_1(vertical_tile_1_19_to_tile_2_19_1),
		.out_wire_1_2(vertical_tile_1_19_to_tile_2_19_2),
		.out_wire_1_3(vertical_tile_1_19_to_tile_2_19_3),
		.in_wire_1_0(vertical_tile_2_19_to_tile_1_19_0),
		.in_wire_1_1(vertical_tile_2_19_to_tile_1_19_1),
		.in_wire_1_2(vertical_tile_2_19_to_tile_1_19_2),
		.in_wire_1_3(vertical_tile_2_19_to_tile_1_19_3),
		.out_wire_2_0(horizontal_tile_1_19_to_tile_1_18_0),
		.out_wire_2_1(horizontal_tile_1_19_to_tile_1_18_1),
		.out_wire_2_2(horizontal_tile_1_19_to_tile_1_18_2),
		.out_wire_2_3(horizontal_tile_1_19_to_tile_1_18_3),
		.in_wire_2_0(horizontal_tile_1_18_to_tile_1_19_0),
		.in_wire_2_1(horizontal_tile_1_18_to_tile_1_19_1),
		.in_wire_2_2(horizontal_tile_1_18_to_tile_1_19_2),
		.in_wire_2_3(horizontal_tile_1_18_to_tile_1_19_3),
		.out_wire_0_0(horizontal_tile_1_19_to_tile_1_20_0),
		.out_wire_0_1(horizontal_tile_1_19_to_tile_1_20_1),
		.out_wire_0_2(horizontal_tile_1_19_to_tile_1_20_2),
		.out_wire_0_3(horizontal_tile_1_19_to_tile_1_20_3),
		.in_wire_0_0(horizontal_tile_1_20_to_tile_1_19_0),
		.in_wire_0_1(horizontal_tile_1_20_to_tile_1_19_1),
		.in_wire_0_2(horizontal_tile_1_20_to_tile_1_19_2),
		.in_wire_0_3(horizontal_tile_1_20_to_tile_1_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(52)
	);

	pe_tile pe_tile_1_20(
		.out_wire_3_0(vertical_tile_1_20_to_tile_0_20_0),
		.out_wire_3_1(vertical_tile_1_20_to_tile_0_20_1),
		.out_wire_3_2(vertical_tile_1_20_to_tile_0_20_2),
		.out_wire_3_3(vertical_tile_1_20_to_tile_0_20_3),
		.in_wire_3_0(vertical_tile_0_20_to_tile_1_20_0),
		.in_wire_3_1(vertical_tile_0_20_to_tile_1_20_1),
		.in_wire_3_2(vertical_tile_0_20_to_tile_1_20_2),
		.in_wire_3_3(vertical_tile_0_20_to_tile_1_20_3),
		.out_wire_1_0(vertical_tile_1_20_to_tile_2_20_0),
		.out_wire_1_1(vertical_tile_1_20_to_tile_2_20_1),
		.out_wire_1_2(vertical_tile_1_20_to_tile_2_20_2),
		.out_wire_1_3(vertical_tile_1_20_to_tile_2_20_3),
		.in_wire_1_0(vertical_tile_2_20_to_tile_1_20_0),
		.in_wire_1_1(vertical_tile_2_20_to_tile_1_20_1),
		.in_wire_1_2(vertical_tile_2_20_to_tile_1_20_2),
		.in_wire_1_3(vertical_tile_2_20_to_tile_1_20_3),
		.out_wire_2_0(horizontal_tile_1_20_to_tile_1_19_0),
		.out_wire_2_1(horizontal_tile_1_20_to_tile_1_19_1),
		.out_wire_2_2(horizontal_tile_1_20_to_tile_1_19_2),
		.out_wire_2_3(horizontal_tile_1_20_to_tile_1_19_3),
		.in_wire_2_0(horizontal_tile_1_19_to_tile_1_20_0),
		.in_wire_2_1(horizontal_tile_1_19_to_tile_1_20_1),
		.in_wire_2_2(horizontal_tile_1_19_to_tile_1_20_2),
		.in_wire_2_3(horizontal_tile_1_19_to_tile_1_20_3),
		.out_wire_0_0(horizontal_tile_1_20_to_tile_1_21_0),
		.out_wire_0_1(horizontal_tile_1_20_to_tile_1_21_1),
		.out_wire_0_2(horizontal_tile_1_20_to_tile_1_21_2),
		.out_wire_0_3(horizontal_tile_1_20_to_tile_1_21_3),
		.in_wire_0_0(horizontal_tile_1_21_to_tile_1_20_0),
		.in_wire_0_1(horizontal_tile_1_21_to_tile_1_20_1),
		.in_wire_0_2(horizontal_tile_1_21_to_tile_1_20_2),
		.in_wire_0_3(horizontal_tile_1_21_to_tile_1_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(53)
	);

	pe_tile pe_tile_1_21(
		.out_wire_3_0(vertical_tile_1_21_to_tile_0_21_0),
		.out_wire_3_1(vertical_tile_1_21_to_tile_0_21_1),
		.out_wire_3_2(vertical_tile_1_21_to_tile_0_21_2),
		.out_wire_3_3(vertical_tile_1_21_to_tile_0_21_3),
		.in_wire_3_0(vertical_tile_0_21_to_tile_1_21_0),
		.in_wire_3_1(vertical_tile_0_21_to_tile_1_21_1),
		.in_wire_3_2(vertical_tile_0_21_to_tile_1_21_2),
		.in_wire_3_3(vertical_tile_0_21_to_tile_1_21_3),
		.out_wire_1_0(vertical_tile_1_21_to_tile_2_21_0),
		.out_wire_1_1(vertical_tile_1_21_to_tile_2_21_1),
		.out_wire_1_2(vertical_tile_1_21_to_tile_2_21_2),
		.out_wire_1_3(vertical_tile_1_21_to_tile_2_21_3),
		.in_wire_1_0(vertical_tile_2_21_to_tile_1_21_0),
		.in_wire_1_1(vertical_tile_2_21_to_tile_1_21_1),
		.in_wire_1_2(vertical_tile_2_21_to_tile_1_21_2),
		.in_wire_1_3(vertical_tile_2_21_to_tile_1_21_3),
		.out_wire_2_0(horizontal_tile_1_21_to_tile_1_20_0),
		.out_wire_2_1(horizontal_tile_1_21_to_tile_1_20_1),
		.out_wire_2_2(horizontal_tile_1_21_to_tile_1_20_2),
		.out_wire_2_3(horizontal_tile_1_21_to_tile_1_20_3),
		.in_wire_2_0(horizontal_tile_1_20_to_tile_1_21_0),
		.in_wire_2_1(horizontal_tile_1_20_to_tile_1_21_1),
		.in_wire_2_2(horizontal_tile_1_20_to_tile_1_21_2),
		.in_wire_2_3(horizontal_tile_1_20_to_tile_1_21_3),
		.out_wire_0_0(horizontal_tile_1_21_to_tile_1_22_0),
		.out_wire_0_1(horizontal_tile_1_21_to_tile_1_22_1),
		.out_wire_0_2(horizontal_tile_1_21_to_tile_1_22_2),
		.out_wire_0_3(horizontal_tile_1_21_to_tile_1_22_3),
		.in_wire_0_0(horizontal_tile_1_22_to_tile_1_21_0),
		.in_wire_0_1(horizontal_tile_1_22_to_tile_1_21_1),
		.in_wire_0_2(horizontal_tile_1_22_to_tile_1_21_2),
		.in_wire_0_3(horizontal_tile_1_22_to_tile_1_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(54)
	);

	pe_tile pe_tile_1_22(
		.out_wire_3_0(vertical_tile_1_22_to_tile_0_22_0),
		.out_wire_3_1(vertical_tile_1_22_to_tile_0_22_1),
		.out_wire_3_2(vertical_tile_1_22_to_tile_0_22_2),
		.out_wire_3_3(vertical_tile_1_22_to_tile_0_22_3),
		.in_wire_3_0(vertical_tile_0_22_to_tile_1_22_0),
		.in_wire_3_1(vertical_tile_0_22_to_tile_1_22_1),
		.in_wire_3_2(vertical_tile_0_22_to_tile_1_22_2),
		.in_wire_3_3(vertical_tile_0_22_to_tile_1_22_3),
		.out_wire_1_0(vertical_tile_1_22_to_tile_2_22_0),
		.out_wire_1_1(vertical_tile_1_22_to_tile_2_22_1),
		.out_wire_1_2(vertical_tile_1_22_to_tile_2_22_2),
		.out_wire_1_3(vertical_tile_1_22_to_tile_2_22_3),
		.in_wire_1_0(vertical_tile_2_22_to_tile_1_22_0),
		.in_wire_1_1(vertical_tile_2_22_to_tile_1_22_1),
		.in_wire_1_2(vertical_tile_2_22_to_tile_1_22_2),
		.in_wire_1_3(vertical_tile_2_22_to_tile_1_22_3),
		.out_wire_2_0(horizontal_tile_1_22_to_tile_1_21_0),
		.out_wire_2_1(horizontal_tile_1_22_to_tile_1_21_1),
		.out_wire_2_2(horizontal_tile_1_22_to_tile_1_21_2),
		.out_wire_2_3(horizontal_tile_1_22_to_tile_1_21_3),
		.in_wire_2_0(horizontal_tile_1_21_to_tile_1_22_0),
		.in_wire_2_1(horizontal_tile_1_21_to_tile_1_22_1),
		.in_wire_2_2(horizontal_tile_1_21_to_tile_1_22_2),
		.in_wire_2_3(horizontal_tile_1_21_to_tile_1_22_3),
		.out_wire_0_0(horizontal_tile_1_22_to_tile_1_23_0),
		.out_wire_0_1(horizontal_tile_1_22_to_tile_1_23_1),
		.out_wire_0_2(horizontal_tile_1_22_to_tile_1_23_2),
		.out_wire_0_3(horizontal_tile_1_22_to_tile_1_23_3),
		.in_wire_0_0(horizontal_tile_1_23_to_tile_1_22_0),
		.in_wire_0_1(horizontal_tile_1_23_to_tile_1_22_1),
		.in_wire_0_2(horizontal_tile_1_23_to_tile_1_22_2),
		.in_wire_0_3(horizontal_tile_1_23_to_tile_1_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(55)
	);

	pe_tile pe_tile_1_23(
		.out_wire_3_0(vertical_tile_1_23_to_tile_0_23_0),
		.out_wire_3_1(vertical_tile_1_23_to_tile_0_23_1),
		.out_wire_3_2(vertical_tile_1_23_to_tile_0_23_2),
		.out_wire_3_3(vertical_tile_1_23_to_tile_0_23_3),
		.in_wire_3_0(vertical_tile_0_23_to_tile_1_23_0),
		.in_wire_3_1(vertical_tile_0_23_to_tile_1_23_1),
		.in_wire_3_2(vertical_tile_0_23_to_tile_1_23_2),
		.in_wire_3_3(vertical_tile_0_23_to_tile_1_23_3),
		.out_wire_1_0(vertical_tile_1_23_to_tile_2_23_0),
		.out_wire_1_1(vertical_tile_1_23_to_tile_2_23_1),
		.out_wire_1_2(vertical_tile_1_23_to_tile_2_23_2),
		.out_wire_1_3(vertical_tile_1_23_to_tile_2_23_3),
		.in_wire_1_0(vertical_tile_2_23_to_tile_1_23_0),
		.in_wire_1_1(vertical_tile_2_23_to_tile_1_23_1),
		.in_wire_1_2(vertical_tile_2_23_to_tile_1_23_2),
		.in_wire_1_3(vertical_tile_2_23_to_tile_1_23_3),
		.out_wire_2_0(horizontal_tile_1_23_to_tile_1_22_0),
		.out_wire_2_1(horizontal_tile_1_23_to_tile_1_22_1),
		.out_wire_2_2(horizontal_tile_1_23_to_tile_1_22_2),
		.out_wire_2_3(horizontal_tile_1_23_to_tile_1_22_3),
		.in_wire_2_0(horizontal_tile_1_22_to_tile_1_23_0),
		.in_wire_2_1(horizontal_tile_1_22_to_tile_1_23_1),
		.in_wire_2_2(horizontal_tile_1_22_to_tile_1_23_2),
		.in_wire_2_3(horizontal_tile_1_22_to_tile_1_23_3),
		.out_wire_0_0(horizontal_tile_1_23_to_tile_1_24_0),
		.out_wire_0_1(horizontal_tile_1_23_to_tile_1_24_1),
		.out_wire_0_2(horizontal_tile_1_23_to_tile_1_24_2),
		.out_wire_0_3(horizontal_tile_1_23_to_tile_1_24_3),
		.in_wire_0_0(horizontal_tile_1_24_to_tile_1_23_0),
		.in_wire_0_1(horizontal_tile_1_24_to_tile_1_23_1),
		.in_wire_0_2(horizontal_tile_1_24_to_tile_1_23_2),
		.in_wire_0_3(horizontal_tile_1_24_to_tile_1_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(56)
	);

	pe_tile pe_tile_1_24(
		.out_wire_3_0(vertical_tile_1_24_to_tile_0_24_0),
		.out_wire_3_1(vertical_tile_1_24_to_tile_0_24_1),
		.out_wire_3_2(vertical_tile_1_24_to_tile_0_24_2),
		.out_wire_3_3(vertical_tile_1_24_to_tile_0_24_3),
		.in_wire_3_0(vertical_tile_0_24_to_tile_1_24_0),
		.in_wire_3_1(vertical_tile_0_24_to_tile_1_24_1),
		.in_wire_3_2(vertical_tile_0_24_to_tile_1_24_2),
		.in_wire_3_3(vertical_tile_0_24_to_tile_1_24_3),
		.out_wire_1_0(vertical_tile_1_24_to_tile_2_24_0),
		.out_wire_1_1(vertical_tile_1_24_to_tile_2_24_1),
		.out_wire_1_2(vertical_tile_1_24_to_tile_2_24_2),
		.out_wire_1_3(vertical_tile_1_24_to_tile_2_24_3),
		.in_wire_1_0(vertical_tile_2_24_to_tile_1_24_0),
		.in_wire_1_1(vertical_tile_2_24_to_tile_1_24_1),
		.in_wire_1_2(vertical_tile_2_24_to_tile_1_24_2),
		.in_wire_1_3(vertical_tile_2_24_to_tile_1_24_3),
		.out_wire_2_0(horizontal_tile_1_24_to_tile_1_23_0),
		.out_wire_2_1(horizontal_tile_1_24_to_tile_1_23_1),
		.out_wire_2_2(horizontal_tile_1_24_to_tile_1_23_2),
		.out_wire_2_3(horizontal_tile_1_24_to_tile_1_23_3),
		.in_wire_2_0(horizontal_tile_1_23_to_tile_1_24_0),
		.in_wire_2_1(horizontal_tile_1_23_to_tile_1_24_1),
		.in_wire_2_2(horizontal_tile_1_23_to_tile_1_24_2),
		.in_wire_2_3(horizontal_tile_1_23_to_tile_1_24_3),
		.out_wire_0_0(horizontal_tile_1_24_to_tile_1_25_0),
		.out_wire_0_1(horizontal_tile_1_24_to_tile_1_25_1),
		.out_wire_0_2(horizontal_tile_1_24_to_tile_1_25_2),
		.out_wire_0_3(horizontal_tile_1_24_to_tile_1_25_3),
		.in_wire_0_0(horizontal_tile_1_25_to_tile_1_24_0),
		.in_wire_0_1(horizontal_tile_1_25_to_tile_1_24_1),
		.in_wire_0_2(horizontal_tile_1_25_to_tile_1_24_2),
		.in_wire_0_3(horizontal_tile_1_25_to_tile_1_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(57)
	);

	pe_tile pe_tile_1_25(
		.out_wire_3_0(vertical_tile_1_25_to_tile_0_25_0),
		.out_wire_3_1(vertical_tile_1_25_to_tile_0_25_1),
		.out_wire_3_2(vertical_tile_1_25_to_tile_0_25_2),
		.out_wire_3_3(vertical_tile_1_25_to_tile_0_25_3),
		.in_wire_3_0(vertical_tile_0_25_to_tile_1_25_0),
		.in_wire_3_1(vertical_tile_0_25_to_tile_1_25_1),
		.in_wire_3_2(vertical_tile_0_25_to_tile_1_25_2),
		.in_wire_3_3(vertical_tile_0_25_to_tile_1_25_3),
		.out_wire_1_0(vertical_tile_1_25_to_tile_2_25_0),
		.out_wire_1_1(vertical_tile_1_25_to_tile_2_25_1),
		.out_wire_1_2(vertical_tile_1_25_to_tile_2_25_2),
		.out_wire_1_3(vertical_tile_1_25_to_tile_2_25_3),
		.in_wire_1_0(vertical_tile_2_25_to_tile_1_25_0),
		.in_wire_1_1(vertical_tile_2_25_to_tile_1_25_1),
		.in_wire_1_2(vertical_tile_2_25_to_tile_1_25_2),
		.in_wire_1_3(vertical_tile_2_25_to_tile_1_25_3),
		.out_wire_2_0(horizontal_tile_1_25_to_tile_1_24_0),
		.out_wire_2_1(horizontal_tile_1_25_to_tile_1_24_1),
		.out_wire_2_2(horizontal_tile_1_25_to_tile_1_24_2),
		.out_wire_2_3(horizontal_tile_1_25_to_tile_1_24_3),
		.in_wire_2_0(horizontal_tile_1_24_to_tile_1_25_0),
		.in_wire_2_1(horizontal_tile_1_24_to_tile_1_25_1),
		.in_wire_2_2(horizontal_tile_1_24_to_tile_1_25_2),
		.in_wire_2_3(horizontal_tile_1_24_to_tile_1_25_3),
		.out_wire_0_0(horizontal_tile_1_25_to_tile_1_26_0),
		.out_wire_0_1(horizontal_tile_1_25_to_tile_1_26_1),
		.out_wire_0_2(horizontal_tile_1_25_to_tile_1_26_2),
		.out_wire_0_3(horizontal_tile_1_25_to_tile_1_26_3),
		.in_wire_0_0(horizontal_tile_1_26_to_tile_1_25_0),
		.in_wire_0_1(horizontal_tile_1_26_to_tile_1_25_1),
		.in_wire_0_2(horizontal_tile_1_26_to_tile_1_25_2),
		.in_wire_0_3(horizontal_tile_1_26_to_tile_1_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(58)
	);

	pe_tile pe_tile_1_26(
		.out_wire_3_0(vertical_tile_1_26_to_tile_0_26_0),
		.out_wire_3_1(vertical_tile_1_26_to_tile_0_26_1),
		.out_wire_3_2(vertical_tile_1_26_to_tile_0_26_2),
		.out_wire_3_3(vertical_tile_1_26_to_tile_0_26_3),
		.in_wire_3_0(vertical_tile_0_26_to_tile_1_26_0),
		.in_wire_3_1(vertical_tile_0_26_to_tile_1_26_1),
		.in_wire_3_2(vertical_tile_0_26_to_tile_1_26_2),
		.in_wire_3_3(vertical_tile_0_26_to_tile_1_26_3),
		.out_wire_1_0(vertical_tile_1_26_to_tile_2_26_0),
		.out_wire_1_1(vertical_tile_1_26_to_tile_2_26_1),
		.out_wire_1_2(vertical_tile_1_26_to_tile_2_26_2),
		.out_wire_1_3(vertical_tile_1_26_to_tile_2_26_3),
		.in_wire_1_0(vertical_tile_2_26_to_tile_1_26_0),
		.in_wire_1_1(vertical_tile_2_26_to_tile_1_26_1),
		.in_wire_1_2(vertical_tile_2_26_to_tile_1_26_2),
		.in_wire_1_3(vertical_tile_2_26_to_tile_1_26_3),
		.out_wire_2_0(horizontal_tile_1_26_to_tile_1_25_0),
		.out_wire_2_1(horizontal_tile_1_26_to_tile_1_25_1),
		.out_wire_2_2(horizontal_tile_1_26_to_tile_1_25_2),
		.out_wire_2_3(horizontal_tile_1_26_to_tile_1_25_3),
		.in_wire_2_0(horizontal_tile_1_25_to_tile_1_26_0),
		.in_wire_2_1(horizontal_tile_1_25_to_tile_1_26_1),
		.in_wire_2_2(horizontal_tile_1_25_to_tile_1_26_2),
		.in_wire_2_3(horizontal_tile_1_25_to_tile_1_26_3),
		.out_wire_0_0(horizontal_tile_1_26_to_tile_1_27_0),
		.out_wire_0_1(horizontal_tile_1_26_to_tile_1_27_1),
		.out_wire_0_2(horizontal_tile_1_26_to_tile_1_27_2),
		.out_wire_0_3(horizontal_tile_1_26_to_tile_1_27_3),
		.in_wire_0_0(horizontal_tile_1_27_to_tile_1_26_0),
		.in_wire_0_1(horizontal_tile_1_27_to_tile_1_26_1),
		.in_wire_0_2(horizontal_tile_1_27_to_tile_1_26_2),
		.in_wire_0_3(horizontal_tile_1_27_to_tile_1_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(59)
	);

	pe_tile pe_tile_1_27(
		.out_wire_3_0(vertical_tile_1_27_to_tile_0_27_0),
		.out_wire_3_1(vertical_tile_1_27_to_tile_0_27_1),
		.out_wire_3_2(vertical_tile_1_27_to_tile_0_27_2),
		.out_wire_3_3(vertical_tile_1_27_to_tile_0_27_3),
		.in_wire_3_0(vertical_tile_0_27_to_tile_1_27_0),
		.in_wire_3_1(vertical_tile_0_27_to_tile_1_27_1),
		.in_wire_3_2(vertical_tile_0_27_to_tile_1_27_2),
		.in_wire_3_3(vertical_tile_0_27_to_tile_1_27_3),
		.out_wire_1_0(vertical_tile_1_27_to_tile_2_27_0),
		.out_wire_1_1(vertical_tile_1_27_to_tile_2_27_1),
		.out_wire_1_2(vertical_tile_1_27_to_tile_2_27_2),
		.out_wire_1_3(vertical_tile_1_27_to_tile_2_27_3),
		.in_wire_1_0(vertical_tile_2_27_to_tile_1_27_0),
		.in_wire_1_1(vertical_tile_2_27_to_tile_1_27_1),
		.in_wire_1_2(vertical_tile_2_27_to_tile_1_27_2),
		.in_wire_1_3(vertical_tile_2_27_to_tile_1_27_3),
		.out_wire_2_0(horizontal_tile_1_27_to_tile_1_26_0),
		.out_wire_2_1(horizontal_tile_1_27_to_tile_1_26_1),
		.out_wire_2_2(horizontal_tile_1_27_to_tile_1_26_2),
		.out_wire_2_3(horizontal_tile_1_27_to_tile_1_26_3),
		.in_wire_2_0(horizontal_tile_1_26_to_tile_1_27_0),
		.in_wire_2_1(horizontal_tile_1_26_to_tile_1_27_1),
		.in_wire_2_2(horizontal_tile_1_26_to_tile_1_27_2),
		.in_wire_2_3(horizontal_tile_1_26_to_tile_1_27_3),
		.out_wire_0_0(horizontal_tile_1_27_to_tile_1_28_0),
		.out_wire_0_1(horizontal_tile_1_27_to_tile_1_28_1),
		.out_wire_0_2(horizontal_tile_1_27_to_tile_1_28_2),
		.out_wire_0_3(horizontal_tile_1_27_to_tile_1_28_3),
		.in_wire_0_0(horizontal_tile_1_28_to_tile_1_27_0),
		.in_wire_0_1(horizontal_tile_1_28_to_tile_1_27_1),
		.in_wire_0_2(horizontal_tile_1_28_to_tile_1_27_2),
		.in_wire_0_3(horizontal_tile_1_28_to_tile_1_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(60)
	);

	pe_tile pe_tile_1_28(
		.out_wire_3_0(vertical_tile_1_28_to_tile_0_28_0),
		.out_wire_3_1(vertical_tile_1_28_to_tile_0_28_1),
		.out_wire_3_2(vertical_tile_1_28_to_tile_0_28_2),
		.out_wire_3_3(vertical_tile_1_28_to_tile_0_28_3),
		.in_wire_3_0(vertical_tile_0_28_to_tile_1_28_0),
		.in_wire_3_1(vertical_tile_0_28_to_tile_1_28_1),
		.in_wire_3_2(vertical_tile_0_28_to_tile_1_28_2),
		.in_wire_3_3(vertical_tile_0_28_to_tile_1_28_3),
		.out_wire_1_0(vertical_tile_1_28_to_tile_2_28_0),
		.out_wire_1_1(vertical_tile_1_28_to_tile_2_28_1),
		.out_wire_1_2(vertical_tile_1_28_to_tile_2_28_2),
		.out_wire_1_3(vertical_tile_1_28_to_tile_2_28_3),
		.in_wire_1_0(vertical_tile_2_28_to_tile_1_28_0),
		.in_wire_1_1(vertical_tile_2_28_to_tile_1_28_1),
		.in_wire_1_2(vertical_tile_2_28_to_tile_1_28_2),
		.in_wire_1_3(vertical_tile_2_28_to_tile_1_28_3),
		.out_wire_2_0(horizontal_tile_1_28_to_tile_1_27_0),
		.out_wire_2_1(horizontal_tile_1_28_to_tile_1_27_1),
		.out_wire_2_2(horizontal_tile_1_28_to_tile_1_27_2),
		.out_wire_2_3(horizontal_tile_1_28_to_tile_1_27_3),
		.in_wire_2_0(horizontal_tile_1_27_to_tile_1_28_0),
		.in_wire_2_1(horizontal_tile_1_27_to_tile_1_28_1),
		.in_wire_2_2(horizontal_tile_1_27_to_tile_1_28_2),
		.in_wire_2_3(horizontal_tile_1_27_to_tile_1_28_3),
		.out_wire_0_0(horizontal_tile_1_28_to_tile_1_29_0),
		.out_wire_0_1(horizontal_tile_1_28_to_tile_1_29_1),
		.out_wire_0_2(horizontal_tile_1_28_to_tile_1_29_2),
		.out_wire_0_3(horizontal_tile_1_28_to_tile_1_29_3),
		.in_wire_0_0(horizontal_tile_1_29_to_tile_1_28_0),
		.in_wire_0_1(horizontal_tile_1_29_to_tile_1_28_1),
		.in_wire_0_2(horizontal_tile_1_29_to_tile_1_28_2),
		.in_wire_0_3(horizontal_tile_1_29_to_tile_1_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(61)
	);

	pe_tile pe_tile_1_29(
		.out_wire_3_0(vertical_tile_1_29_to_tile_0_29_0),
		.out_wire_3_1(vertical_tile_1_29_to_tile_0_29_1),
		.out_wire_3_2(vertical_tile_1_29_to_tile_0_29_2),
		.out_wire_3_3(vertical_tile_1_29_to_tile_0_29_3),
		.in_wire_3_0(vertical_tile_0_29_to_tile_1_29_0),
		.in_wire_3_1(vertical_tile_0_29_to_tile_1_29_1),
		.in_wire_3_2(vertical_tile_0_29_to_tile_1_29_2),
		.in_wire_3_3(vertical_tile_0_29_to_tile_1_29_3),
		.out_wire_1_0(vertical_tile_1_29_to_tile_2_29_0),
		.out_wire_1_1(vertical_tile_1_29_to_tile_2_29_1),
		.out_wire_1_2(vertical_tile_1_29_to_tile_2_29_2),
		.out_wire_1_3(vertical_tile_1_29_to_tile_2_29_3),
		.in_wire_1_0(vertical_tile_2_29_to_tile_1_29_0),
		.in_wire_1_1(vertical_tile_2_29_to_tile_1_29_1),
		.in_wire_1_2(vertical_tile_2_29_to_tile_1_29_2),
		.in_wire_1_3(vertical_tile_2_29_to_tile_1_29_3),
		.out_wire_2_0(horizontal_tile_1_29_to_tile_1_28_0),
		.out_wire_2_1(horizontal_tile_1_29_to_tile_1_28_1),
		.out_wire_2_2(horizontal_tile_1_29_to_tile_1_28_2),
		.out_wire_2_3(horizontal_tile_1_29_to_tile_1_28_3),
		.in_wire_2_0(horizontal_tile_1_28_to_tile_1_29_0),
		.in_wire_2_1(horizontal_tile_1_28_to_tile_1_29_1),
		.in_wire_2_2(horizontal_tile_1_28_to_tile_1_29_2),
		.in_wire_2_3(horizontal_tile_1_28_to_tile_1_29_3),
		.out_wire_0_0(horizontal_tile_1_29_to_tile_1_30_0),
		.out_wire_0_1(horizontal_tile_1_29_to_tile_1_30_1),
		.out_wire_0_2(horizontal_tile_1_29_to_tile_1_30_2),
		.out_wire_0_3(horizontal_tile_1_29_to_tile_1_30_3),
		.in_wire_0_0(horizontal_tile_1_30_to_tile_1_29_0),
		.in_wire_0_1(horizontal_tile_1_30_to_tile_1_29_1),
		.in_wire_0_2(horizontal_tile_1_30_to_tile_1_29_2),
		.in_wire_0_3(horizontal_tile_1_30_to_tile_1_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(62)
	);

	pe_tile pe_tile_1_30(
		.out_wire_3_0(vertical_tile_1_30_to_tile_0_30_0),
		.out_wire_3_1(vertical_tile_1_30_to_tile_0_30_1),
		.out_wire_3_2(vertical_tile_1_30_to_tile_0_30_2),
		.out_wire_3_3(vertical_tile_1_30_to_tile_0_30_3),
		.in_wire_3_0(vertical_tile_0_30_to_tile_1_30_0),
		.in_wire_3_1(vertical_tile_0_30_to_tile_1_30_1),
		.in_wire_3_2(vertical_tile_0_30_to_tile_1_30_2),
		.in_wire_3_3(vertical_tile_0_30_to_tile_1_30_3),
		.out_wire_1_0(vertical_tile_1_30_to_tile_2_30_0),
		.out_wire_1_1(vertical_tile_1_30_to_tile_2_30_1),
		.out_wire_1_2(vertical_tile_1_30_to_tile_2_30_2),
		.out_wire_1_3(vertical_tile_1_30_to_tile_2_30_3),
		.in_wire_1_0(vertical_tile_2_30_to_tile_1_30_0),
		.in_wire_1_1(vertical_tile_2_30_to_tile_1_30_1),
		.in_wire_1_2(vertical_tile_2_30_to_tile_1_30_2),
		.in_wire_1_3(vertical_tile_2_30_to_tile_1_30_3),
		.out_wire_2_0(horizontal_tile_1_30_to_tile_1_29_0),
		.out_wire_2_1(horizontal_tile_1_30_to_tile_1_29_1),
		.out_wire_2_2(horizontal_tile_1_30_to_tile_1_29_2),
		.out_wire_2_3(horizontal_tile_1_30_to_tile_1_29_3),
		.in_wire_2_0(horizontal_tile_1_29_to_tile_1_30_0),
		.in_wire_2_1(horizontal_tile_1_29_to_tile_1_30_1),
		.in_wire_2_2(horizontal_tile_1_29_to_tile_1_30_2),
		.in_wire_2_3(horizontal_tile_1_29_to_tile_1_30_3),
		.out_wire_0_0(horizontal_tile_1_30_to_tile_1_31_0),
		.out_wire_0_1(horizontal_tile_1_30_to_tile_1_31_1),
		.out_wire_0_2(horizontal_tile_1_30_to_tile_1_31_2),
		.out_wire_0_3(horizontal_tile_1_30_to_tile_1_31_3),
		.in_wire_0_0(horizontal_tile_1_31_to_tile_1_30_0),
		.in_wire_0_1(horizontal_tile_1_31_to_tile_1_30_1),
		.in_wire_0_2(horizontal_tile_1_31_to_tile_1_30_2),
		.in_wire_0_3(horizontal_tile_1_31_to_tile_1_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(63)
	);

	pe_tile_right pe_tile_1_31(
		.out_wire_3_0(vertical_tile_1_31_to_tile_0_31_0),
		.out_wire_3_1(vertical_tile_1_31_to_tile_0_31_1),
		.out_wire_3_2(vertical_tile_1_31_to_tile_0_31_2),
		.out_wire_3_3(vertical_tile_1_31_to_tile_0_31_3),
		.in_wire_3_0(vertical_tile_0_31_to_tile_1_31_0),
		.in_wire_3_1(vertical_tile_0_31_to_tile_1_31_1),
		.in_wire_3_2(vertical_tile_0_31_to_tile_1_31_2),
		.in_wire_3_3(vertical_tile_0_31_to_tile_1_31_3),
		.out_wire_1_0(vertical_tile_1_31_to_tile_2_31_0),
		.out_wire_1_1(vertical_tile_1_31_to_tile_2_31_1),
		.out_wire_1_2(vertical_tile_1_31_to_tile_2_31_2),
		.out_wire_1_3(vertical_tile_1_31_to_tile_2_31_3),
		.in_wire_1_0(vertical_tile_2_31_to_tile_1_31_0),
		.in_wire_1_1(vertical_tile_2_31_to_tile_1_31_1),
		.in_wire_1_2(vertical_tile_2_31_to_tile_1_31_2),
		.in_wire_1_3(vertical_tile_2_31_to_tile_1_31_3),
		.out_wire_2_0(horizontal_tile_1_31_to_tile_1_30_0),
		.out_wire_2_1(horizontal_tile_1_31_to_tile_1_30_1),
		.out_wire_2_2(horizontal_tile_1_31_to_tile_1_30_2),
		.out_wire_2_3(horizontal_tile_1_31_to_tile_1_30_3),
		.in_wire_2_0(horizontal_tile_1_30_to_tile_1_31_0),
		.in_wire_2_1(horizontal_tile_1_30_to_tile_1_31_1),
		.in_wire_2_2(horizontal_tile_1_30_to_tile_1_31_2),
		.in_wire_2_3(horizontal_tile_1_30_to_tile_1_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(64)
	);

	pe_tile_left pe_tile_2_0(
		.out_wire_3_0(vertical_tile_2_0_to_tile_1_0_0),
		.out_wire_3_1(vertical_tile_2_0_to_tile_1_0_1),
		.out_wire_3_2(vertical_tile_2_0_to_tile_1_0_2),
		.out_wire_3_3(vertical_tile_2_0_to_tile_1_0_3),
		.in_wire_3_0(vertical_tile_1_0_to_tile_2_0_0),
		.in_wire_3_1(vertical_tile_1_0_to_tile_2_0_1),
		.in_wire_3_2(vertical_tile_1_0_to_tile_2_0_2),
		.in_wire_3_3(vertical_tile_1_0_to_tile_2_0_3),
		.out_wire_1_0(vertical_tile_2_0_to_tile_3_0_0),
		.out_wire_1_1(vertical_tile_2_0_to_tile_3_0_1),
		.out_wire_1_2(vertical_tile_2_0_to_tile_3_0_2),
		.out_wire_1_3(vertical_tile_2_0_to_tile_3_0_3),
		.in_wire_1_0(vertical_tile_3_0_to_tile_2_0_0),
		.in_wire_1_1(vertical_tile_3_0_to_tile_2_0_1),
		.in_wire_1_2(vertical_tile_3_0_to_tile_2_0_2),
		.in_wire_1_3(vertical_tile_3_0_to_tile_2_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_2_0_to_tile_2_1_0),
		.out_wire_0_1(horizontal_tile_2_0_to_tile_2_1_1),
		.out_wire_0_2(horizontal_tile_2_0_to_tile_2_1_2),
		.out_wire_0_3(horizontal_tile_2_0_to_tile_2_1_3),
		.in_wire_0_0(horizontal_tile_2_1_to_tile_2_0_0),
		.in_wire_0_1(horizontal_tile_2_1_to_tile_2_0_1),
		.in_wire_0_2(horizontal_tile_2_1_to_tile_2_0_2),
		.in_wire_0_3(horizontal_tile_2_1_to_tile_2_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(65)
	);

	pe_tile pe_tile_2_1(
		.out_wire_3_0(vertical_tile_2_1_to_tile_1_1_0),
		.out_wire_3_1(vertical_tile_2_1_to_tile_1_1_1),
		.out_wire_3_2(vertical_tile_2_1_to_tile_1_1_2),
		.out_wire_3_3(vertical_tile_2_1_to_tile_1_1_3),
		.in_wire_3_0(vertical_tile_1_1_to_tile_2_1_0),
		.in_wire_3_1(vertical_tile_1_1_to_tile_2_1_1),
		.in_wire_3_2(vertical_tile_1_1_to_tile_2_1_2),
		.in_wire_3_3(vertical_tile_1_1_to_tile_2_1_3),
		.out_wire_1_0(vertical_tile_2_1_to_tile_3_1_0),
		.out_wire_1_1(vertical_tile_2_1_to_tile_3_1_1),
		.out_wire_1_2(vertical_tile_2_1_to_tile_3_1_2),
		.out_wire_1_3(vertical_tile_2_1_to_tile_3_1_3),
		.in_wire_1_0(vertical_tile_3_1_to_tile_2_1_0),
		.in_wire_1_1(vertical_tile_3_1_to_tile_2_1_1),
		.in_wire_1_2(vertical_tile_3_1_to_tile_2_1_2),
		.in_wire_1_3(vertical_tile_3_1_to_tile_2_1_3),
		.out_wire_2_0(horizontal_tile_2_1_to_tile_2_0_0),
		.out_wire_2_1(horizontal_tile_2_1_to_tile_2_0_1),
		.out_wire_2_2(horizontal_tile_2_1_to_tile_2_0_2),
		.out_wire_2_3(horizontal_tile_2_1_to_tile_2_0_3),
		.in_wire_2_0(horizontal_tile_2_0_to_tile_2_1_0),
		.in_wire_2_1(horizontal_tile_2_0_to_tile_2_1_1),
		.in_wire_2_2(horizontal_tile_2_0_to_tile_2_1_2),
		.in_wire_2_3(horizontal_tile_2_0_to_tile_2_1_3),
		.out_wire_0_0(horizontal_tile_2_1_to_tile_2_2_0),
		.out_wire_0_1(horizontal_tile_2_1_to_tile_2_2_1),
		.out_wire_0_2(horizontal_tile_2_1_to_tile_2_2_2),
		.out_wire_0_3(horizontal_tile_2_1_to_tile_2_2_3),
		.in_wire_0_0(horizontal_tile_2_2_to_tile_2_1_0),
		.in_wire_0_1(horizontal_tile_2_2_to_tile_2_1_1),
		.in_wire_0_2(horizontal_tile_2_2_to_tile_2_1_2),
		.in_wire_0_3(horizontal_tile_2_2_to_tile_2_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(66)
	);

	pe_tile pe_tile_2_2(
		.out_wire_3_0(vertical_tile_2_2_to_tile_1_2_0),
		.out_wire_3_1(vertical_tile_2_2_to_tile_1_2_1),
		.out_wire_3_2(vertical_tile_2_2_to_tile_1_2_2),
		.out_wire_3_3(vertical_tile_2_2_to_tile_1_2_3),
		.in_wire_3_0(vertical_tile_1_2_to_tile_2_2_0),
		.in_wire_3_1(vertical_tile_1_2_to_tile_2_2_1),
		.in_wire_3_2(vertical_tile_1_2_to_tile_2_2_2),
		.in_wire_3_3(vertical_tile_1_2_to_tile_2_2_3),
		.out_wire_1_0(vertical_tile_2_2_to_tile_3_2_0),
		.out_wire_1_1(vertical_tile_2_2_to_tile_3_2_1),
		.out_wire_1_2(vertical_tile_2_2_to_tile_3_2_2),
		.out_wire_1_3(vertical_tile_2_2_to_tile_3_2_3),
		.in_wire_1_0(vertical_tile_3_2_to_tile_2_2_0),
		.in_wire_1_1(vertical_tile_3_2_to_tile_2_2_1),
		.in_wire_1_2(vertical_tile_3_2_to_tile_2_2_2),
		.in_wire_1_3(vertical_tile_3_2_to_tile_2_2_3),
		.out_wire_2_0(horizontal_tile_2_2_to_tile_2_1_0),
		.out_wire_2_1(horizontal_tile_2_2_to_tile_2_1_1),
		.out_wire_2_2(horizontal_tile_2_2_to_tile_2_1_2),
		.out_wire_2_3(horizontal_tile_2_2_to_tile_2_1_3),
		.in_wire_2_0(horizontal_tile_2_1_to_tile_2_2_0),
		.in_wire_2_1(horizontal_tile_2_1_to_tile_2_2_1),
		.in_wire_2_2(horizontal_tile_2_1_to_tile_2_2_2),
		.in_wire_2_3(horizontal_tile_2_1_to_tile_2_2_3),
		.out_wire_0_0(horizontal_tile_2_2_to_tile_2_3_0),
		.out_wire_0_1(horizontal_tile_2_2_to_tile_2_3_1),
		.out_wire_0_2(horizontal_tile_2_2_to_tile_2_3_2),
		.out_wire_0_3(horizontal_tile_2_2_to_tile_2_3_3),
		.in_wire_0_0(horizontal_tile_2_3_to_tile_2_2_0),
		.in_wire_0_1(horizontal_tile_2_3_to_tile_2_2_1),
		.in_wire_0_2(horizontal_tile_2_3_to_tile_2_2_2),
		.in_wire_0_3(horizontal_tile_2_3_to_tile_2_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(67)
	);

	pe_tile pe_tile_2_3(
		.out_wire_3_0(vertical_tile_2_3_to_tile_1_3_0),
		.out_wire_3_1(vertical_tile_2_3_to_tile_1_3_1),
		.out_wire_3_2(vertical_tile_2_3_to_tile_1_3_2),
		.out_wire_3_3(vertical_tile_2_3_to_tile_1_3_3),
		.in_wire_3_0(vertical_tile_1_3_to_tile_2_3_0),
		.in_wire_3_1(vertical_tile_1_3_to_tile_2_3_1),
		.in_wire_3_2(vertical_tile_1_3_to_tile_2_3_2),
		.in_wire_3_3(vertical_tile_1_3_to_tile_2_3_3),
		.out_wire_1_0(vertical_tile_2_3_to_tile_3_3_0),
		.out_wire_1_1(vertical_tile_2_3_to_tile_3_3_1),
		.out_wire_1_2(vertical_tile_2_3_to_tile_3_3_2),
		.out_wire_1_3(vertical_tile_2_3_to_tile_3_3_3),
		.in_wire_1_0(vertical_tile_3_3_to_tile_2_3_0),
		.in_wire_1_1(vertical_tile_3_3_to_tile_2_3_1),
		.in_wire_1_2(vertical_tile_3_3_to_tile_2_3_2),
		.in_wire_1_3(vertical_tile_3_3_to_tile_2_3_3),
		.out_wire_2_0(horizontal_tile_2_3_to_tile_2_2_0),
		.out_wire_2_1(horizontal_tile_2_3_to_tile_2_2_1),
		.out_wire_2_2(horizontal_tile_2_3_to_tile_2_2_2),
		.out_wire_2_3(horizontal_tile_2_3_to_tile_2_2_3),
		.in_wire_2_0(horizontal_tile_2_2_to_tile_2_3_0),
		.in_wire_2_1(horizontal_tile_2_2_to_tile_2_3_1),
		.in_wire_2_2(horizontal_tile_2_2_to_tile_2_3_2),
		.in_wire_2_3(horizontal_tile_2_2_to_tile_2_3_3),
		.out_wire_0_0(horizontal_tile_2_3_to_tile_2_4_0),
		.out_wire_0_1(horizontal_tile_2_3_to_tile_2_4_1),
		.out_wire_0_2(horizontal_tile_2_3_to_tile_2_4_2),
		.out_wire_0_3(horizontal_tile_2_3_to_tile_2_4_3),
		.in_wire_0_0(horizontal_tile_2_4_to_tile_2_3_0),
		.in_wire_0_1(horizontal_tile_2_4_to_tile_2_3_1),
		.in_wire_0_2(horizontal_tile_2_4_to_tile_2_3_2),
		.in_wire_0_3(horizontal_tile_2_4_to_tile_2_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(68)
	);

	pe_tile pe_tile_2_4(
		.out_wire_3_0(vertical_tile_2_4_to_tile_1_4_0),
		.out_wire_3_1(vertical_tile_2_4_to_tile_1_4_1),
		.out_wire_3_2(vertical_tile_2_4_to_tile_1_4_2),
		.out_wire_3_3(vertical_tile_2_4_to_tile_1_4_3),
		.in_wire_3_0(vertical_tile_1_4_to_tile_2_4_0),
		.in_wire_3_1(vertical_tile_1_4_to_tile_2_4_1),
		.in_wire_3_2(vertical_tile_1_4_to_tile_2_4_2),
		.in_wire_3_3(vertical_tile_1_4_to_tile_2_4_3),
		.out_wire_1_0(vertical_tile_2_4_to_tile_3_4_0),
		.out_wire_1_1(vertical_tile_2_4_to_tile_3_4_1),
		.out_wire_1_2(vertical_tile_2_4_to_tile_3_4_2),
		.out_wire_1_3(vertical_tile_2_4_to_tile_3_4_3),
		.in_wire_1_0(vertical_tile_3_4_to_tile_2_4_0),
		.in_wire_1_1(vertical_tile_3_4_to_tile_2_4_1),
		.in_wire_1_2(vertical_tile_3_4_to_tile_2_4_2),
		.in_wire_1_3(vertical_tile_3_4_to_tile_2_4_3),
		.out_wire_2_0(horizontal_tile_2_4_to_tile_2_3_0),
		.out_wire_2_1(horizontal_tile_2_4_to_tile_2_3_1),
		.out_wire_2_2(horizontal_tile_2_4_to_tile_2_3_2),
		.out_wire_2_3(horizontal_tile_2_4_to_tile_2_3_3),
		.in_wire_2_0(horizontal_tile_2_3_to_tile_2_4_0),
		.in_wire_2_1(horizontal_tile_2_3_to_tile_2_4_1),
		.in_wire_2_2(horizontal_tile_2_3_to_tile_2_4_2),
		.in_wire_2_3(horizontal_tile_2_3_to_tile_2_4_3),
		.out_wire_0_0(horizontal_tile_2_4_to_tile_2_5_0),
		.out_wire_0_1(horizontal_tile_2_4_to_tile_2_5_1),
		.out_wire_0_2(horizontal_tile_2_4_to_tile_2_5_2),
		.out_wire_0_3(horizontal_tile_2_4_to_tile_2_5_3),
		.in_wire_0_0(horizontal_tile_2_5_to_tile_2_4_0),
		.in_wire_0_1(horizontal_tile_2_5_to_tile_2_4_1),
		.in_wire_0_2(horizontal_tile_2_5_to_tile_2_4_2),
		.in_wire_0_3(horizontal_tile_2_5_to_tile_2_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(69)
	);

	pe_tile pe_tile_2_5(
		.out_wire_3_0(vertical_tile_2_5_to_tile_1_5_0),
		.out_wire_3_1(vertical_tile_2_5_to_tile_1_5_1),
		.out_wire_3_2(vertical_tile_2_5_to_tile_1_5_2),
		.out_wire_3_3(vertical_tile_2_5_to_tile_1_5_3),
		.in_wire_3_0(vertical_tile_1_5_to_tile_2_5_0),
		.in_wire_3_1(vertical_tile_1_5_to_tile_2_5_1),
		.in_wire_3_2(vertical_tile_1_5_to_tile_2_5_2),
		.in_wire_3_3(vertical_tile_1_5_to_tile_2_5_3),
		.out_wire_1_0(vertical_tile_2_5_to_tile_3_5_0),
		.out_wire_1_1(vertical_tile_2_5_to_tile_3_5_1),
		.out_wire_1_2(vertical_tile_2_5_to_tile_3_5_2),
		.out_wire_1_3(vertical_tile_2_5_to_tile_3_5_3),
		.in_wire_1_0(vertical_tile_3_5_to_tile_2_5_0),
		.in_wire_1_1(vertical_tile_3_5_to_tile_2_5_1),
		.in_wire_1_2(vertical_tile_3_5_to_tile_2_5_2),
		.in_wire_1_3(vertical_tile_3_5_to_tile_2_5_3),
		.out_wire_2_0(horizontal_tile_2_5_to_tile_2_4_0),
		.out_wire_2_1(horizontal_tile_2_5_to_tile_2_4_1),
		.out_wire_2_2(horizontal_tile_2_5_to_tile_2_4_2),
		.out_wire_2_3(horizontal_tile_2_5_to_tile_2_4_3),
		.in_wire_2_0(horizontal_tile_2_4_to_tile_2_5_0),
		.in_wire_2_1(horizontal_tile_2_4_to_tile_2_5_1),
		.in_wire_2_2(horizontal_tile_2_4_to_tile_2_5_2),
		.in_wire_2_3(horizontal_tile_2_4_to_tile_2_5_3),
		.out_wire_0_0(horizontal_tile_2_5_to_tile_2_6_0),
		.out_wire_0_1(horizontal_tile_2_5_to_tile_2_6_1),
		.out_wire_0_2(horizontal_tile_2_5_to_tile_2_6_2),
		.out_wire_0_3(horizontal_tile_2_5_to_tile_2_6_3),
		.in_wire_0_0(horizontal_tile_2_6_to_tile_2_5_0),
		.in_wire_0_1(horizontal_tile_2_6_to_tile_2_5_1),
		.in_wire_0_2(horizontal_tile_2_6_to_tile_2_5_2),
		.in_wire_0_3(horizontal_tile_2_6_to_tile_2_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(70)
	);

	pe_tile pe_tile_2_6(
		.out_wire_3_0(vertical_tile_2_6_to_tile_1_6_0),
		.out_wire_3_1(vertical_tile_2_6_to_tile_1_6_1),
		.out_wire_3_2(vertical_tile_2_6_to_tile_1_6_2),
		.out_wire_3_3(vertical_tile_2_6_to_tile_1_6_3),
		.in_wire_3_0(vertical_tile_1_6_to_tile_2_6_0),
		.in_wire_3_1(vertical_tile_1_6_to_tile_2_6_1),
		.in_wire_3_2(vertical_tile_1_6_to_tile_2_6_2),
		.in_wire_3_3(vertical_tile_1_6_to_tile_2_6_3),
		.out_wire_1_0(vertical_tile_2_6_to_tile_3_6_0),
		.out_wire_1_1(vertical_tile_2_6_to_tile_3_6_1),
		.out_wire_1_2(vertical_tile_2_6_to_tile_3_6_2),
		.out_wire_1_3(vertical_tile_2_6_to_tile_3_6_3),
		.in_wire_1_0(vertical_tile_3_6_to_tile_2_6_0),
		.in_wire_1_1(vertical_tile_3_6_to_tile_2_6_1),
		.in_wire_1_2(vertical_tile_3_6_to_tile_2_6_2),
		.in_wire_1_3(vertical_tile_3_6_to_tile_2_6_3),
		.out_wire_2_0(horizontal_tile_2_6_to_tile_2_5_0),
		.out_wire_2_1(horizontal_tile_2_6_to_tile_2_5_1),
		.out_wire_2_2(horizontal_tile_2_6_to_tile_2_5_2),
		.out_wire_2_3(horizontal_tile_2_6_to_tile_2_5_3),
		.in_wire_2_0(horizontal_tile_2_5_to_tile_2_6_0),
		.in_wire_2_1(horizontal_tile_2_5_to_tile_2_6_1),
		.in_wire_2_2(horizontal_tile_2_5_to_tile_2_6_2),
		.in_wire_2_3(horizontal_tile_2_5_to_tile_2_6_3),
		.out_wire_0_0(horizontal_tile_2_6_to_tile_2_7_0),
		.out_wire_0_1(horizontal_tile_2_6_to_tile_2_7_1),
		.out_wire_0_2(horizontal_tile_2_6_to_tile_2_7_2),
		.out_wire_0_3(horizontal_tile_2_6_to_tile_2_7_3),
		.in_wire_0_0(horizontal_tile_2_7_to_tile_2_6_0),
		.in_wire_0_1(horizontal_tile_2_7_to_tile_2_6_1),
		.in_wire_0_2(horizontal_tile_2_7_to_tile_2_6_2),
		.in_wire_0_3(horizontal_tile_2_7_to_tile_2_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(71)
	);

	pe_tile pe_tile_2_7(
		.out_wire_3_0(vertical_tile_2_7_to_tile_1_7_0),
		.out_wire_3_1(vertical_tile_2_7_to_tile_1_7_1),
		.out_wire_3_2(vertical_tile_2_7_to_tile_1_7_2),
		.out_wire_3_3(vertical_tile_2_7_to_tile_1_7_3),
		.in_wire_3_0(vertical_tile_1_7_to_tile_2_7_0),
		.in_wire_3_1(vertical_tile_1_7_to_tile_2_7_1),
		.in_wire_3_2(vertical_tile_1_7_to_tile_2_7_2),
		.in_wire_3_3(vertical_tile_1_7_to_tile_2_7_3),
		.out_wire_1_0(vertical_tile_2_7_to_tile_3_7_0),
		.out_wire_1_1(vertical_tile_2_7_to_tile_3_7_1),
		.out_wire_1_2(vertical_tile_2_7_to_tile_3_7_2),
		.out_wire_1_3(vertical_tile_2_7_to_tile_3_7_3),
		.in_wire_1_0(vertical_tile_3_7_to_tile_2_7_0),
		.in_wire_1_1(vertical_tile_3_7_to_tile_2_7_1),
		.in_wire_1_2(vertical_tile_3_7_to_tile_2_7_2),
		.in_wire_1_3(vertical_tile_3_7_to_tile_2_7_3),
		.out_wire_2_0(horizontal_tile_2_7_to_tile_2_6_0),
		.out_wire_2_1(horizontal_tile_2_7_to_tile_2_6_1),
		.out_wire_2_2(horizontal_tile_2_7_to_tile_2_6_2),
		.out_wire_2_3(horizontal_tile_2_7_to_tile_2_6_3),
		.in_wire_2_0(horizontal_tile_2_6_to_tile_2_7_0),
		.in_wire_2_1(horizontal_tile_2_6_to_tile_2_7_1),
		.in_wire_2_2(horizontal_tile_2_6_to_tile_2_7_2),
		.in_wire_2_3(horizontal_tile_2_6_to_tile_2_7_3),
		.out_wire_0_0(horizontal_tile_2_7_to_tile_2_8_0),
		.out_wire_0_1(horizontal_tile_2_7_to_tile_2_8_1),
		.out_wire_0_2(horizontal_tile_2_7_to_tile_2_8_2),
		.out_wire_0_3(horizontal_tile_2_7_to_tile_2_8_3),
		.in_wire_0_0(horizontal_tile_2_8_to_tile_2_7_0),
		.in_wire_0_1(horizontal_tile_2_8_to_tile_2_7_1),
		.in_wire_0_2(horizontal_tile_2_8_to_tile_2_7_2),
		.in_wire_0_3(horizontal_tile_2_8_to_tile_2_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(72)
	);

	pe_tile pe_tile_2_8(
		.out_wire_3_0(vertical_tile_2_8_to_tile_1_8_0),
		.out_wire_3_1(vertical_tile_2_8_to_tile_1_8_1),
		.out_wire_3_2(vertical_tile_2_8_to_tile_1_8_2),
		.out_wire_3_3(vertical_tile_2_8_to_tile_1_8_3),
		.in_wire_3_0(vertical_tile_1_8_to_tile_2_8_0),
		.in_wire_3_1(vertical_tile_1_8_to_tile_2_8_1),
		.in_wire_3_2(vertical_tile_1_8_to_tile_2_8_2),
		.in_wire_3_3(vertical_tile_1_8_to_tile_2_8_3),
		.out_wire_1_0(vertical_tile_2_8_to_tile_3_8_0),
		.out_wire_1_1(vertical_tile_2_8_to_tile_3_8_1),
		.out_wire_1_2(vertical_tile_2_8_to_tile_3_8_2),
		.out_wire_1_3(vertical_tile_2_8_to_tile_3_8_3),
		.in_wire_1_0(vertical_tile_3_8_to_tile_2_8_0),
		.in_wire_1_1(vertical_tile_3_8_to_tile_2_8_1),
		.in_wire_1_2(vertical_tile_3_8_to_tile_2_8_2),
		.in_wire_1_3(vertical_tile_3_8_to_tile_2_8_3),
		.out_wire_2_0(horizontal_tile_2_8_to_tile_2_7_0),
		.out_wire_2_1(horizontal_tile_2_8_to_tile_2_7_1),
		.out_wire_2_2(horizontal_tile_2_8_to_tile_2_7_2),
		.out_wire_2_3(horizontal_tile_2_8_to_tile_2_7_3),
		.in_wire_2_0(horizontal_tile_2_7_to_tile_2_8_0),
		.in_wire_2_1(horizontal_tile_2_7_to_tile_2_8_1),
		.in_wire_2_2(horizontal_tile_2_7_to_tile_2_8_2),
		.in_wire_2_3(horizontal_tile_2_7_to_tile_2_8_3),
		.out_wire_0_0(horizontal_tile_2_8_to_tile_2_9_0),
		.out_wire_0_1(horizontal_tile_2_8_to_tile_2_9_1),
		.out_wire_0_2(horizontal_tile_2_8_to_tile_2_9_2),
		.out_wire_0_3(horizontal_tile_2_8_to_tile_2_9_3),
		.in_wire_0_0(horizontal_tile_2_9_to_tile_2_8_0),
		.in_wire_0_1(horizontal_tile_2_9_to_tile_2_8_1),
		.in_wire_0_2(horizontal_tile_2_9_to_tile_2_8_2),
		.in_wire_0_3(horizontal_tile_2_9_to_tile_2_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(73)
	);

	pe_tile pe_tile_2_9(
		.out_wire_3_0(vertical_tile_2_9_to_tile_1_9_0),
		.out_wire_3_1(vertical_tile_2_9_to_tile_1_9_1),
		.out_wire_3_2(vertical_tile_2_9_to_tile_1_9_2),
		.out_wire_3_3(vertical_tile_2_9_to_tile_1_9_3),
		.in_wire_3_0(vertical_tile_1_9_to_tile_2_9_0),
		.in_wire_3_1(vertical_tile_1_9_to_tile_2_9_1),
		.in_wire_3_2(vertical_tile_1_9_to_tile_2_9_2),
		.in_wire_3_3(vertical_tile_1_9_to_tile_2_9_3),
		.out_wire_1_0(vertical_tile_2_9_to_tile_3_9_0),
		.out_wire_1_1(vertical_tile_2_9_to_tile_3_9_1),
		.out_wire_1_2(vertical_tile_2_9_to_tile_3_9_2),
		.out_wire_1_3(vertical_tile_2_9_to_tile_3_9_3),
		.in_wire_1_0(vertical_tile_3_9_to_tile_2_9_0),
		.in_wire_1_1(vertical_tile_3_9_to_tile_2_9_1),
		.in_wire_1_2(vertical_tile_3_9_to_tile_2_9_2),
		.in_wire_1_3(vertical_tile_3_9_to_tile_2_9_3),
		.out_wire_2_0(horizontal_tile_2_9_to_tile_2_8_0),
		.out_wire_2_1(horizontal_tile_2_9_to_tile_2_8_1),
		.out_wire_2_2(horizontal_tile_2_9_to_tile_2_8_2),
		.out_wire_2_3(horizontal_tile_2_9_to_tile_2_8_3),
		.in_wire_2_0(horizontal_tile_2_8_to_tile_2_9_0),
		.in_wire_2_1(horizontal_tile_2_8_to_tile_2_9_1),
		.in_wire_2_2(horizontal_tile_2_8_to_tile_2_9_2),
		.in_wire_2_3(horizontal_tile_2_8_to_tile_2_9_3),
		.out_wire_0_0(horizontal_tile_2_9_to_tile_2_10_0),
		.out_wire_0_1(horizontal_tile_2_9_to_tile_2_10_1),
		.out_wire_0_2(horizontal_tile_2_9_to_tile_2_10_2),
		.out_wire_0_3(horizontal_tile_2_9_to_tile_2_10_3),
		.in_wire_0_0(horizontal_tile_2_10_to_tile_2_9_0),
		.in_wire_0_1(horizontal_tile_2_10_to_tile_2_9_1),
		.in_wire_0_2(horizontal_tile_2_10_to_tile_2_9_2),
		.in_wire_0_3(horizontal_tile_2_10_to_tile_2_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(74)
	);

	pe_tile pe_tile_2_10(
		.out_wire_3_0(vertical_tile_2_10_to_tile_1_10_0),
		.out_wire_3_1(vertical_tile_2_10_to_tile_1_10_1),
		.out_wire_3_2(vertical_tile_2_10_to_tile_1_10_2),
		.out_wire_3_3(vertical_tile_2_10_to_tile_1_10_3),
		.in_wire_3_0(vertical_tile_1_10_to_tile_2_10_0),
		.in_wire_3_1(vertical_tile_1_10_to_tile_2_10_1),
		.in_wire_3_2(vertical_tile_1_10_to_tile_2_10_2),
		.in_wire_3_3(vertical_tile_1_10_to_tile_2_10_3),
		.out_wire_1_0(vertical_tile_2_10_to_tile_3_10_0),
		.out_wire_1_1(vertical_tile_2_10_to_tile_3_10_1),
		.out_wire_1_2(vertical_tile_2_10_to_tile_3_10_2),
		.out_wire_1_3(vertical_tile_2_10_to_tile_3_10_3),
		.in_wire_1_0(vertical_tile_3_10_to_tile_2_10_0),
		.in_wire_1_1(vertical_tile_3_10_to_tile_2_10_1),
		.in_wire_1_2(vertical_tile_3_10_to_tile_2_10_2),
		.in_wire_1_3(vertical_tile_3_10_to_tile_2_10_3),
		.out_wire_2_0(horizontal_tile_2_10_to_tile_2_9_0),
		.out_wire_2_1(horizontal_tile_2_10_to_tile_2_9_1),
		.out_wire_2_2(horizontal_tile_2_10_to_tile_2_9_2),
		.out_wire_2_3(horizontal_tile_2_10_to_tile_2_9_3),
		.in_wire_2_0(horizontal_tile_2_9_to_tile_2_10_0),
		.in_wire_2_1(horizontal_tile_2_9_to_tile_2_10_1),
		.in_wire_2_2(horizontal_tile_2_9_to_tile_2_10_2),
		.in_wire_2_3(horizontal_tile_2_9_to_tile_2_10_3),
		.out_wire_0_0(horizontal_tile_2_10_to_tile_2_11_0),
		.out_wire_0_1(horizontal_tile_2_10_to_tile_2_11_1),
		.out_wire_0_2(horizontal_tile_2_10_to_tile_2_11_2),
		.out_wire_0_3(horizontal_tile_2_10_to_tile_2_11_3),
		.in_wire_0_0(horizontal_tile_2_11_to_tile_2_10_0),
		.in_wire_0_1(horizontal_tile_2_11_to_tile_2_10_1),
		.in_wire_0_2(horizontal_tile_2_11_to_tile_2_10_2),
		.in_wire_0_3(horizontal_tile_2_11_to_tile_2_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(75)
	);

	pe_tile pe_tile_2_11(
		.out_wire_3_0(vertical_tile_2_11_to_tile_1_11_0),
		.out_wire_3_1(vertical_tile_2_11_to_tile_1_11_1),
		.out_wire_3_2(vertical_tile_2_11_to_tile_1_11_2),
		.out_wire_3_3(vertical_tile_2_11_to_tile_1_11_3),
		.in_wire_3_0(vertical_tile_1_11_to_tile_2_11_0),
		.in_wire_3_1(vertical_tile_1_11_to_tile_2_11_1),
		.in_wire_3_2(vertical_tile_1_11_to_tile_2_11_2),
		.in_wire_3_3(vertical_tile_1_11_to_tile_2_11_3),
		.out_wire_1_0(vertical_tile_2_11_to_tile_3_11_0),
		.out_wire_1_1(vertical_tile_2_11_to_tile_3_11_1),
		.out_wire_1_2(vertical_tile_2_11_to_tile_3_11_2),
		.out_wire_1_3(vertical_tile_2_11_to_tile_3_11_3),
		.in_wire_1_0(vertical_tile_3_11_to_tile_2_11_0),
		.in_wire_1_1(vertical_tile_3_11_to_tile_2_11_1),
		.in_wire_1_2(vertical_tile_3_11_to_tile_2_11_2),
		.in_wire_1_3(vertical_tile_3_11_to_tile_2_11_3),
		.out_wire_2_0(horizontal_tile_2_11_to_tile_2_10_0),
		.out_wire_2_1(horizontal_tile_2_11_to_tile_2_10_1),
		.out_wire_2_2(horizontal_tile_2_11_to_tile_2_10_2),
		.out_wire_2_3(horizontal_tile_2_11_to_tile_2_10_3),
		.in_wire_2_0(horizontal_tile_2_10_to_tile_2_11_0),
		.in_wire_2_1(horizontal_tile_2_10_to_tile_2_11_1),
		.in_wire_2_2(horizontal_tile_2_10_to_tile_2_11_2),
		.in_wire_2_3(horizontal_tile_2_10_to_tile_2_11_3),
		.out_wire_0_0(horizontal_tile_2_11_to_tile_2_12_0),
		.out_wire_0_1(horizontal_tile_2_11_to_tile_2_12_1),
		.out_wire_0_2(horizontal_tile_2_11_to_tile_2_12_2),
		.out_wire_0_3(horizontal_tile_2_11_to_tile_2_12_3),
		.in_wire_0_0(horizontal_tile_2_12_to_tile_2_11_0),
		.in_wire_0_1(horizontal_tile_2_12_to_tile_2_11_1),
		.in_wire_0_2(horizontal_tile_2_12_to_tile_2_11_2),
		.in_wire_0_3(horizontal_tile_2_12_to_tile_2_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(76)
	);

	pe_tile pe_tile_2_12(
		.out_wire_3_0(vertical_tile_2_12_to_tile_1_12_0),
		.out_wire_3_1(vertical_tile_2_12_to_tile_1_12_1),
		.out_wire_3_2(vertical_tile_2_12_to_tile_1_12_2),
		.out_wire_3_3(vertical_tile_2_12_to_tile_1_12_3),
		.in_wire_3_0(vertical_tile_1_12_to_tile_2_12_0),
		.in_wire_3_1(vertical_tile_1_12_to_tile_2_12_1),
		.in_wire_3_2(vertical_tile_1_12_to_tile_2_12_2),
		.in_wire_3_3(vertical_tile_1_12_to_tile_2_12_3),
		.out_wire_1_0(vertical_tile_2_12_to_tile_3_12_0),
		.out_wire_1_1(vertical_tile_2_12_to_tile_3_12_1),
		.out_wire_1_2(vertical_tile_2_12_to_tile_3_12_2),
		.out_wire_1_3(vertical_tile_2_12_to_tile_3_12_3),
		.in_wire_1_0(vertical_tile_3_12_to_tile_2_12_0),
		.in_wire_1_1(vertical_tile_3_12_to_tile_2_12_1),
		.in_wire_1_2(vertical_tile_3_12_to_tile_2_12_2),
		.in_wire_1_3(vertical_tile_3_12_to_tile_2_12_3),
		.out_wire_2_0(horizontal_tile_2_12_to_tile_2_11_0),
		.out_wire_2_1(horizontal_tile_2_12_to_tile_2_11_1),
		.out_wire_2_2(horizontal_tile_2_12_to_tile_2_11_2),
		.out_wire_2_3(horizontal_tile_2_12_to_tile_2_11_3),
		.in_wire_2_0(horizontal_tile_2_11_to_tile_2_12_0),
		.in_wire_2_1(horizontal_tile_2_11_to_tile_2_12_1),
		.in_wire_2_2(horizontal_tile_2_11_to_tile_2_12_2),
		.in_wire_2_3(horizontal_tile_2_11_to_tile_2_12_3),
		.out_wire_0_0(horizontal_tile_2_12_to_tile_2_13_0),
		.out_wire_0_1(horizontal_tile_2_12_to_tile_2_13_1),
		.out_wire_0_2(horizontal_tile_2_12_to_tile_2_13_2),
		.out_wire_0_3(horizontal_tile_2_12_to_tile_2_13_3),
		.in_wire_0_0(horizontal_tile_2_13_to_tile_2_12_0),
		.in_wire_0_1(horizontal_tile_2_13_to_tile_2_12_1),
		.in_wire_0_2(horizontal_tile_2_13_to_tile_2_12_2),
		.in_wire_0_3(horizontal_tile_2_13_to_tile_2_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(77)
	);

	pe_tile pe_tile_2_13(
		.out_wire_3_0(vertical_tile_2_13_to_tile_1_13_0),
		.out_wire_3_1(vertical_tile_2_13_to_tile_1_13_1),
		.out_wire_3_2(vertical_tile_2_13_to_tile_1_13_2),
		.out_wire_3_3(vertical_tile_2_13_to_tile_1_13_3),
		.in_wire_3_0(vertical_tile_1_13_to_tile_2_13_0),
		.in_wire_3_1(vertical_tile_1_13_to_tile_2_13_1),
		.in_wire_3_2(vertical_tile_1_13_to_tile_2_13_2),
		.in_wire_3_3(vertical_tile_1_13_to_tile_2_13_3),
		.out_wire_1_0(vertical_tile_2_13_to_tile_3_13_0),
		.out_wire_1_1(vertical_tile_2_13_to_tile_3_13_1),
		.out_wire_1_2(vertical_tile_2_13_to_tile_3_13_2),
		.out_wire_1_3(vertical_tile_2_13_to_tile_3_13_3),
		.in_wire_1_0(vertical_tile_3_13_to_tile_2_13_0),
		.in_wire_1_1(vertical_tile_3_13_to_tile_2_13_1),
		.in_wire_1_2(vertical_tile_3_13_to_tile_2_13_2),
		.in_wire_1_3(vertical_tile_3_13_to_tile_2_13_3),
		.out_wire_2_0(horizontal_tile_2_13_to_tile_2_12_0),
		.out_wire_2_1(horizontal_tile_2_13_to_tile_2_12_1),
		.out_wire_2_2(horizontal_tile_2_13_to_tile_2_12_2),
		.out_wire_2_3(horizontal_tile_2_13_to_tile_2_12_3),
		.in_wire_2_0(horizontal_tile_2_12_to_tile_2_13_0),
		.in_wire_2_1(horizontal_tile_2_12_to_tile_2_13_1),
		.in_wire_2_2(horizontal_tile_2_12_to_tile_2_13_2),
		.in_wire_2_3(horizontal_tile_2_12_to_tile_2_13_3),
		.out_wire_0_0(horizontal_tile_2_13_to_tile_2_14_0),
		.out_wire_0_1(horizontal_tile_2_13_to_tile_2_14_1),
		.out_wire_0_2(horizontal_tile_2_13_to_tile_2_14_2),
		.out_wire_0_3(horizontal_tile_2_13_to_tile_2_14_3),
		.in_wire_0_0(horizontal_tile_2_14_to_tile_2_13_0),
		.in_wire_0_1(horizontal_tile_2_14_to_tile_2_13_1),
		.in_wire_0_2(horizontal_tile_2_14_to_tile_2_13_2),
		.in_wire_0_3(horizontal_tile_2_14_to_tile_2_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(78)
	);

	pe_tile pe_tile_2_14(
		.out_wire_3_0(vertical_tile_2_14_to_tile_1_14_0),
		.out_wire_3_1(vertical_tile_2_14_to_tile_1_14_1),
		.out_wire_3_2(vertical_tile_2_14_to_tile_1_14_2),
		.out_wire_3_3(vertical_tile_2_14_to_tile_1_14_3),
		.in_wire_3_0(vertical_tile_1_14_to_tile_2_14_0),
		.in_wire_3_1(vertical_tile_1_14_to_tile_2_14_1),
		.in_wire_3_2(vertical_tile_1_14_to_tile_2_14_2),
		.in_wire_3_3(vertical_tile_1_14_to_tile_2_14_3),
		.out_wire_1_0(vertical_tile_2_14_to_tile_3_14_0),
		.out_wire_1_1(vertical_tile_2_14_to_tile_3_14_1),
		.out_wire_1_2(vertical_tile_2_14_to_tile_3_14_2),
		.out_wire_1_3(vertical_tile_2_14_to_tile_3_14_3),
		.in_wire_1_0(vertical_tile_3_14_to_tile_2_14_0),
		.in_wire_1_1(vertical_tile_3_14_to_tile_2_14_1),
		.in_wire_1_2(vertical_tile_3_14_to_tile_2_14_2),
		.in_wire_1_3(vertical_tile_3_14_to_tile_2_14_3),
		.out_wire_2_0(horizontal_tile_2_14_to_tile_2_13_0),
		.out_wire_2_1(horizontal_tile_2_14_to_tile_2_13_1),
		.out_wire_2_2(horizontal_tile_2_14_to_tile_2_13_2),
		.out_wire_2_3(horizontal_tile_2_14_to_tile_2_13_3),
		.in_wire_2_0(horizontal_tile_2_13_to_tile_2_14_0),
		.in_wire_2_1(horizontal_tile_2_13_to_tile_2_14_1),
		.in_wire_2_2(horizontal_tile_2_13_to_tile_2_14_2),
		.in_wire_2_3(horizontal_tile_2_13_to_tile_2_14_3),
		.out_wire_0_0(horizontal_tile_2_14_to_tile_2_15_0),
		.out_wire_0_1(horizontal_tile_2_14_to_tile_2_15_1),
		.out_wire_0_2(horizontal_tile_2_14_to_tile_2_15_2),
		.out_wire_0_3(horizontal_tile_2_14_to_tile_2_15_3),
		.in_wire_0_0(horizontal_tile_2_15_to_tile_2_14_0),
		.in_wire_0_1(horizontal_tile_2_15_to_tile_2_14_1),
		.in_wire_0_2(horizontal_tile_2_15_to_tile_2_14_2),
		.in_wire_0_3(horizontal_tile_2_15_to_tile_2_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(79)
	);

	pe_tile pe_tile_2_15(
		.out_wire_3_0(vertical_tile_2_15_to_tile_1_15_0),
		.out_wire_3_1(vertical_tile_2_15_to_tile_1_15_1),
		.out_wire_3_2(vertical_tile_2_15_to_tile_1_15_2),
		.out_wire_3_3(vertical_tile_2_15_to_tile_1_15_3),
		.in_wire_3_0(vertical_tile_1_15_to_tile_2_15_0),
		.in_wire_3_1(vertical_tile_1_15_to_tile_2_15_1),
		.in_wire_3_2(vertical_tile_1_15_to_tile_2_15_2),
		.in_wire_3_3(vertical_tile_1_15_to_tile_2_15_3),
		.out_wire_1_0(vertical_tile_2_15_to_tile_3_15_0),
		.out_wire_1_1(vertical_tile_2_15_to_tile_3_15_1),
		.out_wire_1_2(vertical_tile_2_15_to_tile_3_15_2),
		.out_wire_1_3(vertical_tile_2_15_to_tile_3_15_3),
		.in_wire_1_0(vertical_tile_3_15_to_tile_2_15_0),
		.in_wire_1_1(vertical_tile_3_15_to_tile_2_15_1),
		.in_wire_1_2(vertical_tile_3_15_to_tile_2_15_2),
		.in_wire_1_3(vertical_tile_3_15_to_tile_2_15_3),
		.out_wire_2_0(horizontal_tile_2_15_to_tile_2_14_0),
		.out_wire_2_1(horizontal_tile_2_15_to_tile_2_14_1),
		.out_wire_2_2(horizontal_tile_2_15_to_tile_2_14_2),
		.out_wire_2_3(horizontal_tile_2_15_to_tile_2_14_3),
		.in_wire_2_0(horizontal_tile_2_14_to_tile_2_15_0),
		.in_wire_2_1(horizontal_tile_2_14_to_tile_2_15_1),
		.in_wire_2_2(horizontal_tile_2_14_to_tile_2_15_2),
		.in_wire_2_3(horizontal_tile_2_14_to_tile_2_15_3),
		.out_wire_0_0(horizontal_tile_2_15_to_tile_2_16_0),
		.out_wire_0_1(horizontal_tile_2_15_to_tile_2_16_1),
		.out_wire_0_2(horizontal_tile_2_15_to_tile_2_16_2),
		.out_wire_0_3(horizontal_tile_2_15_to_tile_2_16_3),
		.in_wire_0_0(horizontal_tile_2_16_to_tile_2_15_0),
		.in_wire_0_1(horizontal_tile_2_16_to_tile_2_15_1),
		.in_wire_0_2(horizontal_tile_2_16_to_tile_2_15_2),
		.in_wire_0_3(horizontal_tile_2_16_to_tile_2_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(80)
	);

	pe_tile pe_tile_2_16(
		.out_wire_3_0(vertical_tile_2_16_to_tile_1_16_0),
		.out_wire_3_1(vertical_tile_2_16_to_tile_1_16_1),
		.out_wire_3_2(vertical_tile_2_16_to_tile_1_16_2),
		.out_wire_3_3(vertical_tile_2_16_to_tile_1_16_3),
		.in_wire_3_0(vertical_tile_1_16_to_tile_2_16_0),
		.in_wire_3_1(vertical_tile_1_16_to_tile_2_16_1),
		.in_wire_3_2(vertical_tile_1_16_to_tile_2_16_2),
		.in_wire_3_3(vertical_tile_1_16_to_tile_2_16_3),
		.out_wire_1_0(vertical_tile_2_16_to_tile_3_16_0),
		.out_wire_1_1(vertical_tile_2_16_to_tile_3_16_1),
		.out_wire_1_2(vertical_tile_2_16_to_tile_3_16_2),
		.out_wire_1_3(vertical_tile_2_16_to_tile_3_16_3),
		.in_wire_1_0(vertical_tile_3_16_to_tile_2_16_0),
		.in_wire_1_1(vertical_tile_3_16_to_tile_2_16_1),
		.in_wire_1_2(vertical_tile_3_16_to_tile_2_16_2),
		.in_wire_1_3(vertical_tile_3_16_to_tile_2_16_3),
		.out_wire_2_0(horizontal_tile_2_16_to_tile_2_15_0),
		.out_wire_2_1(horizontal_tile_2_16_to_tile_2_15_1),
		.out_wire_2_2(horizontal_tile_2_16_to_tile_2_15_2),
		.out_wire_2_3(horizontal_tile_2_16_to_tile_2_15_3),
		.in_wire_2_0(horizontal_tile_2_15_to_tile_2_16_0),
		.in_wire_2_1(horizontal_tile_2_15_to_tile_2_16_1),
		.in_wire_2_2(horizontal_tile_2_15_to_tile_2_16_2),
		.in_wire_2_3(horizontal_tile_2_15_to_tile_2_16_3),
		.out_wire_0_0(horizontal_tile_2_16_to_tile_2_17_0),
		.out_wire_0_1(horizontal_tile_2_16_to_tile_2_17_1),
		.out_wire_0_2(horizontal_tile_2_16_to_tile_2_17_2),
		.out_wire_0_3(horizontal_tile_2_16_to_tile_2_17_3),
		.in_wire_0_0(horizontal_tile_2_17_to_tile_2_16_0),
		.in_wire_0_1(horizontal_tile_2_17_to_tile_2_16_1),
		.in_wire_0_2(horizontal_tile_2_17_to_tile_2_16_2),
		.in_wire_0_3(horizontal_tile_2_17_to_tile_2_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(81)
	);

	pe_tile pe_tile_2_17(
		.out_wire_3_0(vertical_tile_2_17_to_tile_1_17_0),
		.out_wire_3_1(vertical_tile_2_17_to_tile_1_17_1),
		.out_wire_3_2(vertical_tile_2_17_to_tile_1_17_2),
		.out_wire_3_3(vertical_tile_2_17_to_tile_1_17_3),
		.in_wire_3_0(vertical_tile_1_17_to_tile_2_17_0),
		.in_wire_3_1(vertical_tile_1_17_to_tile_2_17_1),
		.in_wire_3_2(vertical_tile_1_17_to_tile_2_17_2),
		.in_wire_3_3(vertical_tile_1_17_to_tile_2_17_3),
		.out_wire_1_0(vertical_tile_2_17_to_tile_3_17_0),
		.out_wire_1_1(vertical_tile_2_17_to_tile_3_17_1),
		.out_wire_1_2(vertical_tile_2_17_to_tile_3_17_2),
		.out_wire_1_3(vertical_tile_2_17_to_tile_3_17_3),
		.in_wire_1_0(vertical_tile_3_17_to_tile_2_17_0),
		.in_wire_1_1(vertical_tile_3_17_to_tile_2_17_1),
		.in_wire_1_2(vertical_tile_3_17_to_tile_2_17_2),
		.in_wire_1_3(vertical_tile_3_17_to_tile_2_17_3),
		.out_wire_2_0(horizontal_tile_2_17_to_tile_2_16_0),
		.out_wire_2_1(horizontal_tile_2_17_to_tile_2_16_1),
		.out_wire_2_2(horizontal_tile_2_17_to_tile_2_16_2),
		.out_wire_2_3(horizontal_tile_2_17_to_tile_2_16_3),
		.in_wire_2_0(horizontal_tile_2_16_to_tile_2_17_0),
		.in_wire_2_1(horizontal_tile_2_16_to_tile_2_17_1),
		.in_wire_2_2(horizontal_tile_2_16_to_tile_2_17_2),
		.in_wire_2_3(horizontal_tile_2_16_to_tile_2_17_3),
		.out_wire_0_0(horizontal_tile_2_17_to_tile_2_18_0),
		.out_wire_0_1(horizontal_tile_2_17_to_tile_2_18_1),
		.out_wire_0_2(horizontal_tile_2_17_to_tile_2_18_2),
		.out_wire_0_3(horizontal_tile_2_17_to_tile_2_18_3),
		.in_wire_0_0(horizontal_tile_2_18_to_tile_2_17_0),
		.in_wire_0_1(horizontal_tile_2_18_to_tile_2_17_1),
		.in_wire_0_2(horizontal_tile_2_18_to_tile_2_17_2),
		.in_wire_0_3(horizontal_tile_2_18_to_tile_2_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(82)
	);

	pe_tile pe_tile_2_18(
		.out_wire_3_0(vertical_tile_2_18_to_tile_1_18_0),
		.out_wire_3_1(vertical_tile_2_18_to_tile_1_18_1),
		.out_wire_3_2(vertical_tile_2_18_to_tile_1_18_2),
		.out_wire_3_3(vertical_tile_2_18_to_tile_1_18_3),
		.in_wire_3_0(vertical_tile_1_18_to_tile_2_18_0),
		.in_wire_3_1(vertical_tile_1_18_to_tile_2_18_1),
		.in_wire_3_2(vertical_tile_1_18_to_tile_2_18_2),
		.in_wire_3_3(vertical_tile_1_18_to_tile_2_18_3),
		.out_wire_1_0(vertical_tile_2_18_to_tile_3_18_0),
		.out_wire_1_1(vertical_tile_2_18_to_tile_3_18_1),
		.out_wire_1_2(vertical_tile_2_18_to_tile_3_18_2),
		.out_wire_1_3(vertical_tile_2_18_to_tile_3_18_3),
		.in_wire_1_0(vertical_tile_3_18_to_tile_2_18_0),
		.in_wire_1_1(vertical_tile_3_18_to_tile_2_18_1),
		.in_wire_1_2(vertical_tile_3_18_to_tile_2_18_2),
		.in_wire_1_3(vertical_tile_3_18_to_tile_2_18_3),
		.out_wire_2_0(horizontal_tile_2_18_to_tile_2_17_0),
		.out_wire_2_1(horizontal_tile_2_18_to_tile_2_17_1),
		.out_wire_2_2(horizontal_tile_2_18_to_tile_2_17_2),
		.out_wire_2_3(horizontal_tile_2_18_to_tile_2_17_3),
		.in_wire_2_0(horizontal_tile_2_17_to_tile_2_18_0),
		.in_wire_2_1(horizontal_tile_2_17_to_tile_2_18_1),
		.in_wire_2_2(horizontal_tile_2_17_to_tile_2_18_2),
		.in_wire_2_3(horizontal_tile_2_17_to_tile_2_18_3),
		.out_wire_0_0(horizontal_tile_2_18_to_tile_2_19_0),
		.out_wire_0_1(horizontal_tile_2_18_to_tile_2_19_1),
		.out_wire_0_2(horizontal_tile_2_18_to_tile_2_19_2),
		.out_wire_0_3(horizontal_tile_2_18_to_tile_2_19_3),
		.in_wire_0_0(horizontal_tile_2_19_to_tile_2_18_0),
		.in_wire_0_1(horizontal_tile_2_19_to_tile_2_18_1),
		.in_wire_0_2(horizontal_tile_2_19_to_tile_2_18_2),
		.in_wire_0_3(horizontal_tile_2_19_to_tile_2_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(83)
	);

	pe_tile pe_tile_2_19(
		.out_wire_3_0(vertical_tile_2_19_to_tile_1_19_0),
		.out_wire_3_1(vertical_tile_2_19_to_tile_1_19_1),
		.out_wire_3_2(vertical_tile_2_19_to_tile_1_19_2),
		.out_wire_3_3(vertical_tile_2_19_to_tile_1_19_3),
		.in_wire_3_0(vertical_tile_1_19_to_tile_2_19_0),
		.in_wire_3_1(vertical_tile_1_19_to_tile_2_19_1),
		.in_wire_3_2(vertical_tile_1_19_to_tile_2_19_2),
		.in_wire_3_3(vertical_tile_1_19_to_tile_2_19_3),
		.out_wire_1_0(vertical_tile_2_19_to_tile_3_19_0),
		.out_wire_1_1(vertical_tile_2_19_to_tile_3_19_1),
		.out_wire_1_2(vertical_tile_2_19_to_tile_3_19_2),
		.out_wire_1_3(vertical_tile_2_19_to_tile_3_19_3),
		.in_wire_1_0(vertical_tile_3_19_to_tile_2_19_0),
		.in_wire_1_1(vertical_tile_3_19_to_tile_2_19_1),
		.in_wire_1_2(vertical_tile_3_19_to_tile_2_19_2),
		.in_wire_1_3(vertical_tile_3_19_to_tile_2_19_3),
		.out_wire_2_0(horizontal_tile_2_19_to_tile_2_18_0),
		.out_wire_2_1(horizontal_tile_2_19_to_tile_2_18_1),
		.out_wire_2_2(horizontal_tile_2_19_to_tile_2_18_2),
		.out_wire_2_3(horizontal_tile_2_19_to_tile_2_18_3),
		.in_wire_2_0(horizontal_tile_2_18_to_tile_2_19_0),
		.in_wire_2_1(horizontal_tile_2_18_to_tile_2_19_1),
		.in_wire_2_2(horizontal_tile_2_18_to_tile_2_19_2),
		.in_wire_2_3(horizontal_tile_2_18_to_tile_2_19_3),
		.out_wire_0_0(horizontal_tile_2_19_to_tile_2_20_0),
		.out_wire_0_1(horizontal_tile_2_19_to_tile_2_20_1),
		.out_wire_0_2(horizontal_tile_2_19_to_tile_2_20_2),
		.out_wire_0_3(horizontal_tile_2_19_to_tile_2_20_3),
		.in_wire_0_0(horizontal_tile_2_20_to_tile_2_19_0),
		.in_wire_0_1(horizontal_tile_2_20_to_tile_2_19_1),
		.in_wire_0_2(horizontal_tile_2_20_to_tile_2_19_2),
		.in_wire_0_3(horizontal_tile_2_20_to_tile_2_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(84)
	);

	pe_tile pe_tile_2_20(
		.out_wire_3_0(vertical_tile_2_20_to_tile_1_20_0),
		.out_wire_3_1(vertical_tile_2_20_to_tile_1_20_1),
		.out_wire_3_2(vertical_tile_2_20_to_tile_1_20_2),
		.out_wire_3_3(vertical_tile_2_20_to_tile_1_20_3),
		.in_wire_3_0(vertical_tile_1_20_to_tile_2_20_0),
		.in_wire_3_1(vertical_tile_1_20_to_tile_2_20_1),
		.in_wire_3_2(vertical_tile_1_20_to_tile_2_20_2),
		.in_wire_3_3(vertical_tile_1_20_to_tile_2_20_3),
		.out_wire_1_0(vertical_tile_2_20_to_tile_3_20_0),
		.out_wire_1_1(vertical_tile_2_20_to_tile_3_20_1),
		.out_wire_1_2(vertical_tile_2_20_to_tile_3_20_2),
		.out_wire_1_3(vertical_tile_2_20_to_tile_3_20_3),
		.in_wire_1_0(vertical_tile_3_20_to_tile_2_20_0),
		.in_wire_1_1(vertical_tile_3_20_to_tile_2_20_1),
		.in_wire_1_2(vertical_tile_3_20_to_tile_2_20_2),
		.in_wire_1_3(vertical_tile_3_20_to_tile_2_20_3),
		.out_wire_2_0(horizontal_tile_2_20_to_tile_2_19_0),
		.out_wire_2_1(horizontal_tile_2_20_to_tile_2_19_1),
		.out_wire_2_2(horizontal_tile_2_20_to_tile_2_19_2),
		.out_wire_2_3(horizontal_tile_2_20_to_tile_2_19_3),
		.in_wire_2_0(horizontal_tile_2_19_to_tile_2_20_0),
		.in_wire_2_1(horizontal_tile_2_19_to_tile_2_20_1),
		.in_wire_2_2(horizontal_tile_2_19_to_tile_2_20_2),
		.in_wire_2_3(horizontal_tile_2_19_to_tile_2_20_3),
		.out_wire_0_0(horizontal_tile_2_20_to_tile_2_21_0),
		.out_wire_0_1(horizontal_tile_2_20_to_tile_2_21_1),
		.out_wire_0_2(horizontal_tile_2_20_to_tile_2_21_2),
		.out_wire_0_3(horizontal_tile_2_20_to_tile_2_21_3),
		.in_wire_0_0(horizontal_tile_2_21_to_tile_2_20_0),
		.in_wire_0_1(horizontal_tile_2_21_to_tile_2_20_1),
		.in_wire_0_2(horizontal_tile_2_21_to_tile_2_20_2),
		.in_wire_0_3(horizontal_tile_2_21_to_tile_2_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(85)
	);

	pe_tile pe_tile_2_21(
		.out_wire_3_0(vertical_tile_2_21_to_tile_1_21_0),
		.out_wire_3_1(vertical_tile_2_21_to_tile_1_21_1),
		.out_wire_3_2(vertical_tile_2_21_to_tile_1_21_2),
		.out_wire_3_3(vertical_tile_2_21_to_tile_1_21_3),
		.in_wire_3_0(vertical_tile_1_21_to_tile_2_21_0),
		.in_wire_3_1(vertical_tile_1_21_to_tile_2_21_1),
		.in_wire_3_2(vertical_tile_1_21_to_tile_2_21_2),
		.in_wire_3_3(vertical_tile_1_21_to_tile_2_21_3),
		.out_wire_1_0(vertical_tile_2_21_to_tile_3_21_0),
		.out_wire_1_1(vertical_tile_2_21_to_tile_3_21_1),
		.out_wire_1_2(vertical_tile_2_21_to_tile_3_21_2),
		.out_wire_1_3(vertical_tile_2_21_to_tile_3_21_3),
		.in_wire_1_0(vertical_tile_3_21_to_tile_2_21_0),
		.in_wire_1_1(vertical_tile_3_21_to_tile_2_21_1),
		.in_wire_1_2(vertical_tile_3_21_to_tile_2_21_2),
		.in_wire_1_3(vertical_tile_3_21_to_tile_2_21_3),
		.out_wire_2_0(horizontal_tile_2_21_to_tile_2_20_0),
		.out_wire_2_1(horizontal_tile_2_21_to_tile_2_20_1),
		.out_wire_2_2(horizontal_tile_2_21_to_tile_2_20_2),
		.out_wire_2_3(horizontal_tile_2_21_to_tile_2_20_3),
		.in_wire_2_0(horizontal_tile_2_20_to_tile_2_21_0),
		.in_wire_2_1(horizontal_tile_2_20_to_tile_2_21_1),
		.in_wire_2_2(horizontal_tile_2_20_to_tile_2_21_2),
		.in_wire_2_3(horizontal_tile_2_20_to_tile_2_21_3),
		.out_wire_0_0(horizontal_tile_2_21_to_tile_2_22_0),
		.out_wire_0_1(horizontal_tile_2_21_to_tile_2_22_1),
		.out_wire_0_2(horizontal_tile_2_21_to_tile_2_22_2),
		.out_wire_0_3(horizontal_tile_2_21_to_tile_2_22_3),
		.in_wire_0_0(horizontal_tile_2_22_to_tile_2_21_0),
		.in_wire_0_1(horizontal_tile_2_22_to_tile_2_21_1),
		.in_wire_0_2(horizontal_tile_2_22_to_tile_2_21_2),
		.in_wire_0_3(horizontal_tile_2_22_to_tile_2_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(86)
	);

	pe_tile pe_tile_2_22(
		.out_wire_3_0(vertical_tile_2_22_to_tile_1_22_0),
		.out_wire_3_1(vertical_tile_2_22_to_tile_1_22_1),
		.out_wire_3_2(vertical_tile_2_22_to_tile_1_22_2),
		.out_wire_3_3(vertical_tile_2_22_to_tile_1_22_3),
		.in_wire_3_0(vertical_tile_1_22_to_tile_2_22_0),
		.in_wire_3_1(vertical_tile_1_22_to_tile_2_22_1),
		.in_wire_3_2(vertical_tile_1_22_to_tile_2_22_2),
		.in_wire_3_3(vertical_tile_1_22_to_tile_2_22_3),
		.out_wire_1_0(vertical_tile_2_22_to_tile_3_22_0),
		.out_wire_1_1(vertical_tile_2_22_to_tile_3_22_1),
		.out_wire_1_2(vertical_tile_2_22_to_tile_3_22_2),
		.out_wire_1_3(vertical_tile_2_22_to_tile_3_22_3),
		.in_wire_1_0(vertical_tile_3_22_to_tile_2_22_0),
		.in_wire_1_1(vertical_tile_3_22_to_tile_2_22_1),
		.in_wire_1_2(vertical_tile_3_22_to_tile_2_22_2),
		.in_wire_1_3(vertical_tile_3_22_to_tile_2_22_3),
		.out_wire_2_0(horizontal_tile_2_22_to_tile_2_21_0),
		.out_wire_2_1(horizontal_tile_2_22_to_tile_2_21_1),
		.out_wire_2_2(horizontal_tile_2_22_to_tile_2_21_2),
		.out_wire_2_3(horizontal_tile_2_22_to_tile_2_21_3),
		.in_wire_2_0(horizontal_tile_2_21_to_tile_2_22_0),
		.in_wire_2_1(horizontal_tile_2_21_to_tile_2_22_1),
		.in_wire_2_2(horizontal_tile_2_21_to_tile_2_22_2),
		.in_wire_2_3(horizontal_tile_2_21_to_tile_2_22_3),
		.out_wire_0_0(horizontal_tile_2_22_to_tile_2_23_0),
		.out_wire_0_1(horizontal_tile_2_22_to_tile_2_23_1),
		.out_wire_0_2(horizontal_tile_2_22_to_tile_2_23_2),
		.out_wire_0_3(horizontal_tile_2_22_to_tile_2_23_3),
		.in_wire_0_0(horizontal_tile_2_23_to_tile_2_22_0),
		.in_wire_0_1(horizontal_tile_2_23_to_tile_2_22_1),
		.in_wire_0_2(horizontal_tile_2_23_to_tile_2_22_2),
		.in_wire_0_3(horizontal_tile_2_23_to_tile_2_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(87)
	);

	pe_tile pe_tile_2_23(
		.out_wire_3_0(vertical_tile_2_23_to_tile_1_23_0),
		.out_wire_3_1(vertical_tile_2_23_to_tile_1_23_1),
		.out_wire_3_2(vertical_tile_2_23_to_tile_1_23_2),
		.out_wire_3_3(vertical_tile_2_23_to_tile_1_23_3),
		.in_wire_3_0(vertical_tile_1_23_to_tile_2_23_0),
		.in_wire_3_1(vertical_tile_1_23_to_tile_2_23_1),
		.in_wire_3_2(vertical_tile_1_23_to_tile_2_23_2),
		.in_wire_3_3(vertical_tile_1_23_to_tile_2_23_3),
		.out_wire_1_0(vertical_tile_2_23_to_tile_3_23_0),
		.out_wire_1_1(vertical_tile_2_23_to_tile_3_23_1),
		.out_wire_1_2(vertical_tile_2_23_to_tile_3_23_2),
		.out_wire_1_3(vertical_tile_2_23_to_tile_3_23_3),
		.in_wire_1_0(vertical_tile_3_23_to_tile_2_23_0),
		.in_wire_1_1(vertical_tile_3_23_to_tile_2_23_1),
		.in_wire_1_2(vertical_tile_3_23_to_tile_2_23_2),
		.in_wire_1_3(vertical_tile_3_23_to_tile_2_23_3),
		.out_wire_2_0(horizontal_tile_2_23_to_tile_2_22_0),
		.out_wire_2_1(horizontal_tile_2_23_to_tile_2_22_1),
		.out_wire_2_2(horizontal_tile_2_23_to_tile_2_22_2),
		.out_wire_2_3(horizontal_tile_2_23_to_tile_2_22_3),
		.in_wire_2_0(horizontal_tile_2_22_to_tile_2_23_0),
		.in_wire_2_1(horizontal_tile_2_22_to_tile_2_23_1),
		.in_wire_2_2(horizontal_tile_2_22_to_tile_2_23_2),
		.in_wire_2_3(horizontal_tile_2_22_to_tile_2_23_3),
		.out_wire_0_0(horizontal_tile_2_23_to_tile_2_24_0),
		.out_wire_0_1(horizontal_tile_2_23_to_tile_2_24_1),
		.out_wire_0_2(horizontal_tile_2_23_to_tile_2_24_2),
		.out_wire_0_3(horizontal_tile_2_23_to_tile_2_24_3),
		.in_wire_0_0(horizontal_tile_2_24_to_tile_2_23_0),
		.in_wire_0_1(horizontal_tile_2_24_to_tile_2_23_1),
		.in_wire_0_2(horizontal_tile_2_24_to_tile_2_23_2),
		.in_wire_0_3(horizontal_tile_2_24_to_tile_2_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(88)
	);

	pe_tile pe_tile_2_24(
		.out_wire_3_0(vertical_tile_2_24_to_tile_1_24_0),
		.out_wire_3_1(vertical_tile_2_24_to_tile_1_24_1),
		.out_wire_3_2(vertical_tile_2_24_to_tile_1_24_2),
		.out_wire_3_3(vertical_tile_2_24_to_tile_1_24_3),
		.in_wire_3_0(vertical_tile_1_24_to_tile_2_24_0),
		.in_wire_3_1(vertical_tile_1_24_to_tile_2_24_1),
		.in_wire_3_2(vertical_tile_1_24_to_tile_2_24_2),
		.in_wire_3_3(vertical_tile_1_24_to_tile_2_24_3),
		.out_wire_1_0(vertical_tile_2_24_to_tile_3_24_0),
		.out_wire_1_1(vertical_tile_2_24_to_tile_3_24_1),
		.out_wire_1_2(vertical_tile_2_24_to_tile_3_24_2),
		.out_wire_1_3(vertical_tile_2_24_to_tile_3_24_3),
		.in_wire_1_0(vertical_tile_3_24_to_tile_2_24_0),
		.in_wire_1_1(vertical_tile_3_24_to_tile_2_24_1),
		.in_wire_1_2(vertical_tile_3_24_to_tile_2_24_2),
		.in_wire_1_3(vertical_tile_3_24_to_tile_2_24_3),
		.out_wire_2_0(horizontal_tile_2_24_to_tile_2_23_0),
		.out_wire_2_1(horizontal_tile_2_24_to_tile_2_23_1),
		.out_wire_2_2(horizontal_tile_2_24_to_tile_2_23_2),
		.out_wire_2_3(horizontal_tile_2_24_to_tile_2_23_3),
		.in_wire_2_0(horizontal_tile_2_23_to_tile_2_24_0),
		.in_wire_2_1(horizontal_tile_2_23_to_tile_2_24_1),
		.in_wire_2_2(horizontal_tile_2_23_to_tile_2_24_2),
		.in_wire_2_3(horizontal_tile_2_23_to_tile_2_24_3),
		.out_wire_0_0(horizontal_tile_2_24_to_tile_2_25_0),
		.out_wire_0_1(horizontal_tile_2_24_to_tile_2_25_1),
		.out_wire_0_2(horizontal_tile_2_24_to_tile_2_25_2),
		.out_wire_0_3(horizontal_tile_2_24_to_tile_2_25_3),
		.in_wire_0_0(horizontal_tile_2_25_to_tile_2_24_0),
		.in_wire_0_1(horizontal_tile_2_25_to_tile_2_24_1),
		.in_wire_0_2(horizontal_tile_2_25_to_tile_2_24_2),
		.in_wire_0_3(horizontal_tile_2_25_to_tile_2_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(89)
	);

	pe_tile pe_tile_2_25(
		.out_wire_3_0(vertical_tile_2_25_to_tile_1_25_0),
		.out_wire_3_1(vertical_tile_2_25_to_tile_1_25_1),
		.out_wire_3_2(vertical_tile_2_25_to_tile_1_25_2),
		.out_wire_3_3(vertical_tile_2_25_to_tile_1_25_3),
		.in_wire_3_0(vertical_tile_1_25_to_tile_2_25_0),
		.in_wire_3_1(vertical_tile_1_25_to_tile_2_25_1),
		.in_wire_3_2(vertical_tile_1_25_to_tile_2_25_2),
		.in_wire_3_3(vertical_tile_1_25_to_tile_2_25_3),
		.out_wire_1_0(vertical_tile_2_25_to_tile_3_25_0),
		.out_wire_1_1(vertical_tile_2_25_to_tile_3_25_1),
		.out_wire_1_2(vertical_tile_2_25_to_tile_3_25_2),
		.out_wire_1_3(vertical_tile_2_25_to_tile_3_25_3),
		.in_wire_1_0(vertical_tile_3_25_to_tile_2_25_0),
		.in_wire_1_1(vertical_tile_3_25_to_tile_2_25_1),
		.in_wire_1_2(vertical_tile_3_25_to_tile_2_25_2),
		.in_wire_1_3(vertical_tile_3_25_to_tile_2_25_3),
		.out_wire_2_0(horizontal_tile_2_25_to_tile_2_24_0),
		.out_wire_2_1(horizontal_tile_2_25_to_tile_2_24_1),
		.out_wire_2_2(horizontal_tile_2_25_to_tile_2_24_2),
		.out_wire_2_3(horizontal_tile_2_25_to_tile_2_24_3),
		.in_wire_2_0(horizontal_tile_2_24_to_tile_2_25_0),
		.in_wire_2_1(horizontal_tile_2_24_to_tile_2_25_1),
		.in_wire_2_2(horizontal_tile_2_24_to_tile_2_25_2),
		.in_wire_2_3(horizontal_tile_2_24_to_tile_2_25_3),
		.out_wire_0_0(horizontal_tile_2_25_to_tile_2_26_0),
		.out_wire_0_1(horizontal_tile_2_25_to_tile_2_26_1),
		.out_wire_0_2(horizontal_tile_2_25_to_tile_2_26_2),
		.out_wire_0_3(horizontal_tile_2_25_to_tile_2_26_3),
		.in_wire_0_0(horizontal_tile_2_26_to_tile_2_25_0),
		.in_wire_0_1(horizontal_tile_2_26_to_tile_2_25_1),
		.in_wire_0_2(horizontal_tile_2_26_to_tile_2_25_2),
		.in_wire_0_3(horizontal_tile_2_26_to_tile_2_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(90)
	);

	pe_tile pe_tile_2_26(
		.out_wire_3_0(vertical_tile_2_26_to_tile_1_26_0),
		.out_wire_3_1(vertical_tile_2_26_to_tile_1_26_1),
		.out_wire_3_2(vertical_tile_2_26_to_tile_1_26_2),
		.out_wire_3_3(vertical_tile_2_26_to_tile_1_26_3),
		.in_wire_3_0(vertical_tile_1_26_to_tile_2_26_0),
		.in_wire_3_1(vertical_tile_1_26_to_tile_2_26_1),
		.in_wire_3_2(vertical_tile_1_26_to_tile_2_26_2),
		.in_wire_3_3(vertical_tile_1_26_to_tile_2_26_3),
		.out_wire_1_0(vertical_tile_2_26_to_tile_3_26_0),
		.out_wire_1_1(vertical_tile_2_26_to_tile_3_26_1),
		.out_wire_1_2(vertical_tile_2_26_to_tile_3_26_2),
		.out_wire_1_3(vertical_tile_2_26_to_tile_3_26_3),
		.in_wire_1_0(vertical_tile_3_26_to_tile_2_26_0),
		.in_wire_1_1(vertical_tile_3_26_to_tile_2_26_1),
		.in_wire_1_2(vertical_tile_3_26_to_tile_2_26_2),
		.in_wire_1_3(vertical_tile_3_26_to_tile_2_26_3),
		.out_wire_2_0(horizontal_tile_2_26_to_tile_2_25_0),
		.out_wire_2_1(horizontal_tile_2_26_to_tile_2_25_1),
		.out_wire_2_2(horizontal_tile_2_26_to_tile_2_25_2),
		.out_wire_2_3(horizontal_tile_2_26_to_tile_2_25_3),
		.in_wire_2_0(horizontal_tile_2_25_to_tile_2_26_0),
		.in_wire_2_1(horizontal_tile_2_25_to_tile_2_26_1),
		.in_wire_2_2(horizontal_tile_2_25_to_tile_2_26_2),
		.in_wire_2_3(horizontal_tile_2_25_to_tile_2_26_3),
		.out_wire_0_0(horizontal_tile_2_26_to_tile_2_27_0),
		.out_wire_0_1(horizontal_tile_2_26_to_tile_2_27_1),
		.out_wire_0_2(horizontal_tile_2_26_to_tile_2_27_2),
		.out_wire_0_3(horizontal_tile_2_26_to_tile_2_27_3),
		.in_wire_0_0(horizontal_tile_2_27_to_tile_2_26_0),
		.in_wire_0_1(horizontal_tile_2_27_to_tile_2_26_1),
		.in_wire_0_2(horizontal_tile_2_27_to_tile_2_26_2),
		.in_wire_0_3(horizontal_tile_2_27_to_tile_2_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(91)
	);

	pe_tile pe_tile_2_27(
		.out_wire_3_0(vertical_tile_2_27_to_tile_1_27_0),
		.out_wire_3_1(vertical_tile_2_27_to_tile_1_27_1),
		.out_wire_3_2(vertical_tile_2_27_to_tile_1_27_2),
		.out_wire_3_3(vertical_tile_2_27_to_tile_1_27_3),
		.in_wire_3_0(vertical_tile_1_27_to_tile_2_27_0),
		.in_wire_3_1(vertical_tile_1_27_to_tile_2_27_1),
		.in_wire_3_2(vertical_tile_1_27_to_tile_2_27_2),
		.in_wire_3_3(vertical_tile_1_27_to_tile_2_27_3),
		.out_wire_1_0(vertical_tile_2_27_to_tile_3_27_0),
		.out_wire_1_1(vertical_tile_2_27_to_tile_3_27_1),
		.out_wire_1_2(vertical_tile_2_27_to_tile_3_27_2),
		.out_wire_1_3(vertical_tile_2_27_to_tile_3_27_3),
		.in_wire_1_0(vertical_tile_3_27_to_tile_2_27_0),
		.in_wire_1_1(vertical_tile_3_27_to_tile_2_27_1),
		.in_wire_1_2(vertical_tile_3_27_to_tile_2_27_2),
		.in_wire_1_3(vertical_tile_3_27_to_tile_2_27_3),
		.out_wire_2_0(horizontal_tile_2_27_to_tile_2_26_0),
		.out_wire_2_1(horizontal_tile_2_27_to_tile_2_26_1),
		.out_wire_2_2(horizontal_tile_2_27_to_tile_2_26_2),
		.out_wire_2_3(horizontal_tile_2_27_to_tile_2_26_3),
		.in_wire_2_0(horizontal_tile_2_26_to_tile_2_27_0),
		.in_wire_2_1(horizontal_tile_2_26_to_tile_2_27_1),
		.in_wire_2_2(horizontal_tile_2_26_to_tile_2_27_2),
		.in_wire_2_3(horizontal_tile_2_26_to_tile_2_27_3),
		.out_wire_0_0(horizontal_tile_2_27_to_tile_2_28_0),
		.out_wire_0_1(horizontal_tile_2_27_to_tile_2_28_1),
		.out_wire_0_2(horizontal_tile_2_27_to_tile_2_28_2),
		.out_wire_0_3(horizontal_tile_2_27_to_tile_2_28_3),
		.in_wire_0_0(horizontal_tile_2_28_to_tile_2_27_0),
		.in_wire_0_1(horizontal_tile_2_28_to_tile_2_27_1),
		.in_wire_0_2(horizontal_tile_2_28_to_tile_2_27_2),
		.in_wire_0_3(horizontal_tile_2_28_to_tile_2_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(92)
	);

	pe_tile pe_tile_2_28(
		.out_wire_3_0(vertical_tile_2_28_to_tile_1_28_0),
		.out_wire_3_1(vertical_tile_2_28_to_tile_1_28_1),
		.out_wire_3_2(vertical_tile_2_28_to_tile_1_28_2),
		.out_wire_3_3(vertical_tile_2_28_to_tile_1_28_3),
		.in_wire_3_0(vertical_tile_1_28_to_tile_2_28_0),
		.in_wire_3_1(vertical_tile_1_28_to_tile_2_28_1),
		.in_wire_3_2(vertical_tile_1_28_to_tile_2_28_2),
		.in_wire_3_3(vertical_tile_1_28_to_tile_2_28_3),
		.out_wire_1_0(vertical_tile_2_28_to_tile_3_28_0),
		.out_wire_1_1(vertical_tile_2_28_to_tile_3_28_1),
		.out_wire_1_2(vertical_tile_2_28_to_tile_3_28_2),
		.out_wire_1_3(vertical_tile_2_28_to_tile_3_28_3),
		.in_wire_1_0(vertical_tile_3_28_to_tile_2_28_0),
		.in_wire_1_1(vertical_tile_3_28_to_tile_2_28_1),
		.in_wire_1_2(vertical_tile_3_28_to_tile_2_28_2),
		.in_wire_1_3(vertical_tile_3_28_to_tile_2_28_3),
		.out_wire_2_0(horizontal_tile_2_28_to_tile_2_27_0),
		.out_wire_2_1(horizontal_tile_2_28_to_tile_2_27_1),
		.out_wire_2_2(horizontal_tile_2_28_to_tile_2_27_2),
		.out_wire_2_3(horizontal_tile_2_28_to_tile_2_27_3),
		.in_wire_2_0(horizontal_tile_2_27_to_tile_2_28_0),
		.in_wire_2_1(horizontal_tile_2_27_to_tile_2_28_1),
		.in_wire_2_2(horizontal_tile_2_27_to_tile_2_28_2),
		.in_wire_2_3(horizontal_tile_2_27_to_tile_2_28_3),
		.out_wire_0_0(horizontal_tile_2_28_to_tile_2_29_0),
		.out_wire_0_1(horizontal_tile_2_28_to_tile_2_29_1),
		.out_wire_0_2(horizontal_tile_2_28_to_tile_2_29_2),
		.out_wire_0_3(horizontal_tile_2_28_to_tile_2_29_3),
		.in_wire_0_0(horizontal_tile_2_29_to_tile_2_28_0),
		.in_wire_0_1(horizontal_tile_2_29_to_tile_2_28_1),
		.in_wire_0_2(horizontal_tile_2_29_to_tile_2_28_2),
		.in_wire_0_3(horizontal_tile_2_29_to_tile_2_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(93)
	);

	pe_tile pe_tile_2_29(
		.out_wire_3_0(vertical_tile_2_29_to_tile_1_29_0),
		.out_wire_3_1(vertical_tile_2_29_to_tile_1_29_1),
		.out_wire_3_2(vertical_tile_2_29_to_tile_1_29_2),
		.out_wire_3_3(vertical_tile_2_29_to_tile_1_29_3),
		.in_wire_3_0(vertical_tile_1_29_to_tile_2_29_0),
		.in_wire_3_1(vertical_tile_1_29_to_tile_2_29_1),
		.in_wire_3_2(vertical_tile_1_29_to_tile_2_29_2),
		.in_wire_3_3(vertical_tile_1_29_to_tile_2_29_3),
		.out_wire_1_0(vertical_tile_2_29_to_tile_3_29_0),
		.out_wire_1_1(vertical_tile_2_29_to_tile_3_29_1),
		.out_wire_1_2(vertical_tile_2_29_to_tile_3_29_2),
		.out_wire_1_3(vertical_tile_2_29_to_tile_3_29_3),
		.in_wire_1_0(vertical_tile_3_29_to_tile_2_29_0),
		.in_wire_1_1(vertical_tile_3_29_to_tile_2_29_1),
		.in_wire_1_2(vertical_tile_3_29_to_tile_2_29_2),
		.in_wire_1_3(vertical_tile_3_29_to_tile_2_29_3),
		.out_wire_2_0(horizontal_tile_2_29_to_tile_2_28_0),
		.out_wire_2_1(horizontal_tile_2_29_to_tile_2_28_1),
		.out_wire_2_2(horizontal_tile_2_29_to_tile_2_28_2),
		.out_wire_2_3(horizontal_tile_2_29_to_tile_2_28_3),
		.in_wire_2_0(horizontal_tile_2_28_to_tile_2_29_0),
		.in_wire_2_1(horizontal_tile_2_28_to_tile_2_29_1),
		.in_wire_2_2(horizontal_tile_2_28_to_tile_2_29_2),
		.in_wire_2_3(horizontal_tile_2_28_to_tile_2_29_3),
		.out_wire_0_0(horizontal_tile_2_29_to_tile_2_30_0),
		.out_wire_0_1(horizontal_tile_2_29_to_tile_2_30_1),
		.out_wire_0_2(horizontal_tile_2_29_to_tile_2_30_2),
		.out_wire_0_3(horizontal_tile_2_29_to_tile_2_30_3),
		.in_wire_0_0(horizontal_tile_2_30_to_tile_2_29_0),
		.in_wire_0_1(horizontal_tile_2_30_to_tile_2_29_1),
		.in_wire_0_2(horizontal_tile_2_30_to_tile_2_29_2),
		.in_wire_0_3(horizontal_tile_2_30_to_tile_2_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(94)
	);

	pe_tile pe_tile_2_30(
		.out_wire_3_0(vertical_tile_2_30_to_tile_1_30_0),
		.out_wire_3_1(vertical_tile_2_30_to_tile_1_30_1),
		.out_wire_3_2(vertical_tile_2_30_to_tile_1_30_2),
		.out_wire_3_3(vertical_tile_2_30_to_tile_1_30_3),
		.in_wire_3_0(vertical_tile_1_30_to_tile_2_30_0),
		.in_wire_3_1(vertical_tile_1_30_to_tile_2_30_1),
		.in_wire_3_2(vertical_tile_1_30_to_tile_2_30_2),
		.in_wire_3_3(vertical_tile_1_30_to_tile_2_30_3),
		.out_wire_1_0(vertical_tile_2_30_to_tile_3_30_0),
		.out_wire_1_1(vertical_tile_2_30_to_tile_3_30_1),
		.out_wire_1_2(vertical_tile_2_30_to_tile_3_30_2),
		.out_wire_1_3(vertical_tile_2_30_to_tile_3_30_3),
		.in_wire_1_0(vertical_tile_3_30_to_tile_2_30_0),
		.in_wire_1_1(vertical_tile_3_30_to_tile_2_30_1),
		.in_wire_1_2(vertical_tile_3_30_to_tile_2_30_2),
		.in_wire_1_3(vertical_tile_3_30_to_tile_2_30_3),
		.out_wire_2_0(horizontal_tile_2_30_to_tile_2_29_0),
		.out_wire_2_1(horizontal_tile_2_30_to_tile_2_29_1),
		.out_wire_2_2(horizontal_tile_2_30_to_tile_2_29_2),
		.out_wire_2_3(horizontal_tile_2_30_to_tile_2_29_3),
		.in_wire_2_0(horizontal_tile_2_29_to_tile_2_30_0),
		.in_wire_2_1(horizontal_tile_2_29_to_tile_2_30_1),
		.in_wire_2_2(horizontal_tile_2_29_to_tile_2_30_2),
		.in_wire_2_3(horizontal_tile_2_29_to_tile_2_30_3),
		.out_wire_0_0(horizontal_tile_2_30_to_tile_2_31_0),
		.out_wire_0_1(horizontal_tile_2_30_to_tile_2_31_1),
		.out_wire_0_2(horizontal_tile_2_30_to_tile_2_31_2),
		.out_wire_0_3(horizontal_tile_2_30_to_tile_2_31_3),
		.in_wire_0_0(horizontal_tile_2_31_to_tile_2_30_0),
		.in_wire_0_1(horizontal_tile_2_31_to_tile_2_30_1),
		.in_wire_0_2(horizontal_tile_2_31_to_tile_2_30_2),
		.in_wire_0_3(horizontal_tile_2_31_to_tile_2_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(95)
	);

	pe_tile_right pe_tile_2_31(
		.out_wire_3_0(vertical_tile_2_31_to_tile_1_31_0),
		.out_wire_3_1(vertical_tile_2_31_to_tile_1_31_1),
		.out_wire_3_2(vertical_tile_2_31_to_tile_1_31_2),
		.out_wire_3_3(vertical_tile_2_31_to_tile_1_31_3),
		.in_wire_3_0(vertical_tile_1_31_to_tile_2_31_0),
		.in_wire_3_1(vertical_tile_1_31_to_tile_2_31_1),
		.in_wire_3_2(vertical_tile_1_31_to_tile_2_31_2),
		.in_wire_3_3(vertical_tile_1_31_to_tile_2_31_3),
		.out_wire_1_0(vertical_tile_2_31_to_tile_3_31_0),
		.out_wire_1_1(vertical_tile_2_31_to_tile_3_31_1),
		.out_wire_1_2(vertical_tile_2_31_to_tile_3_31_2),
		.out_wire_1_3(vertical_tile_2_31_to_tile_3_31_3),
		.in_wire_1_0(vertical_tile_3_31_to_tile_2_31_0),
		.in_wire_1_1(vertical_tile_3_31_to_tile_2_31_1),
		.in_wire_1_2(vertical_tile_3_31_to_tile_2_31_2),
		.in_wire_1_3(vertical_tile_3_31_to_tile_2_31_3),
		.out_wire_2_0(horizontal_tile_2_31_to_tile_2_30_0),
		.out_wire_2_1(horizontal_tile_2_31_to_tile_2_30_1),
		.out_wire_2_2(horizontal_tile_2_31_to_tile_2_30_2),
		.out_wire_2_3(horizontal_tile_2_31_to_tile_2_30_3),
		.in_wire_2_0(horizontal_tile_2_30_to_tile_2_31_0),
		.in_wire_2_1(horizontal_tile_2_30_to_tile_2_31_1),
		.in_wire_2_2(horizontal_tile_2_30_to_tile_2_31_2),
		.in_wire_2_3(horizontal_tile_2_30_to_tile_2_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(96)
	);

	pe_tile_left pe_tile_3_0(
		.out_wire_3_0(vertical_tile_3_0_to_tile_2_0_0),
		.out_wire_3_1(vertical_tile_3_0_to_tile_2_0_1),
		.out_wire_3_2(vertical_tile_3_0_to_tile_2_0_2),
		.out_wire_3_3(vertical_tile_3_0_to_tile_2_0_3),
		.in_wire_3_0(vertical_tile_2_0_to_tile_3_0_0),
		.in_wire_3_1(vertical_tile_2_0_to_tile_3_0_1),
		.in_wire_3_2(vertical_tile_2_0_to_tile_3_0_2),
		.in_wire_3_3(vertical_tile_2_0_to_tile_3_0_3),
		.out_wire_1_0(vertical_tile_3_0_to_tile_4_0_0),
		.out_wire_1_1(vertical_tile_3_0_to_tile_4_0_1),
		.out_wire_1_2(vertical_tile_3_0_to_tile_4_0_2),
		.out_wire_1_3(vertical_tile_3_0_to_tile_4_0_3),
		.in_wire_1_0(vertical_tile_4_0_to_tile_3_0_0),
		.in_wire_1_1(vertical_tile_4_0_to_tile_3_0_1),
		.in_wire_1_2(vertical_tile_4_0_to_tile_3_0_2),
		.in_wire_1_3(vertical_tile_4_0_to_tile_3_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_3_0_to_tile_3_1_0),
		.out_wire_0_1(horizontal_tile_3_0_to_tile_3_1_1),
		.out_wire_0_2(horizontal_tile_3_0_to_tile_3_1_2),
		.out_wire_0_3(horizontal_tile_3_0_to_tile_3_1_3),
		.in_wire_0_0(horizontal_tile_3_1_to_tile_3_0_0),
		.in_wire_0_1(horizontal_tile_3_1_to_tile_3_0_1),
		.in_wire_0_2(horizontal_tile_3_1_to_tile_3_0_2),
		.in_wire_0_3(horizontal_tile_3_1_to_tile_3_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(97)
	);

	pe_tile pe_tile_3_1(
		.out_wire_3_0(vertical_tile_3_1_to_tile_2_1_0),
		.out_wire_3_1(vertical_tile_3_1_to_tile_2_1_1),
		.out_wire_3_2(vertical_tile_3_1_to_tile_2_1_2),
		.out_wire_3_3(vertical_tile_3_1_to_tile_2_1_3),
		.in_wire_3_0(vertical_tile_2_1_to_tile_3_1_0),
		.in_wire_3_1(vertical_tile_2_1_to_tile_3_1_1),
		.in_wire_3_2(vertical_tile_2_1_to_tile_3_1_2),
		.in_wire_3_3(vertical_tile_2_1_to_tile_3_1_3),
		.out_wire_1_0(vertical_tile_3_1_to_tile_4_1_0),
		.out_wire_1_1(vertical_tile_3_1_to_tile_4_1_1),
		.out_wire_1_2(vertical_tile_3_1_to_tile_4_1_2),
		.out_wire_1_3(vertical_tile_3_1_to_tile_4_1_3),
		.in_wire_1_0(vertical_tile_4_1_to_tile_3_1_0),
		.in_wire_1_1(vertical_tile_4_1_to_tile_3_1_1),
		.in_wire_1_2(vertical_tile_4_1_to_tile_3_1_2),
		.in_wire_1_3(vertical_tile_4_1_to_tile_3_1_3),
		.out_wire_2_0(horizontal_tile_3_1_to_tile_3_0_0),
		.out_wire_2_1(horizontal_tile_3_1_to_tile_3_0_1),
		.out_wire_2_2(horizontal_tile_3_1_to_tile_3_0_2),
		.out_wire_2_3(horizontal_tile_3_1_to_tile_3_0_3),
		.in_wire_2_0(horizontal_tile_3_0_to_tile_3_1_0),
		.in_wire_2_1(horizontal_tile_3_0_to_tile_3_1_1),
		.in_wire_2_2(horizontal_tile_3_0_to_tile_3_1_2),
		.in_wire_2_3(horizontal_tile_3_0_to_tile_3_1_3),
		.out_wire_0_0(horizontal_tile_3_1_to_tile_3_2_0),
		.out_wire_0_1(horizontal_tile_3_1_to_tile_3_2_1),
		.out_wire_0_2(horizontal_tile_3_1_to_tile_3_2_2),
		.out_wire_0_3(horizontal_tile_3_1_to_tile_3_2_3),
		.in_wire_0_0(horizontal_tile_3_2_to_tile_3_1_0),
		.in_wire_0_1(horizontal_tile_3_2_to_tile_3_1_1),
		.in_wire_0_2(horizontal_tile_3_2_to_tile_3_1_2),
		.in_wire_0_3(horizontal_tile_3_2_to_tile_3_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(98)
	);

	pe_tile pe_tile_3_2(
		.out_wire_3_0(vertical_tile_3_2_to_tile_2_2_0),
		.out_wire_3_1(vertical_tile_3_2_to_tile_2_2_1),
		.out_wire_3_2(vertical_tile_3_2_to_tile_2_2_2),
		.out_wire_3_3(vertical_tile_3_2_to_tile_2_2_3),
		.in_wire_3_0(vertical_tile_2_2_to_tile_3_2_0),
		.in_wire_3_1(vertical_tile_2_2_to_tile_3_2_1),
		.in_wire_3_2(vertical_tile_2_2_to_tile_3_2_2),
		.in_wire_3_3(vertical_tile_2_2_to_tile_3_2_3),
		.out_wire_1_0(vertical_tile_3_2_to_tile_4_2_0),
		.out_wire_1_1(vertical_tile_3_2_to_tile_4_2_1),
		.out_wire_1_2(vertical_tile_3_2_to_tile_4_2_2),
		.out_wire_1_3(vertical_tile_3_2_to_tile_4_2_3),
		.in_wire_1_0(vertical_tile_4_2_to_tile_3_2_0),
		.in_wire_1_1(vertical_tile_4_2_to_tile_3_2_1),
		.in_wire_1_2(vertical_tile_4_2_to_tile_3_2_2),
		.in_wire_1_3(vertical_tile_4_2_to_tile_3_2_3),
		.out_wire_2_0(horizontal_tile_3_2_to_tile_3_1_0),
		.out_wire_2_1(horizontal_tile_3_2_to_tile_3_1_1),
		.out_wire_2_2(horizontal_tile_3_2_to_tile_3_1_2),
		.out_wire_2_3(horizontal_tile_3_2_to_tile_3_1_3),
		.in_wire_2_0(horizontal_tile_3_1_to_tile_3_2_0),
		.in_wire_2_1(horizontal_tile_3_1_to_tile_3_2_1),
		.in_wire_2_2(horizontal_tile_3_1_to_tile_3_2_2),
		.in_wire_2_3(horizontal_tile_3_1_to_tile_3_2_3),
		.out_wire_0_0(horizontal_tile_3_2_to_tile_3_3_0),
		.out_wire_0_1(horizontal_tile_3_2_to_tile_3_3_1),
		.out_wire_0_2(horizontal_tile_3_2_to_tile_3_3_2),
		.out_wire_0_3(horizontal_tile_3_2_to_tile_3_3_3),
		.in_wire_0_0(horizontal_tile_3_3_to_tile_3_2_0),
		.in_wire_0_1(horizontal_tile_3_3_to_tile_3_2_1),
		.in_wire_0_2(horizontal_tile_3_3_to_tile_3_2_2),
		.in_wire_0_3(horizontal_tile_3_3_to_tile_3_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(99)
	);

	pe_tile pe_tile_3_3(
		.out_wire_3_0(vertical_tile_3_3_to_tile_2_3_0),
		.out_wire_3_1(vertical_tile_3_3_to_tile_2_3_1),
		.out_wire_3_2(vertical_tile_3_3_to_tile_2_3_2),
		.out_wire_3_3(vertical_tile_3_3_to_tile_2_3_3),
		.in_wire_3_0(vertical_tile_2_3_to_tile_3_3_0),
		.in_wire_3_1(vertical_tile_2_3_to_tile_3_3_1),
		.in_wire_3_2(vertical_tile_2_3_to_tile_3_3_2),
		.in_wire_3_3(vertical_tile_2_3_to_tile_3_3_3),
		.out_wire_1_0(vertical_tile_3_3_to_tile_4_3_0),
		.out_wire_1_1(vertical_tile_3_3_to_tile_4_3_1),
		.out_wire_1_2(vertical_tile_3_3_to_tile_4_3_2),
		.out_wire_1_3(vertical_tile_3_3_to_tile_4_3_3),
		.in_wire_1_0(vertical_tile_4_3_to_tile_3_3_0),
		.in_wire_1_1(vertical_tile_4_3_to_tile_3_3_1),
		.in_wire_1_2(vertical_tile_4_3_to_tile_3_3_2),
		.in_wire_1_3(vertical_tile_4_3_to_tile_3_3_3),
		.out_wire_2_0(horizontal_tile_3_3_to_tile_3_2_0),
		.out_wire_2_1(horizontal_tile_3_3_to_tile_3_2_1),
		.out_wire_2_2(horizontal_tile_3_3_to_tile_3_2_2),
		.out_wire_2_3(horizontal_tile_3_3_to_tile_3_2_3),
		.in_wire_2_0(horizontal_tile_3_2_to_tile_3_3_0),
		.in_wire_2_1(horizontal_tile_3_2_to_tile_3_3_1),
		.in_wire_2_2(horizontal_tile_3_2_to_tile_3_3_2),
		.in_wire_2_3(horizontal_tile_3_2_to_tile_3_3_3),
		.out_wire_0_0(horizontal_tile_3_3_to_tile_3_4_0),
		.out_wire_0_1(horizontal_tile_3_3_to_tile_3_4_1),
		.out_wire_0_2(horizontal_tile_3_3_to_tile_3_4_2),
		.out_wire_0_3(horizontal_tile_3_3_to_tile_3_4_3),
		.in_wire_0_0(horizontal_tile_3_4_to_tile_3_3_0),
		.in_wire_0_1(horizontal_tile_3_4_to_tile_3_3_1),
		.in_wire_0_2(horizontal_tile_3_4_to_tile_3_3_2),
		.in_wire_0_3(horizontal_tile_3_4_to_tile_3_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(100)
	);

	pe_tile pe_tile_3_4(
		.out_wire_3_0(vertical_tile_3_4_to_tile_2_4_0),
		.out_wire_3_1(vertical_tile_3_4_to_tile_2_4_1),
		.out_wire_3_2(vertical_tile_3_4_to_tile_2_4_2),
		.out_wire_3_3(vertical_tile_3_4_to_tile_2_4_3),
		.in_wire_3_0(vertical_tile_2_4_to_tile_3_4_0),
		.in_wire_3_1(vertical_tile_2_4_to_tile_3_4_1),
		.in_wire_3_2(vertical_tile_2_4_to_tile_3_4_2),
		.in_wire_3_3(vertical_tile_2_4_to_tile_3_4_3),
		.out_wire_1_0(vertical_tile_3_4_to_tile_4_4_0),
		.out_wire_1_1(vertical_tile_3_4_to_tile_4_4_1),
		.out_wire_1_2(vertical_tile_3_4_to_tile_4_4_2),
		.out_wire_1_3(vertical_tile_3_4_to_tile_4_4_3),
		.in_wire_1_0(vertical_tile_4_4_to_tile_3_4_0),
		.in_wire_1_1(vertical_tile_4_4_to_tile_3_4_1),
		.in_wire_1_2(vertical_tile_4_4_to_tile_3_4_2),
		.in_wire_1_3(vertical_tile_4_4_to_tile_3_4_3),
		.out_wire_2_0(horizontal_tile_3_4_to_tile_3_3_0),
		.out_wire_2_1(horizontal_tile_3_4_to_tile_3_3_1),
		.out_wire_2_2(horizontal_tile_3_4_to_tile_3_3_2),
		.out_wire_2_3(horizontal_tile_3_4_to_tile_3_3_3),
		.in_wire_2_0(horizontal_tile_3_3_to_tile_3_4_0),
		.in_wire_2_1(horizontal_tile_3_3_to_tile_3_4_1),
		.in_wire_2_2(horizontal_tile_3_3_to_tile_3_4_2),
		.in_wire_2_3(horizontal_tile_3_3_to_tile_3_4_3),
		.out_wire_0_0(horizontal_tile_3_4_to_tile_3_5_0),
		.out_wire_0_1(horizontal_tile_3_4_to_tile_3_5_1),
		.out_wire_0_2(horizontal_tile_3_4_to_tile_3_5_2),
		.out_wire_0_3(horizontal_tile_3_4_to_tile_3_5_3),
		.in_wire_0_0(horizontal_tile_3_5_to_tile_3_4_0),
		.in_wire_0_1(horizontal_tile_3_5_to_tile_3_4_1),
		.in_wire_0_2(horizontal_tile_3_5_to_tile_3_4_2),
		.in_wire_0_3(horizontal_tile_3_5_to_tile_3_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(101)
	);

	pe_tile pe_tile_3_5(
		.out_wire_3_0(vertical_tile_3_5_to_tile_2_5_0),
		.out_wire_3_1(vertical_tile_3_5_to_tile_2_5_1),
		.out_wire_3_2(vertical_tile_3_5_to_tile_2_5_2),
		.out_wire_3_3(vertical_tile_3_5_to_tile_2_5_3),
		.in_wire_3_0(vertical_tile_2_5_to_tile_3_5_0),
		.in_wire_3_1(vertical_tile_2_5_to_tile_3_5_1),
		.in_wire_3_2(vertical_tile_2_5_to_tile_3_5_2),
		.in_wire_3_3(vertical_tile_2_5_to_tile_3_5_3),
		.out_wire_1_0(vertical_tile_3_5_to_tile_4_5_0),
		.out_wire_1_1(vertical_tile_3_5_to_tile_4_5_1),
		.out_wire_1_2(vertical_tile_3_5_to_tile_4_5_2),
		.out_wire_1_3(vertical_tile_3_5_to_tile_4_5_3),
		.in_wire_1_0(vertical_tile_4_5_to_tile_3_5_0),
		.in_wire_1_1(vertical_tile_4_5_to_tile_3_5_1),
		.in_wire_1_2(vertical_tile_4_5_to_tile_3_5_2),
		.in_wire_1_3(vertical_tile_4_5_to_tile_3_5_3),
		.out_wire_2_0(horizontal_tile_3_5_to_tile_3_4_0),
		.out_wire_2_1(horizontal_tile_3_5_to_tile_3_4_1),
		.out_wire_2_2(horizontal_tile_3_5_to_tile_3_4_2),
		.out_wire_2_3(horizontal_tile_3_5_to_tile_3_4_3),
		.in_wire_2_0(horizontal_tile_3_4_to_tile_3_5_0),
		.in_wire_2_1(horizontal_tile_3_4_to_tile_3_5_1),
		.in_wire_2_2(horizontal_tile_3_4_to_tile_3_5_2),
		.in_wire_2_3(horizontal_tile_3_4_to_tile_3_5_3),
		.out_wire_0_0(horizontal_tile_3_5_to_tile_3_6_0),
		.out_wire_0_1(horizontal_tile_3_5_to_tile_3_6_1),
		.out_wire_0_2(horizontal_tile_3_5_to_tile_3_6_2),
		.out_wire_0_3(horizontal_tile_3_5_to_tile_3_6_3),
		.in_wire_0_0(horizontal_tile_3_6_to_tile_3_5_0),
		.in_wire_0_1(horizontal_tile_3_6_to_tile_3_5_1),
		.in_wire_0_2(horizontal_tile_3_6_to_tile_3_5_2),
		.in_wire_0_3(horizontal_tile_3_6_to_tile_3_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(102)
	);

	pe_tile pe_tile_3_6(
		.out_wire_3_0(vertical_tile_3_6_to_tile_2_6_0),
		.out_wire_3_1(vertical_tile_3_6_to_tile_2_6_1),
		.out_wire_3_2(vertical_tile_3_6_to_tile_2_6_2),
		.out_wire_3_3(vertical_tile_3_6_to_tile_2_6_3),
		.in_wire_3_0(vertical_tile_2_6_to_tile_3_6_0),
		.in_wire_3_1(vertical_tile_2_6_to_tile_3_6_1),
		.in_wire_3_2(vertical_tile_2_6_to_tile_3_6_2),
		.in_wire_3_3(vertical_tile_2_6_to_tile_3_6_3),
		.out_wire_1_0(vertical_tile_3_6_to_tile_4_6_0),
		.out_wire_1_1(vertical_tile_3_6_to_tile_4_6_1),
		.out_wire_1_2(vertical_tile_3_6_to_tile_4_6_2),
		.out_wire_1_3(vertical_tile_3_6_to_tile_4_6_3),
		.in_wire_1_0(vertical_tile_4_6_to_tile_3_6_0),
		.in_wire_1_1(vertical_tile_4_6_to_tile_3_6_1),
		.in_wire_1_2(vertical_tile_4_6_to_tile_3_6_2),
		.in_wire_1_3(vertical_tile_4_6_to_tile_3_6_3),
		.out_wire_2_0(horizontal_tile_3_6_to_tile_3_5_0),
		.out_wire_2_1(horizontal_tile_3_6_to_tile_3_5_1),
		.out_wire_2_2(horizontal_tile_3_6_to_tile_3_5_2),
		.out_wire_2_3(horizontal_tile_3_6_to_tile_3_5_3),
		.in_wire_2_0(horizontal_tile_3_5_to_tile_3_6_0),
		.in_wire_2_1(horizontal_tile_3_5_to_tile_3_6_1),
		.in_wire_2_2(horizontal_tile_3_5_to_tile_3_6_2),
		.in_wire_2_3(horizontal_tile_3_5_to_tile_3_6_3),
		.out_wire_0_0(horizontal_tile_3_6_to_tile_3_7_0),
		.out_wire_0_1(horizontal_tile_3_6_to_tile_3_7_1),
		.out_wire_0_2(horizontal_tile_3_6_to_tile_3_7_2),
		.out_wire_0_3(horizontal_tile_3_6_to_tile_3_7_3),
		.in_wire_0_0(horizontal_tile_3_7_to_tile_3_6_0),
		.in_wire_0_1(horizontal_tile_3_7_to_tile_3_6_1),
		.in_wire_0_2(horizontal_tile_3_7_to_tile_3_6_2),
		.in_wire_0_3(horizontal_tile_3_7_to_tile_3_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(103)
	);

	pe_tile pe_tile_3_7(
		.out_wire_3_0(vertical_tile_3_7_to_tile_2_7_0),
		.out_wire_3_1(vertical_tile_3_7_to_tile_2_7_1),
		.out_wire_3_2(vertical_tile_3_7_to_tile_2_7_2),
		.out_wire_3_3(vertical_tile_3_7_to_tile_2_7_3),
		.in_wire_3_0(vertical_tile_2_7_to_tile_3_7_0),
		.in_wire_3_1(vertical_tile_2_7_to_tile_3_7_1),
		.in_wire_3_2(vertical_tile_2_7_to_tile_3_7_2),
		.in_wire_3_3(vertical_tile_2_7_to_tile_3_7_3),
		.out_wire_1_0(vertical_tile_3_7_to_tile_4_7_0),
		.out_wire_1_1(vertical_tile_3_7_to_tile_4_7_1),
		.out_wire_1_2(vertical_tile_3_7_to_tile_4_7_2),
		.out_wire_1_3(vertical_tile_3_7_to_tile_4_7_3),
		.in_wire_1_0(vertical_tile_4_7_to_tile_3_7_0),
		.in_wire_1_1(vertical_tile_4_7_to_tile_3_7_1),
		.in_wire_1_2(vertical_tile_4_7_to_tile_3_7_2),
		.in_wire_1_3(vertical_tile_4_7_to_tile_3_7_3),
		.out_wire_2_0(horizontal_tile_3_7_to_tile_3_6_0),
		.out_wire_2_1(horizontal_tile_3_7_to_tile_3_6_1),
		.out_wire_2_2(horizontal_tile_3_7_to_tile_3_6_2),
		.out_wire_2_3(horizontal_tile_3_7_to_tile_3_6_3),
		.in_wire_2_0(horizontal_tile_3_6_to_tile_3_7_0),
		.in_wire_2_1(horizontal_tile_3_6_to_tile_3_7_1),
		.in_wire_2_2(horizontal_tile_3_6_to_tile_3_7_2),
		.in_wire_2_3(horizontal_tile_3_6_to_tile_3_7_3),
		.out_wire_0_0(horizontal_tile_3_7_to_tile_3_8_0),
		.out_wire_0_1(horizontal_tile_3_7_to_tile_3_8_1),
		.out_wire_0_2(horizontal_tile_3_7_to_tile_3_8_2),
		.out_wire_0_3(horizontal_tile_3_7_to_tile_3_8_3),
		.in_wire_0_0(horizontal_tile_3_8_to_tile_3_7_0),
		.in_wire_0_1(horizontal_tile_3_8_to_tile_3_7_1),
		.in_wire_0_2(horizontal_tile_3_8_to_tile_3_7_2),
		.in_wire_0_3(horizontal_tile_3_8_to_tile_3_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(104)
	);

	pe_tile pe_tile_3_8(
		.out_wire_3_0(vertical_tile_3_8_to_tile_2_8_0),
		.out_wire_3_1(vertical_tile_3_8_to_tile_2_8_1),
		.out_wire_3_2(vertical_tile_3_8_to_tile_2_8_2),
		.out_wire_3_3(vertical_tile_3_8_to_tile_2_8_3),
		.in_wire_3_0(vertical_tile_2_8_to_tile_3_8_0),
		.in_wire_3_1(vertical_tile_2_8_to_tile_3_8_1),
		.in_wire_3_2(vertical_tile_2_8_to_tile_3_8_2),
		.in_wire_3_3(vertical_tile_2_8_to_tile_3_8_3),
		.out_wire_1_0(vertical_tile_3_8_to_tile_4_8_0),
		.out_wire_1_1(vertical_tile_3_8_to_tile_4_8_1),
		.out_wire_1_2(vertical_tile_3_8_to_tile_4_8_2),
		.out_wire_1_3(vertical_tile_3_8_to_tile_4_8_3),
		.in_wire_1_0(vertical_tile_4_8_to_tile_3_8_0),
		.in_wire_1_1(vertical_tile_4_8_to_tile_3_8_1),
		.in_wire_1_2(vertical_tile_4_8_to_tile_3_8_2),
		.in_wire_1_3(vertical_tile_4_8_to_tile_3_8_3),
		.out_wire_2_0(horizontal_tile_3_8_to_tile_3_7_0),
		.out_wire_2_1(horizontal_tile_3_8_to_tile_3_7_1),
		.out_wire_2_2(horizontal_tile_3_8_to_tile_3_7_2),
		.out_wire_2_3(horizontal_tile_3_8_to_tile_3_7_3),
		.in_wire_2_0(horizontal_tile_3_7_to_tile_3_8_0),
		.in_wire_2_1(horizontal_tile_3_7_to_tile_3_8_1),
		.in_wire_2_2(horizontal_tile_3_7_to_tile_3_8_2),
		.in_wire_2_3(horizontal_tile_3_7_to_tile_3_8_3),
		.out_wire_0_0(horizontal_tile_3_8_to_tile_3_9_0),
		.out_wire_0_1(horizontal_tile_3_8_to_tile_3_9_1),
		.out_wire_0_2(horizontal_tile_3_8_to_tile_3_9_2),
		.out_wire_0_3(horizontal_tile_3_8_to_tile_3_9_3),
		.in_wire_0_0(horizontal_tile_3_9_to_tile_3_8_0),
		.in_wire_0_1(horizontal_tile_3_9_to_tile_3_8_1),
		.in_wire_0_2(horizontal_tile_3_9_to_tile_3_8_2),
		.in_wire_0_3(horizontal_tile_3_9_to_tile_3_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(105)
	);

	pe_tile pe_tile_3_9(
		.out_wire_3_0(vertical_tile_3_9_to_tile_2_9_0),
		.out_wire_3_1(vertical_tile_3_9_to_tile_2_9_1),
		.out_wire_3_2(vertical_tile_3_9_to_tile_2_9_2),
		.out_wire_3_3(vertical_tile_3_9_to_tile_2_9_3),
		.in_wire_3_0(vertical_tile_2_9_to_tile_3_9_0),
		.in_wire_3_1(vertical_tile_2_9_to_tile_3_9_1),
		.in_wire_3_2(vertical_tile_2_9_to_tile_3_9_2),
		.in_wire_3_3(vertical_tile_2_9_to_tile_3_9_3),
		.out_wire_1_0(vertical_tile_3_9_to_tile_4_9_0),
		.out_wire_1_1(vertical_tile_3_9_to_tile_4_9_1),
		.out_wire_1_2(vertical_tile_3_9_to_tile_4_9_2),
		.out_wire_1_3(vertical_tile_3_9_to_tile_4_9_3),
		.in_wire_1_0(vertical_tile_4_9_to_tile_3_9_0),
		.in_wire_1_1(vertical_tile_4_9_to_tile_3_9_1),
		.in_wire_1_2(vertical_tile_4_9_to_tile_3_9_2),
		.in_wire_1_3(vertical_tile_4_9_to_tile_3_9_3),
		.out_wire_2_0(horizontal_tile_3_9_to_tile_3_8_0),
		.out_wire_2_1(horizontal_tile_3_9_to_tile_3_8_1),
		.out_wire_2_2(horizontal_tile_3_9_to_tile_3_8_2),
		.out_wire_2_3(horizontal_tile_3_9_to_tile_3_8_3),
		.in_wire_2_0(horizontal_tile_3_8_to_tile_3_9_0),
		.in_wire_2_1(horizontal_tile_3_8_to_tile_3_9_1),
		.in_wire_2_2(horizontal_tile_3_8_to_tile_3_9_2),
		.in_wire_2_3(horizontal_tile_3_8_to_tile_3_9_3),
		.out_wire_0_0(horizontal_tile_3_9_to_tile_3_10_0),
		.out_wire_0_1(horizontal_tile_3_9_to_tile_3_10_1),
		.out_wire_0_2(horizontal_tile_3_9_to_tile_3_10_2),
		.out_wire_0_3(horizontal_tile_3_9_to_tile_3_10_3),
		.in_wire_0_0(horizontal_tile_3_10_to_tile_3_9_0),
		.in_wire_0_1(horizontal_tile_3_10_to_tile_3_9_1),
		.in_wire_0_2(horizontal_tile_3_10_to_tile_3_9_2),
		.in_wire_0_3(horizontal_tile_3_10_to_tile_3_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(106)
	);

	pe_tile pe_tile_3_10(
		.out_wire_3_0(vertical_tile_3_10_to_tile_2_10_0),
		.out_wire_3_1(vertical_tile_3_10_to_tile_2_10_1),
		.out_wire_3_2(vertical_tile_3_10_to_tile_2_10_2),
		.out_wire_3_3(vertical_tile_3_10_to_tile_2_10_3),
		.in_wire_3_0(vertical_tile_2_10_to_tile_3_10_0),
		.in_wire_3_1(vertical_tile_2_10_to_tile_3_10_1),
		.in_wire_3_2(vertical_tile_2_10_to_tile_3_10_2),
		.in_wire_3_3(vertical_tile_2_10_to_tile_3_10_3),
		.out_wire_1_0(vertical_tile_3_10_to_tile_4_10_0),
		.out_wire_1_1(vertical_tile_3_10_to_tile_4_10_1),
		.out_wire_1_2(vertical_tile_3_10_to_tile_4_10_2),
		.out_wire_1_3(vertical_tile_3_10_to_tile_4_10_3),
		.in_wire_1_0(vertical_tile_4_10_to_tile_3_10_0),
		.in_wire_1_1(vertical_tile_4_10_to_tile_3_10_1),
		.in_wire_1_2(vertical_tile_4_10_to_tile_3_10_2),
		.in_wire_1_3(vertical_tile_4_10_to_tile_3_10_3),
		.out_wire_2_0(horizontal_tile_3_10_to_tile_3_9_0),
		.out_wire_2_1(horizontal_tile_3_10_to_tile_3_9_1),
		.out_wire_2_2(horizontal_tile_3_10_to_tile_3_9_2),
		.out_wire_2_3(horizontal_tile_3_10_to_tile_3_9_3),
		.in_wire_2_0(horizontal_tile_3_9_to_tile_3_10_0),
		.in_wire_2_1(horizontal_tile_3_9_to_tile_3_10_1),
		.in_wire_2_2(horizontal_tile_3_9_to_tile_3_10_2),
		.in_wire_2_3(horizontal_tile_3_9_to_tile_3_10_3),
		.out_wire_0_0(horizontal_tile_3_10_to_tile_3_11_0),
		.out_wire_0_1(horizontal_tile_3_10_to_tile_3_11_1),
		.out_wire_0_2(horizontal_tile_3_10_to_tile_3_11_2),
		.out_wire_0_3(horizontal_tile_3_10_to_tile_3_11_3),
		.in_wire_0_0(horizontal_tile_3_11_to_tile_3_10_0),
		.in_wire_0_1(horizontal_tile_3_11_to_tile_3_10_1),
		.in_wire_0_2(horizontal_tile_3_11_to_tile_3_10_2),
		.in_wire_0_3(horizontal_tile_3_11_to_tile_3_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(107)
	);

	pe_tile pe_tile_3_11(
		.out_wire_3_0(vertical_tile_3_11_to_tile_2_11_0),
		.out_wire_3_1(vertical_tile_3_11_to_tile_2_11_1),
		.out_wire_3_2(vertical_tile_3_11_to_tile_2_11_2),
		.out_wire_3_3(vertical_tile_3_11_to_tile_2_11_3),
		.in_wire_3_0(vertical_tile_2_11_to_tile_3_11_0),
		.in_wire_3_1(vertical_tile_2_11_to_tile_3_11_1),
		.in_wire_3_2(vertical_tile_2_11_to_tile_3_11_2),
		.in_wire_3_3(vertical_tile_2_11_to_tile_3_11_3),
		.out_wire_1_0(vertical_tile_3_11_to_tile_4_11_0),
		.out_wire_1_1(vertical_tile_3_11_to_tile_4_11_1),
		.out_wire_1_2(vertical_tile_3_11_to_tile_4_11_2),
		.out_wire_1_3(vertical_tile_3_11_to_tile_4_11_3),
		.in_wire_1_0(vertical_tile_4_11_to_tile_3_11_0),
		.in_wire_1_1(vertical_tile_4_11_to_tile_3_11_1),
		.in_wire_1_2(vertical_tile_4_11_to_tile_3_11_2),
		.in_wire_1_3(vertical_tile_4_11_to_tile_3_11_3),
		.out_wire_2_0(horizontal_tile_3_11_to_tile_3_10_0),
		.out_wire_2_1(horizontal_tile_3_11_to_tile_3_10_1),
		.out_wire_2_2(horizontal_tile_3_11_to_tile_3_10_2),
		.out_wire_2_3(horizontal_tile_3_11_to_tile_3_10_3),
		.in_wire_2_0(horizontal_tile_3_10_to_tile_3_11_0),
		.in_wire_2_1(horizontal_tile_3_10_to_tile_3_11_1),
		.in_wire_2_2(horizontal_tile_3_10_to_tile_3_11_2),
		.in_wire_2_3(horizontal_tile_3_10_to_tile_3_11_3),
		.out_wire_0_0(horizontal_tile_3_11_to_tile_3_12_0),
		.out_wire_0_1(horizontal_tile_3_11_to_tile_3_12_1),
		.out_wire_0_2(horizontal_tile_3_11_to_tile_3_12_2),
		.out_wire_0_3(horizontal_tile_3_11_to_tile_3_12_3),
		.in_wire_0_0(horizontal_tile_3_12_to_tile_3_11_0),
		.in_wire_0_1(horizontal_tile_3_12_to_tile_3_11_1),
		.in_wire_0_2(horizontal_tile_3_12_to_tile_3_11_2),
		.in_wire_0_3(horizontal_tile_3_12_to_tile_3_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(108)
	);

	pe_tile pe_tile_3_12(
		.out_wire_3_0(vertical_tile_3_12_to_tile_2_12_0),
		.out_wire_3_1(vertical_tile_3_12_to_tile_2_12_1),
		.out_wire_3_2(vertical_tile_3_12_to_tile_2_12_2),
		.out_wire_3_3(vertical_tile_3_12_to_tile_2_12_3),
		.in_wire_3_0(vertical_tile_2_12_to_tile_3_12_0),
		.in_wire_3_1(vertical_tile_2_12_to_tile_3_12_1),
		.in_wire_3_2(vertical_tile_2_12_to_tile_3_12_2),
		.in_wire_3_3(vertical_tile_2_12_to_tile_3_12_3),
		.out_wire_1_0(vertical_tile_3_12_to_tile_4_12_0),
		.out_wire_1_1(vertical_tile_3_12_to_tile_4_12_1),
		.out_wire_1_2(vertical_tile_3_12_to_tile_4_12_2),
		.out_wire_1_3(vertical_tile_3_12_to_tile_4_12_3),
		.in_wire_1_0(vertical_tile_4_12_to_tile_3_12_0),
		.in_wire_1_1(vertical_tile_4_12_to_tile_3_12_1),
		.in_wire_1_2(vertical_tile_4_12_to_tile_3_12_2),
		.in_wire_1_3(vertical_tile_4_12_to_tile_3_12_3),
		.out_wire_2_0(horizontal_tile_3_12_to_tile_3_11_0),
		.out_wire_2_1(horizontal_tile_3_12_to_tile_3_11_1),
		.out_wire_2_2(horizontal_tile_3_12_to_tile_3_11_2),
		.out_wire_2_3(horizontal_tile_3_12_to_tile_3_11_3),
		.in_wire_2_0(horizontal_tile_3_11_to_tile_3_12_0),
		.in_wire_2_1(horizontal_tile_3_11_to_tile_3_12_1),
		.in_wire_2_2(horizontal_tile_3_11_to_tile_3_12_2),
		.in_wire_2_3(horizontal_tile_3_11_to_tile_3_12_3),
		.out_wire_0_0(horizontal_tile_3_12_to_tile_3_13_0),
		.out_wire_0_1(horizontal_tile_3_12_to_tile_3_13_1),
		.out_wire_0_2(horizontal_tile_3_12_to_tile_3_13_2),
		.out_wire_0_3(horizontal_tile_3_12_to_tile_3_13_3),
		.in_wire_0_0(horizontal_tile_3_13_to_tile_3_12_0),
		.in_wire_0_1(horizontal_tile_3_13_to_tile_3_12_1),
		.in_wire_0_2(horizontal_tile_3_13_to_tile_3_12_2),
		.in_wire_0_3(horizontal_tile_3_13_to_tile_3_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(109)
	);

	pe_tile pe_tile_3_13(
		.out_wire_3_0(vertical_tile_3_13_to_tile_2_13_0),
		.out_wire_3_1(vertical_tile_3_13_to_tile_2_13_1),
		.out_wire_3_2(vertical_tile_3_13_to_tile_2_13_2),
		.out_wire_3_3(vertical_tile_3_13_to_tile_2_13_3),
		.in_wire_3_0(vertical_tile_2_13_to_tile_3_13_0),
		.in_wire_3_1(vertical_tile_2_13_to_tile_3_13_1),
		.in_wire_3_2(vertical_tile_2_13_to_tile_3_13_2),
		.in_wire_3_3(vertical_tile_2_13_to_tile_3_13_3),
		.out_wire_1_0(vertical_tile_3_13_to_tile_4_13_0),
		.out_wire_1_1(vertical_tile_3_13_to_tile_4_13_1),
		.out_wire_1_2(vertical_tile_3_13_to_tile_4_13_2),
		.out_wire_1_3(vertical_tile_3_13_to_tile_4_13_3),
		.in_wire_1_0(vertical_tile_4_13_to_tile_3_13_0),
		.in_wire_1_1(vertical_tile_4_13_to_tile_3_13_1),
		.in_wire_1_2(vertical_tile_4_13_to_tile_3_13_2),
		.in_wire_1_3(vertical_tile_4_13_to_tile_3_13_3),
		.out_wire_2_0(horizontal_tile_3_13_to_tile_3_12_0),
		.out_wire_2_1(horizontal_tile_3_13_to_tile_3_12_1),
		.out_wire_2_2(horizontal_tile_3_13_to_tile_3_12_2),
		.out_wire_2_3(horizontal_tile_3_13_to_tile_3_12_3),
		.in_wire_2_0(horizontal_tile_3_12_to_tile_3_13_0),
		.in_wire_2_1(horizontal_tile_3_12_to_tile_3_13_1),
		.in_wire_2_2(horizontal_tile_3_12_to_tile_3_13_2),
		.in_wire_2_3(horizontal_tile_3_12_to_tile_3_13_3),
		.out_wire_0_0(horizontal_tile_3_13_to_tile_3_14_0),
		.out_wire_0_1(horizontal_tile_3_13_to_tile_3_14_1),
		.out_wire_0_2(horizontal_tile_3_13_to_tile_3_14_2),
		.out_wire_0_3(horizontal_tile_3_13_to_tile_3_14_3),
		.in_wire_0_0(horizontal_tile_3_14_to_tile_3_13_0),
		.in_wire_0_1(horizontal_tile_3_14_to_tile_3_13_1),
		.in_wire_0_2(horizontal_tile_3_14_to_tile_3_13_2),
		.in_wire_0_3(horizontal_tile_3_14_to_tile_3_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(110)
	);

	pe_tile pe_tile_3_14(
		.out_wire_3_0(vertical_tile_3_14_to_tile_2_14_0),
		.out_wire_3_1(vertical_tile_3_14_to_tile_2_14_1),
		.out_wire_3_2(vertical_tile_3_14_to_tile_2_14_2),
		.out_wire_3_3(vertical_tile_3_14_to_tile_2_14_3),
		.in_wire_3_0(vertical_tile_2_14_to_tile_3_14_0),
		.in_wire_3_1(vertical_tile_2_14_to_tile_3_14_1),
		.in_wire_3_2(vertical_tile_2_14_to_tile_3_14_2),
		.in_wire_3_3(vertical_tile_2_14_to_tile_3_14_3),
		.out_wire_1_0(vertical_tile_3_14_to_tile_4_14_0),
		.out_wire_1_1(vertical_tile_3_14_to_tile_4_14_1),
		.out_wire_1_2(vertical_tile_3_14_to_tile_4_14_2),
		.out_wire_1_3(vertical_tile_3_14_to_tile_4_14_3),
		.in_wire_1_0(vertical_tile_4_14_to_tile_3_14_0),
		.in_wire_1_1(vertical_tile_4_14_to_tile_3_14_1),
		.in_wire_1_2(vertical_tile_4_14_to_tile_3_14_2),
		.in_wire_1_3(vertical_tile_4_14_to_tile_3_14_3),
		.out_wire_2_0(horizontal_tile_3_14_to_tile_3_13_0),
		.out_wire_2_1(horizontal_tile_3_14_to_tile_3_13_1),
		.out_wire_2_2(horizontal_tile_3_14_to_tile_3_13_2),
		.out_wire_2_3(horizontal_tile_3_14_to_tile_3_13_3),
		.in_wire_2_0(horizontal_tile_3_13_to_tile_3_14_0),
		.in_wire_2_1(horizontal_tile_3_13_to_tile_3_14_1),
		.in_wire_2_2(horizontal_tile_3_13_to_tile_3_14_2),
		.in_wire_2_3(horizontal_tile_3_13_to_tile_3_14_3),
		.out_wire_0_0(horizontal_tile_3_14_to_tile_3_15_0),
		.out_wire_0_1(horizontal_tile_3_14_to_tile_3_15_1),
		.out_wire_0_2(horizontal_tile_3_14_to_tile_3_15_2),
		.out_wire_0_3(horizontal_tile_3_14_to_tile_3_15_3),
		.in_wire_0_0(horizontal_tile_3_15_to_tile_3_14_0),
		.in_wire_0_1(horizontal_tile_3_15_to_tile_3_14_1),
		.in_wire_0_2(horizontal_tile_3_15_to_tile_3_14_2),
		.in_wire_0_3(horizontal_tile_3_15_to_tile_3_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(111)
	);

	pe_tile pe_tile_3_15(
		.out_wire_3_0(vertical_tile_3_15_to_tile_2_15_0),
		.out_wire_3_1(vertical_tile_3_15_to_tile_2_15_1),
		.out_wire_3_2(vertical_tile_3_15_to_tile_2_15_2),
		.out_wire_3_3(vertical_tile_3_15_to_tile_2_15_3),
		.in_wire_3_0(vertical_tile_2_15_to_tile_3_15_0),
		.in_wire_3_1(vertical_tile_2_15_to_tile_3_15_1),
		.in_wire_3_2(vertical_tile_2_15_to_tile_3_15_2),
		.in_wire_3_3(vertical_tile_2_15_to_tile_3_15_3),
		.out_wire_1_0(vertical_tile_3_15_to_tile_4_15_0),
		.out_wire_1_1(vertical_tile_3_15_to_tile_4_15_1),
		.out_wire_1_2(vertical_tile_3_15_to_tile_4_15_2),
		.out_wire_1_3(vertical_tile_3_15_to_tile_4_15_3),
		.in_wire_1_0(vertical_tile_4_15_to_tile_3_15_0),
		.in_wire_1_1(vertical_tile_4_15_to_tile_3_15_1),
		.in_wire_1_2(vertical_tile_4_15_to_tile_3_15_2),
		.in_wire_1_3(vertical_tile_4_15_to_tile_3_15_3),
		.out_wire_2_0(horizontal_tile_3_15_to_tile_3_14_0),
		.out_wire_2_1(horizontal_tile_3_15_to_tile_3_14_1),
		.out_wire_2_2(horizontal_tile_3_15_to_tile_3_14_2),
		.out_wire_2_3(horizontal_tile_3_15_to_tile_3_14_3),
		.in_wire_2_0(horizontal_tile_3_14_to_tile_3_15_0),
		.in_wire_2_1(horizontal_tile_3_14_to_tile_3_15_1),
		.in_wire_2_2(horizontal_tile_3_14_to_tile_3_15_2),
		.in_wire_2_3(horizontal_tile_3_14_to_tile_3_15_3),
		.out_wire_0_0(horizontal_tile_3_15_to_tile_3_16_0),
		.out_wire_0_1(horizontal_tile_3_15_to_tile_3_16_1),
		.out_wire_0_2(horizontal_tile_3_15_to_tile_3_16_2),
		.out_wire_0_3(horizontal_tile_3_15_to_tile_3_16_3),
		.in_wire_0_0(horizontal_tile_3_16_to_tile_3_15_0),
		.in_wire_0_1(horizontal_tile_3_16_to_tile_3_15_1),
		.in_wire_0_2(horizontal_tile_3_16_to_tile_3_15_2),
		.in_wire_0_3(horizontal_tile_3_16_to_tile_3_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(112)
	);

	pe_tile pe_tile_3_16(
		.out_wire_3_0(vertical_tile_3_16_to_tile_2_16_0),
		.out_wire_3_1(vertical_tile_3_16_to_tile_2_16_1),
		.out_wire_3_2(vertical_tile_3_16_to_tile_2_16_2),
		.out_wire_3_3(vertical_tile_3_16_to_tile_2_16_3),
		.in_wire_3_0(vertical_tile_2_16_to_tile_3_16_0),
		.in_wire_3_1(vertical_tile_2_16_to_tile_3_16_1),
		.in_wire_3_2(vertical_tile_2_16_to_tile_3_16_2),
		.in_wire_3_3(vertical_tile_2_16_to_tile_3_16_3),
		.out_wire_1_0(vertical_tile_3_16_to_tile_4_16_0),
		.out_wire_1_1(vertical_tile_3_16_to_tile_4_16_1),
		.out_wire_1_2(vertical_tile_3_16_to_tile_4_16_2),
		.out_wire_1_3(vertical_tile_3_16_to_tile_4_16_3),
		.in_wire_1_0(vertical_tile_4_16_to_tile_3_16_0),
		.in_wire_1_1(vertical_tile_4_16_to_tile_3_16_1),
		.in_wire_1_2(vertical_tile_4_16_to_tile_3_16_2),
		.in_wire_1_3(vertical_tile_4_16_to_tile_3_16_3),
		.out_wire_2_0(horizontal_tile_3_16_to_tile_3_15_0),
		.out_wire_2_1(horizontal_tile_3_16_to_tile_3_15_1),
		.out_wire_2_2(horizontal_tile_3_16_to_tile_3_15_2),
		.out_wire_2_3(horizontal_tile_3_16_to_tile_3_15_3),
		.in_wire_2_0(horizontal_tile_3_15_to_tile_3_16_0),
		.in_wire_2_1(horizontal_tile_3_15_to_tile_3_16_1),
		.in_wire_2_2(horizontal_tile_3_15_to_tile_3_16_2),
		.in_wire_2_3(horizontal_tile_3_15_to_tile_3_16_3),
		.out_wire_0_0(horizontal_tile_3_16_to_tile_3_17_0),
		.out_wire_0_1(horizontal_tile_3_16_to_tile_3_17_1),
		.out_wire_0_2(horizontal_tile_3_16_to_tile_3_17_2),
		.out_wire_0_3(horizontal_tile_3_16_to_tile_3_17_3),
		.in_wire_0_0(horizontal_tile_3_17_to_tile_3_16_0),
		.in_wire_0_1(horizontal_tile_3_17_to_tile_3_16_1),
		.in_wire_0_2(horizontal_tile_3_17_to_tile_3_16_2),
		.in_wire_0_3(horizontal_tile_3_17_to_tile_3_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(113)
	);

	pe_tile pe_tile_3_17(
		.out_wire_3_0(vertical_tile_3_17_to_tile_2_17_0),
		.out_wire_3_1(vertical_tile_3_17_to_tile_2_17_1),
		.out_wire_3_2(vertical_tile_3_17_to_tile_2_17_2),
		.out_wire_3_3(vertical_tile_3_17_to_tile_2_17_3),
		.in_wire_3_0(vertical_tile_2_17_to_tile_3_17_0),
		.in_wire_3_1(vertical_tile_2_17_to_tile_3_17_1),
		.in_wire_3_2(vertical_tile_2_17_to_tile_3_17_2),
		.in_wire_3_3(vertical_tile_2_17_to_tile_3_17_3),
		.out_wire_1_0(vertical_tile_3_17_to_tile_4_17_0),
		.out_wire_1_1(vertical_tile_3_17_to_tile_4_17_1),
		.out_wire_1_2(vertical_tile_3_17_to_tile_4_17_2),
		.out_wire_1_3(vertical_tile_3_17_to_tile_4_17_3),
		.in_wire_1_0(vertical_tile_4_17_to_tile_3_17_0),
		.in_wire_1_1(vertical_tile_4_17_to_tile_3_17_1),
		.in_wire_1_2(vertical_tile_4_17_to_tile_3_17_2),
		.in_wire_1_3(vertical_tile_4_17_to_tile_3_17_3),
		.out_wire_2_0(horizontal_tile_3_17_to_tile_3_16_0),
		.out_wire_2_1(horizontal_tile_3_17_to_tile_3_16_1),
		.out_wire_2_2(horizontal_tile_3_17_to_tile_3_16_2),
		.out_wire_2_3(horizontal_tile_3_17_to_tile_3_16_3),
		.in_wire_2_0(horizontal_tile_3_16_to_tile_3_17_0),
		.in_wire_2_1(horizontal_tile_3_16_to_tile_3_17_1),
		.in_wire_2_2(horizontal_tile_3_16_to_tile_3_17_2),
		.in_wire_2_3(horizontal_tile_3_16_to_tile_3_17_3),
		.out_wire_0_0(horizontal_tile_3_17_to_tile_3_18_0),
		.out_wire_0_1(horizontal_tile_3_17_to_tile_3_18_1),
		.out_wire_0_2(horizontal_tile_3_17_to_tile_3_18_2),
		.out_wire_0_3(horizontal_tile_3_17_to_tile_3_18_3),
		.in_wire_0_0(horizontal_tile_3_18_to_tile_3_17_0),
		.in_wire_0_1(horizontal_tile_3_18_to_tile_3_17_1),
		.in_wire_0_2(horizontal_tile_3_18_to_tile_3_17_2),
		.in_wire_0_3(horizontal_tile_3_18_to_tile_3_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(114)
	);

	pe_tile pe_tile_3_18(
		.out_wire_3_0(vertical_tile_3_18_to_tile_2_18_0),
		.out_wire_3_1(vertical_tile_3_18_to_tile_2_18_1),
		.out_wire_3_2(vertical_tile_3_18_to_tile_2_18_2),
		.out_wire_3_3(vertical_tile_3_18_to_tile_2_18_3),
		.in_wire_3_0(vertical_tile_2_18_to_tile_3_18_0),
		.in_wire_3_1(vertical_tile_2_18_to_tile_3_18_1),
		.in_wire_3_2(vertical_tile_2_18_to_tile_3_18_2),
		.in_wire_3_3(vertical_tile_2_18_to_tile_3_18_3),
		.out_wire_1_0(vertical_tile_3_18_to_tile_4_18_0),
		.out_wire_1_1(vertical_tile_3_18_to_tile_4_18_1),
		.out_wire_1_2(vertical_tile_3_18_to_tile_4_18_2),
		.out_wire_1_3(vertical_tile_3_18_to_tile_4_18_3),
		.in_wire_1_0(vertical_tile_4_18_to_tile_3_18_0),
		.in_wire_1_1(vertical_tile_4_18_to_tile_3_18_1),
		.in_wire_1_2(vertical_tile_4_18_to_tile_3_18_2),
		.in_wire_1_3(vertical_tile_4_18_to_tile_3_18_3),
		.out_wire_2_0(horizontal_tile_3_18_to_tile_3_17_0),
		.out_wire_2_1(horizontal_tile_3_18_to_tile_3_17_1),
		.out_wire_2_2(horizontal_tile_3_18_to_tile_3_17_2),
		.out_wire_2_3(horizontal_tile_3_18_to_tile_3_17_3),
		.in_wire_2_0(horizontal_tile_3_17_to_tile_3_18_0),
		.in_wire_2_1(horizontal_tile_3_17_to_tile_3_18_1),
		.in_wire_2_2(horizontal_tile_3_17_to_tile_3_18_2),
		.in_wire_2_3(horizontal_tile_3_17_to_tile_3_18_3),
		.out_wire_0_0(horizontal_tile_3_18_to_tile_3_19_0),
		.out_wire_0_1(horizontal_tile_3_18_to_tile_3_19_1),
		.out_wire_0_2(horizontal_tile_3_18_to_tile_3_19_2),
		.out_wire_0_3(horizontal_tile_3_18_to_tile_3_19_3),
		.in_wire_0_0(horizontal_tile_3_19_to_tile_3_18_0),
		.in_wire_0_1(horizontal_tile_3_19_to_tile_3_18_1),
		.in_wire_0_2(horizontal_tile_3_19_to_tile_3_18_2),
		.in_wire_0_3(horizontal_tile_3_19_to_tile_3_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(115)
	);

	pe_tile pe_tile_3_19(
		.out_wire_3_0(vertical_tile_3_19_to_tile_2_19_0),
		.out_wire_3_1(vertical_tile_3_19_to_tile_2_19_1),
		.out_wire_3_2(vertical_tile_3_19_to_tile_2_19_2),
		.out_wire_3_3(vertical_tile_3_19_to_tile_2_19_3),
		.in_wire_3_0(vertical_tile_2_19_to_tile_3_19_0),
		.in_wire_3_1(vertical_tile_2_19_to_tile_3_19_1),
		.in_wire_3_2(vertical_tile_2_19_to_tile_3_19_2),
		.in_wire_3_3(vertical_tile_2_19_to_tile_3_19_3),
		.out_wire_1_0(vertical_tile_3_19_to_tile_4_19_0),
		.out_wire_1_1(vertical_tile_3_19_to_tile_4_19_1),
		.out_wire_1_2(vertical_tile_3_19_to_tile_4_19_2),
		.out_wire_1_3(vertical_tile_3_19_to_tile_4_19_3),
		.in_wire_1_0(vertical_tile_4_19_to_tile_3_19_0),
		.in_wire_1_1(vertical_tile_4_19_to_tile_3_19_1),
		.in_wire_1_2(vertical_tile_4_19_to_tile_3_19_2),
		.in_wire_1_3(vertical_tile_4_19_to_tile_3_19_3),
		.out_wire_2_0(horizontal_tile_3_19_to_tile_3_18_0),
		.out_wire_2_1(horizontal_tile_3_19_to_tile_3_18_1),
		.out_wire_2_2(horizontal_tile_3_19_to_tile_3_18_2),
		.out_wire_2_3(horizontal_tile_3_19_to_tile_3_18_3),
		.in_wire_2_0(horizontal_tile_3_18_to_tile_3_19_0),
		.in_wire_2_1(horizontal_tile_3_18_to_tile_3_19_1),
		.in_wire_2_2(horizontal_tile_3_18_to_tile_3_19_2),
		.in_wire_2_3(horizontal_tile_3_18_to_tile_3_19_3),
		.out_wire_0_0(horizontal_tile_3_19_to_tile_3_20_0),
		.out_wire_0_1(horizontal_tile_3_19_to_tile_3_20_1),
		.out_wire_0_2(horizontal_tile_3_19_to_tile_3_20_2),
		.out_wire_0_3(horizontal_tile_3_19_to_tile_3_20_3),
		.in_wire_0_0(horizontal_tile_3_20_to_tile_3_19_0),
		.in_wire_0_1(horizontal_tile_3_20_to_tile_3_19_1),
		.in_wire_0_2(horizontal_tile_3_20_to_tile_3_19_2),
		.in_wire_0_3(horizontal_tile_3_20_to_tile_3_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(116)
	);

	pe_tile pe_tile_3_20(
		.out_wire_3_0(vertical_tile_3_20_to_tile_2_20_0),
		.out_wire_3_1(vertical_tile_3_20_to_tile_2_20_1),
		.out_wire_3_2(vertical_tile_3_20_to_tile_2_20_2),
		.out_wire_3_3(vertical_tile_3_20_to_tile_2_20_3),
		.in_wire_3_0(vertical_tile_2_20_to_tile_3_20_0),
		.in_wire_3_1(vertical_tile_2_20_to_tile_3_20_1),
		.in_wire_3_2(vertical_tile_2_20_to_tile_3_20_2),
		.in_wire_3_3(vertical_tile_2_20_to_tile_3_20_3),
		.out_wire_1_0(vertical_tile_3_20_to_tile_4_20_0),
		.out_wire_1_1(vertical_tile_3_20_to_tile_4_20_1),
		.out_wire_1_2(vertical_tile_3_20_to_tile_4_20_2),
		.out_wire_1_3(vertical_tile_3_20_to_tile_4_20_3),
		.in_wire_1_0(vertical_tile_4_20_to_tile_3_20_0),
		.in_wire_1_1(vertical_tile_4_20_to_tile_3_20_1),
		.in_wire_1_2(vertical_tile_4_20_to_tile_3_20_2),
		.in_wire_1_3(vertical_tile_4_20_to_tile_3_20_3),
		.out_wire_2_0(horizontal_tile_3_20_to_tile_3_19_0),
		.out_wire_2_1(horizontal_tile_3_20_to_tile_3_19_1),
		.out_wire_2_2(horizontal_tile_3_20_to_tile_3_19_2),
		.out_wire_2_3(horizontal_tile_3_20_to_tile_3_19_3),
		.in_wire_2_0(horizontal_tile_3_19_to_tile_3_20_0),
		.in_wire_2_1(horizontal_tile_3_19_to_tile_3_20_1),
		.in_wire_2_2(horizontal_tile_3_19_to_tile_3_20_2),
		.in_wire_2_3(horizontal_tile_3_19_to_tile_3_20_3),
		.out_wire_0_0(horizontal_tile_3_20_to_tile_3_21_0),
		.out_wire_0_1(horizontal_tile_3_20_to_tile_3_21_1),
		.out_wire_0_2(horizontal_tile_3_20_to_tile_3_21_2),
		.out_wire_0_3(horizontal_tile_3_20_to_tile_3_21_3),
		.in_wire_0_0(horizontal_tile_3_21_to_tile_3_20_0),
		.in_wire_0_1(horizontal_tile_3_21_to_tile_3_20_1),
		.in_wire_0_2(horizontal_tile_3_21_to_tile_3_20_2),
		.in_wire_0_3(horizontal_tile_3_21_to_tile_3_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(117)
	);

	pe_tile pe_tile_3_21(
		.out_wire_3_0(vertical_tile_3_21_to_tile_2_21_0),
		.out_wire_3_1(vertical_tile_3_21_to_tile_2_21_1),
		.out_wire_3_2(vertical_tile_3_21_to_tile_2_21_2),
		.out_wire_3_3(vertical_tile_3_21_to_tile_2_21_3),
		.in_wire_3_0(vertical_tile_2_21_to_tile_3_21_0),
		.in_wire_3_1(vertical_tile_2_21_to_tile_3_21_1),
		.in_wire_3_2(vertical_tile_2_21_to_tile_3_21_2),
		.in_wire_3_3(vertical_tile_2_21_to_tile_3_21_3),
		.out_wire_1_0(vertical_tile_3_21_to_tile_4_21_0),
		.out_wire_1_1(vertical_tile_3_21_to_tile_4_21_1),
		.out_wire_1_2(vertical_tile_3_21_to_tile_4_21_2),
		.out_wire_1_3(vertical_tile_3_21_to_tile_4_21_3),
		.in_wire_1_0(vertical_tile_4_21_to_tile_3_21_0),
		.in_wire_1_1(vertical_tile_4_21_to_tile_3_21_1),
		.in_wire_1_2(vertical_tile_4_21_to_tile_3_21_2),
		.in_wire_1_3(vertical_tile_4_21_to_tile_3_21_3),
		.out_wire_2_0(horizontal_tile_3_21_to_tile_3_20_0),
		.out_wire_2_1(horizontal_tile_3_21_to_tile_3_20_1),
		.out_wire_2_2(horizontal_tile_3_21_to_tile_3_20_2),
		.out_wire_2_3(horizontal_tile_3_21_to_tile_3_20_3),
		.in_wire_2_0(horizontal_tile_3_20_to_tile_3_21_0),
		.in_wire_2_1(horizontal_tile_3_20_to_tile_3_21_1),
		.in_wire_2_2(horizontal_tile_3_20_to_tile_3_21_2),
		.in_wire_2_3(horizontal_tile_3_20_to_tile_3_21_3),
		.out_wire_0_0(horizontal_tile_3_21_to_tile_3_22_0),
		.out_wire_0_1(horizontal_tile_3_21_to_tile_3_22_1),
		.out_wire_0_2(horizontal_tile_3_21_to_tile_3_22_2),
		.out_wire_0_3(horizontal_tile_3_21_to_tile_3_22_3),
		.in_wire_0_0(horizontal_tile_3_22_to_tile_3_21_0),
		.in_wire_0_1(horizontal_tile_3_22_to_tile_3_21_1),
		.in_wire_0_2(horizontal_tile_3_22_to_tile_3_21_2),
		.in_wire_0_3(horizontal_tile_3_22_to_tile_3_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(118)
	);

	pe_tile pe_tile_3_22(
		.out_wire_3_0(vertical_tile_3_22_to_tile_2_22_0),
		.out_wire_3_1(vertical_tile_3_22_to_tile_2_22_1),
		.out_wire_3_2(vertical_tile_3_22_to_tile_2_22_2),
		.out_wire_3_3(vertical_tile_3_22_to_tile_2_22_3),
		.in_wire_3_0(vertical_tile_2_22_to_tile_3_22_0),
		.in_wire_3_1(vertical_tile_2_22_to_tile_3_22_1),
		.in_wire_3_2(vertical_tile_2_22_to_tile_3_22_2),
		.in_wire_3_3(vertical_tile_2_22_to_tile_3_22_3),
		.out_wire_1_0(vertical_tile_3_22_to_tile_4_22_0),
		.out_wire_1_1(vertical_tile_3_22_to_tile_4_22_1),
		.out_wire_1_2(vertical_tile_3_22_to_tile_4_22_2),
		.out_wire_1_3(vertical_tile_3_22_to_tile_4_22_3),
		.in_wire_1_0(vertical_tile_4_22_to_tile_3_22_0),
		.in_wire_1_1(vertical_tile_4_22_to_tile_3_22_1),
		.in_wire_1_2(vertical_tile_4_22_to_tile_3_22_2),
		.in_wire_1_3(vertical_tile_4_22_to_tile_3_22_3),
		.out_wire_2_0(horizontal_tile_3_22_to_tile_3_21_0),
		.out_wire_2_1(horizontal_tile_3_22_to_tile_3_21_1),
		.out_wire_2_2(horizontal_tile_3_22_to_tile_3_21_2),
		.out_wire_2_3(horizontal_tile_3_22_to_tile_3_21_3),
		.in_wire_2_0(horizontal_tile_3_21_to_tile_3_22_0),
		.in_wire_2_1(horizontal_tile_3_21_to_tile_3_22_1),
		.in_wire_2_2(horizontal_tile_3_21_to_tile_3_22_2),
		.in_wire_2_3(horizontal_tile_3_21_to_tile_3_22_3),
		.out_wire_0_0(horizontal_tile_3_22_to_tile_3_23_0),
		.out_wire_0_1(horizontal_tile_3_22_to_tile_3_23_1),
		.out_wire_0_2(horizontal_tile_3_22_to_tile_3_23_2),
		.out_wire_0_3(horizontal_tile_3_22_to_tile_3_23_3),
		.in_wire_0_0(horizontal_tile_3_23_to_tile_3_22_0),
		.in_wire_0_1(horizontal_tile_3_23_to_tile_3_22_1),
		.in_wire_0_2(horizontal_tile_3_23_to_tile_3_22_2),
		.in_wire_0_3(horizontal_tile_3_23_to_tile_3_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(119)
	);

	pe_tile pe_tile_3_23(
		.out_wire_3_0(vertical_tile_3_23_to_tile_2_23_0),
		.out_wire_3_1(vertical_tile_3_23_to_tile_2_23_1),
		.out_wire_3_2(vertical_tile_3_23_to_tile_2_23_2),
		.out_wire_3_3(vertical_tile_3_23_to_tile_2_23_3),
		.in_wire_3_0(vertical_tile_2_23_to_tile_3_23_0),
		.in_wire_3_1(vertical_tile_2_23_to_tile_3_23_1),
		.in_wire_3_2(vertical_tile_2_23_to_tile_3_23_2),
		.in_wire_3_3(vertical_tile_2_23_to_tile_3_23_3),
		.out_wire_1_0(vertical_tile_3_23_to_tile_4_23_0),
		.out_wire_1_1(vertical_tile_3_23_to_tile_4_23_1),
		.out_wire_1_2(vertical_tile_3_23_to_tile_4_23_2),
		.out_wire_1_3(vertical_tile_3_23_to_tile_4_23_3),
		.in_wire_1_0(vertical_tile_4_23_to_tile_3_23_0),
		.in_wire_1_1(vertical_tile_4_23_to_tile_3_23_1),
		.in_wire_1_2(vertical_tile_4_23_to_tile_3_23_2),
		.in_wire_1_3(vertical_tile_4_23_to_tile_3_23_3),
		.out_wire_2_0(horizontal_tile_3_23_to_tile_3_22_0),
		.out_wire_2_1(horizontal_tile_3_23_to_tile_3_22_1),
		.out_wire_2_2(horizontal_tile_3_23_to_tile_3_22_2),
		.out_wire_2_3(horizontal_tile_3_23_to_tile_3_22_3),
		.in_wire_2_0(horizontal_tile_3_22_to_tile_3_23_0),
		.in_wire_2_1(horizontal_tile_3_22_to_tile_3_23_1),
		.in_wire_2_2(horizontal_tile_3_22_to_tile_3_23_2),
		.in_wire_2_3(horizontal_tile_3_22_to_tile_3_23_3),
		.out_wire_0_0(horizontal_tile_3_23_to_tile_3_24_0),
		.out_wire_0_1(horizontal_tile_3_23_to_tile_3_24_1),
		.out_wire_0_2(horizontal_tile_3_23_to_tile_3_24_2),
		.out_wire_0_3(horizontal_tile_3_23_to_tile_3_24_3),
		.in_wire_0_0(horizontal_tile_3_24_to_tile_3_23_0),
		.in_wire_0_1(horizontal_tile_3_24_to_tile_3_23_1),
		.in_wire_0_2(horizontal_tile_3_24_to_tile_3_23_2),
		.in_wire_0_3(horizontal_tile_3_24_to_tile_3_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(120)
	);

	pe_tile pe_tile_3_24(
		.out_wire_3_0(vertical_tile_3_24_to_tile_2_24_0),
		.out_wire_3_1(vertical_tile_3_24_to_tile_2_24_1),
		.out_wire_3_2(vertical_tile_3_24_to_tile_2_24_2),
		.out_wire_3_3(vertical_tile_3_24_to_tile_2_24_3),
		.in_wire_3_0(vertical_tile_2_24_to_tile_3_24_0),
		.in_wire_3_1(vertical_tile_2_24_to_tile_3_24_1),
		.in_wire_3_2(vertical_tile_2_24_to_tile_3_24_2),
		.in_wire_3_3(vertical_tile_2_24_to_tile_3_24_3),
		.out_wire_1_0(vertical_tile_3_24_to_tile_4_24_0),
		.out_wire_1_1(vertical_tile_3_24_to_tile_4_24_1),
		.out_wire_1_2(vertical_tile_3_24_to_tile_4_24_2),
		.out_wire_1_3(vertical_tile_3_24_to_tile_4_24_3),
		.in_wire_1_0(vertical_tile_4_24_to_tile_3_24_0),
		.in_wire_1_1(vertical_tile_4_24_to_tile_3_24_1),
		.in_wire_1_2(vertical_tile_4_24_to_tile_3_24_2),
		.in_wire_1_3(vertical_tile_4_24_to_tile_3_24_3),
		.out_wire_2_0(horizontal_tile_3_24_to_tile_3_23_0),
		.out_wire_2_1(horizontal_tile_3_24_to_tile_3_23_1),
		.out_wire_2_2(horizontal_tile_3_24_to_tile_3_23_2),
		.out_wire_2_3(horizontal_tile_3_24_to_tile_3_23_3),
		.in_wire_2_0(horizontal_tile_3_23_to_tile_3_24_0),
		.in_wire_2_1(horizontal_tile_3_23_to_tile_3_24_1),
		.in_wire_2_2(horizontal_tile_3_23_to_tile_3_24_2),
		.in_wire_2_3(horizontal_tile_3_23_to_tile_3_24_3),
		.out_wire_0_0(horizontal_tile_3_24_to_tile_3_25_0),
		.out_wire_0_1(horizontal_tile_3_24_to_tile_3_25_1),
		.out_wire_0_2(horizontal_tile_3_24_to_tile_3_25_2),
		.out_wire_0_3(horizontal_tile_3_24_to_tile_3_25_3),
		.in_wire_0_0(horizontal_tile_3_25_to_tile_3_24_0),
		.in_wire_0_1(horizontal_tile_3_25_to_tile_3_24_1),
		.in_wire_0_2(horizontal_tile_3_25_to_tile_3_24_2),
		.in_wire_0_3(horizontal_tile_3_25_to_tile_3_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(121)
	);

	pe_tile pe_tile_3_25(
		.out_wire_3_0(vertical_tile_3_25_to_tile_2_25_0),
		.out_wire_3_1(vertical_tile_3_25_to_tile_2_25_1),
		.out_wire_3_2(vertical_tile_3_25_to_tile_2_25_2),
		.out_wire_3_3(vertical_tile_3_25_to_tile_2_25_3),
		.in_wire_3_0(vertical_tile_2_25_to_tile_3_25_0),
		.in_wire_3_1(vertical_tile_2_25_to_tile_3_25_1),
		.in_wire_3_2(vertical_tile_2_25_to_tile_3_25_2),
		.in_wire_3_3(vertical_tile_2_25_to_tile_3_25_3),
		.out_wire_1_0(vertical_tile_3_25_to_tile_4_25_0),
		.out_wire_1_1(vertical_tile_3_25_to_tile_4_25_1),
		.out_wire_1_2(vertical_tile_3_25_to_tile_4_25_2),
		.out_wire_1_3(vertical_tile_3_25_to_tile_4_25_3),
		.in_wire_1_0(vertical_tile_4_25_to_tile_3_25_0),
		.in_wire_1_1(vertical_tile_4_25_to_tile_3_25_1),
		.in_wire_1_2(vertical_tile_4_25_to_tile_3_25_2),
		.in_wire_1_3(vertical_tile_4_25_to_tile_3_25_3),
		.out_wire_2_0(horizontal_tile_3_25_to_tile_3_24_0),
		.out_wire_2_1(horizontal_tile_3_25_to_tile_3_24_1),
		.out_wire_2_2(horizontal_tile_3_25_to_tile_3_24_2),
		.out_wire_2_3(horizontal_tile_3_25_to_tile_3_24_3),
		.in_wire_2_0(horizontal_tile_3_24_to_tile_3_25_0),
		.in_wire_2_1(horizontal_tile_3_24_to_tile_3_25_1),
		.in_wire_2_2(horizontal_tile_3_24_to_tile_3_25_2),
		.in_wire_2_3(horizontal_tile_3_24_to_tile_3_25_3),
		.out_wire_0_0(horizontal_tile_3_25_to_tile_3_26_0),
		.out_wire_0_1(horizontal_tile_3_25_to_tile_3_26_1),
		.out_wire_0_2(horizontal_tile_3_25_to_tile_3_26_2),
		.out_wire_0_3(horizontal_tile_3_25_to_tile_3_26_3),
		.in_wire_0_0(horizontal_tile_3_26_to_tile_3_25_0),
		.in_wire_0_1(horizontal_tile_3_26_to_tile_3_25_1),
		.in_wire_0_2(horizontal_tile_3_26_to_tile_3_25_2),
		.in_wire_0_3(horizontal_tile_3_26_to_tile_3_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(122)
	);

	pe_tile pe_tile_3_26(
		.out_wire_3_0(vertical_tile_3_26_to_tile_2_26_0),
		.out_wire_3_1(vertical_tile_3_26_to_tile_2_26_1),
		.out_wire_3_2(vertical_tile_3_26_to_tile_2_26_2),
		.out_wire_3_3(vertical_tile_3_26_to_tile_2_26_3),
		.in_wire_3_0(vertical_tile_2_26_to_tile_3_26_0),
		.in_wire_3_1(vertical_tile_2_26_to_tile_3_26_1),
		.in_wire_3_2(vertical_tile_2_26_to_tile_3_26_2),
		.in_wire_3_3(vertical_tile_2_26_to_tile_3_26_3),
		.out_wire_1_0(vertical_tile_3_26_to_tile_4_26_0),
		.out_wire_1_1(vertical_tile_3_26_to_tile_4_26_1),
		.out_wire_1_2(vertical_tile_3_26_to_tile_4_26_2),
		.out_wire_1_3(vertical_tile_3_26_to_tile_4_26_3),
		.in_wire_1_0(vertical_tile_4_26_to_tile_3_26_0),
		.in_wire_1_1(vertical_tile_4_26_to_tile_3_26_1),
		.in_wire_1_2(vertical_tile_4_26_to_tile_3_26_2),
		.in_wire_1_3(vertical_tile_4_26_to_tile_3_26_3),
		.out_wire_2_0(horizontal_tile_3_26_to_tile_3_25_0),
		.out_wire_2_1(horizontal_tile_3_26_to_tile_3_25_1),
		.out_wire_2_2(horizontal_tile_3_26_to_tile_3_25_2),
		.out_wire_2_3(horizontal_tile_3_26_to_tile_3_25_3),
		.in_wire_2_0(horizontal_tile_3_25_to_tile_3_26_0),
		.in_wire_2_1(horizontal_tile_3_25_to_tile_3_26_1),
		.in_wire_2_2(horizontal_tile_3_25_to_tile_3_26_2),
		.in_wire_2_3(horizontal_tile_3_25_to_tile_3_26_3),
		.out_wire_0_0(horizontal_tile_3_26_to_tile_3_27_0),
		.out_wire_0_1(horizontal_tile_3_26_to_tile_3_27_1),
		.out_wire_0_2(horizontal_tile_3_26_to_tile_3_27_2),
		.out_wire_0_3(horizontal_tile_3_26_to_tile_3_27_3),
		.in_wire_0_0(horizontal_tile_3_27_to_tile_3_26_0),
		.in_wire_0_1(horizontal_tile_3_27_to_tile_3_26_1),
		.in_wire_0_2(horizontal_tile_3_27_to_tile_3_26_2),
		.in_wire_0_3(horizontal_tile_3_27_to_tile_3_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(123)
	);

	pe_tile pe_tile_3_27(
		.out_wire_3_0(vertical_tile_3_27_to_tile_2_27_0),
		.out_wire_3_1(vertical_tile_3_27_to_tile_2_27_1),
		.out_wire_3_2(vertical_tile_3_27_to_tile_2_27_2),
		.out_wire_3_3(vertical_tile_3_27_to_tile_2_27_3),
		.in_wire_3_0(vertical_tile_2_27_to_tile_3_27_0),
		.in_wire_3_1(vertical_tile_2_27_to_tile_3_27_1),
		.in_wire_3_2(vertical_tile_2_27_to_tile_3_27_2),
		.in_wire_3_3(vertical_tile_2_27_to_tile_3_27_3),
		.out_wire_1_0(vertical_tile_3_27_to_tile_4_27_0),
		.out_wire_1_1(vertical_tile_3_27_to_tile_4_27_1),
		.out_wire_1_2(vertical_tile_3_27_to_tile_4_27_2),
		.out_wire_1_3(vertical_tile_3_27_to_tile_4_27_3),
		.in_wire_1_0(vertical_tile_4_27_to_tile_3_27_0),
		.in_wire_1_1(vertical_tile_4_27_to_tile_3_27_1),
		.in_wire_1_2(vertical_tile_4_27_to_tile_3_27_2),
		.in_wire_1_3(vertical_tile_4_27_to_tile_3_27_3),
		.out_wire_2_0(horizontal_tile_3_27_to_tile_3_26_0),
		.out_wire_2_1(horizontal_tile_3_27_to_tile_3_26_1),
		.out_wire_2_2(horizontal_tile_3_27_to_tile_3_26_2),
		.out_wire_2_3(horizontal_tile_3_27_to_tile_3_26_3),
		.in_wire_2_0(horizontal_tile_3_26_to_tile_3_27_0),
		.in_wire_2_1(horizontal_tile_3_26_to_tile_3_27_1),
		.in_wire_2_2(horizontal_tile_3_26_to_tile_3_27_2),
		.in_wire_2_3(horizontal_tile_3_26_to_tile_3_27_3),
		.out_wire_0_0(horizontal_tile_3_27_to_tile_3_28_0),
		.out_wire_0_1(horizontal_tile_3_27_to_tile_3_28_1),
		.out_wire_0_2(horizontal_tile_3_27_to_tile_3_28_2),
		.out_wire_0_3(horizontal_tile_3_27_to_tile_3_28_3),
		.in_wire_0_0(horizontal_tile_3_28_to_tile_3_27_0),
		.in_wire_0_1(horizontal_tile_3_28_to_tile_3_27_1),
		.in_wire_0_2(horizontal_tile_3_28_to_tile_3_27_2),
		.in_wire_0_3(horizontal_tile_3_28_to_tile_3_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(124)
	);

	pe_tile pe_tile_3_28(
		.out_wire_3_0(vertical_tile_3_28_to_tile_2_28_0),
		.out_wire_3_1(vertical_tile_3_28_to_tile_2_28_1),
		.out_wire_3_2(vertical_tile_3_28_to_tile_2_28_2),
		.out_wire_3_3(vertical_tile_3_28_to_tile_2_28_3),
		.in_wire_3_0(vertical_tile_2_28_to_tile_3_28_0),
		.in_wire_3_1(vertical_tile_2_28_to_tile_3_28_1),
		.in_wire_3_2(vertical_tile_2_28_to_tile_3_28_2),
		.in_wire_3_3(vertical_tile_2_28_to_tile_3_28_3),
		.out_wire_1_0(vertical_tile_3_28_to_tile_4_28_0),
		.out_wire_1_1(vertical_tile_3_28_to_tile_4_28_1),
		.out_wire_1_2(vertical_tile_3_28_to_tile_4_28_2),
		.out_wire_1_3(vertical_tile_3_28_to_tile_4_28_3),
		.in_wire_1_0(vertical_tile_4_28_to_tile_3_28_0),
		.in_wire_1_1(vertical_tile_4_28_to_tile_3_28_1),
		.in_wire_1_2(vertical_tile_4_28_to_tile_3_28_2),
		.in_wire_1_3(vertical_tile_4_28_to_tile_3_28_3),
		.out_wire_2_0(horizontal_tile_3_28_to_tile_3_27_0),
		.out_wire_2_1(horizontal_tile_3_28_to_tile_3_27_1),
		.out_wire_2_2(horizontal_tile_3_28_to_tile_3_27_2),
		.out_wire_2_3(horizontal_tile_3_28_to_tile_3_27_3),
		.in_wire_2_0(horizontal_tile_3_27_to_tile_3_28_0),
		.in_wire_2_1(horizontal_tile_3_27_to_tile_3_28_1),
		.in_wire_2_2(horizontal_tile_3_27_to_tile_3_28_2),
		.in_wire_2_3(horizontal_tile_3_27_to_tile_3_28_3),
		.out_wire_0_0(horizontal_tile_3_28_to_tile_3_29_0),
		.out_wire_0_1(horizontal_tile_3_28_to_tile_3_29_1),
		.out_wire_0_2(horizontal_tile_3_28_to_tile_3_29_2),
		.out_wire_0_3(horizontal_tile_3_28_to_tile_3_29_3),
		.in_wire_0_0(horizontal_tile_3_29_to_tile_3_28_0),
		.in_wire_0_1(horizontal_tile_3_29_to_tile_3_28_1),
		.in_wire_0_2(horizontal_tile_3_29_to_tile_3_28_2),
		.in_wire_0_3(horizontal_tile_3_29_to_tile_3_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(125)
	);

	pe_tile pe_tile_3_29(
		.out_wire_3_0(vertical_tile_3_29_to_tile_2_29_0),
		.out_wire_3_1(vertical_tile_3_29_to_tile_2_29_1),
		.out_wire_3_2(vertical_tile_3_29_to_tile_2_29_2),
		.out_wire_3_3(vertical_tile_3_29_to_tile_2_29_3),
		.in_wire_3_0(vertical_tile_2_29_to_tile_3_29_0),
		.in_wire_3_1(vertical_tile_2_29_to_tile_3_29_1),
		.in_wire_3_2(vertical_tile_2_29_to_tile_3_29_2),
		.in_wire_3_3(vertical_tile_2_29_to_tile_3_29_3),
		.out_wire_1_0(vertical_tile_3_29_to_tile_4_29_0),
		.out_wire_1_1(vertical_tile_3_29_to_tile_4_29_1),
		.out_wire_1_2(vertical_tile_3_29_to_tile_4_29_2),
		.out_wire_1_3(vertical_tile_3_29_to_tile_4_29_3),
		.in_wire_1_0(vertical_tile_4_29_to_tile_3_29_0),
		.in_wire_1_1(vertical_tile_4_29_to_tile_3_29_1),
		.in_wire_1_2(vertical_tile_4_29_to_tile_3_29_2),
		.in_wire_1_3(vertical_tile_4_29_to_tile_3_29_3),
		.out_wire_2_0(horizontal_tile_3_29_to_tile_3_28_0),
		.out_wire_2_1(horizontal_tile_3_29_to_tile_3_28_1),
		.out_wire_2_2(horizontal_tile_3_29_to_tile_3_28_2),
		.out_wire_2_3(horizontal_tile_3_29_to_tile_3_28_3),
		.in_wire_2_0(horizontal_tile_3_28_to_tile_3_29_0),
		.in_wire_2_1(horizontal_tile_3_28_to_tile_3_29_1),
		.in_wire_2_2(horizontal_tile_3_28_to_tile_3_29_2),
		.in_wire_2_3(horizontal_tile_3_28_to_tile_3_29_3),
		.out_wire_0_0(horizontal_tile_3_29_to_tile_3_30_0),
		.out_wire_0_1(horizontal_tile_3_29_to_tile_3_30_1),
		.out_wire_0_2(horizontal_tile_3_29_to_tile_3_30_2),
		.out_wire_0_3(horizontal_tile_3_29_to_tile_3_30_3),
		.in_wire_0_0(horizontal_tile_3_30_to_tile_3_29_0),
		.in_wire_0_1(horizontal_tile_3_30_to_tile_3_29_1),
		.in_wire_0_2(horizontal_tile_3_30_to_tile_3_29_2),
		.in_wire_0_3(horizontal_tile_3_30_to_tile_3_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(126)
	);

	pe_tile pe_tile_3_30(
		.out_wire_3_0(vertical_tile_3_30_to_tile_2_30_0),
		.out_wire_3_1(vertical_tile_3_30_to_tile_2_30_1),
		.out_wire_3_2(vertical_tile_3_30_to_tile_2_30_2),
		.out_wire_3_3(vertical_tile_3_30_to_tile_2_30_3),
		.in_wire_3_0(vertical_tile_2_30_to_tile_3_30_0),
		.in_wire_3_1(vertical_tile_2_30_to_tile_3_30_1),
		.in_wire_3_2(vertical_tile_2_30_to_tile_3_30_2),
		.in_wire_3_3(vertical_tile_2_30_to_tile_3_30_3),
		.out_wire_1_0(vertical_tile_3_30_to_tile_4_30_0),
		.out_wire_1_1(vertical_tile_3_30_to_tile_4_30_1),
		.out_wire_1_2(vertical_tile_3_30_to_tile_4_30_2),
		.out_wire_1_3(vertical_tile_3_30_to_tile_4_30_3),
		.in_wire_1_0(vertical_tile_4_30_to_tile_3_30_0),
		.in_wire_1_1(vertical_tile_4_30_to_tile_3_30_1),
		.in_wire_1_2(vertical_tile_4_30_to_tile_3_30_2),
		.in_wire_1_3(vertical_tile_4_30_to_tile_3_30_3),
		.out_wire_2_0(horizontal_tile_3_30_to_tile_3_29_0),
		.out_wire_2_1(horizontal_tile_3_30_to_tile_3_29_1),
		.out_wire_2_2(horizontal_tile_3_30_to_tile_3_29_2),
		.out_wire_2_3(horizontal_tile_3_30_to_tile_3_29_3),
		.in_wire_2_0(horizontal_tile_3_29_to_tile_3_30_0),
		.in_wire_2_1(horizontal_tile_3_29_to_tile_3_30_1),
		.in_wire_2_2(horizontal_tile_3_29_to_tile_3_30_2),
		.in_wire_2_3(horizontal_tile_3_29_to_tile_3_30_3),
		.out_wire_0_0(horizontal_tile_3_30_to_tile_3_31_0),
		.out_wire_0_1(horizontal_tile_3_30_to_tile_3_31_1),
		.out_wire_0_2(horizontal_tile_3_30_to_tile_3_31_2),
		.out_wire_0_3(horizontal_tile_3_30_to_tile_3_31_3),
		.in_wire_0_0(horizontal_tile_3_31_to_tile_3_30_0),
		.in_wire_0_1(horizontal_tile_3_31_to_tile_3_30_1),
		.in_wire_0_2(horizontal_tile_3_31_to_tile_3_30_2),
		.in_wire_0_3(horizontal_tile_3_31_to_tile_3_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(127)
	);

	pe_tile_right pe_tile_3_31(
		.out_wire_3_0(vertical_tile_3_31_to_tile_2_31_0),
		.out_wire_3_1(vertical_tile_3_31_to_tile_2_31_1),
		.out_wire_3_2(vertical_tile_3_31_to_tile_2_31_2),
		.out_wire_3_3(vertical_tile_3_31_to_tile_2_31_3),
		.in_wire_3_0(vertical_tile_2_31_to_tile_3_31_0),
		.in_wire_3_1(vertical_tile_2_31_to_tile_3_31_1),
		.in_wire_3_2(vertical_tile_2_31_to_tile_3_31_2),
		.in_wire_3_3(vertical_tile_2_31_to_tile_3_31_3),
		.out_wire_1_0(vertical_tile_3_31_to_tile_4_31_0),
		.out_wire_1_1(vertical_tile_3_31_to_tile_4_31_1),
		.out_wire_1_2(vertical_tile_3_31_to_tile_4_31_2),
		.out_wire_1_3(vertical_tile_3_31_to_tile_4_31_3),
		.in_wire_1_0(vertical_tile_4_31_to_tile_3_31_0),
		.in_wire_1_1(vertical_tile_4_31_to_tile_3_31_1),
		.in_wire_1_2(vertical_tile_4_31_to_tile_3_31_2),
		.in_wire_1_3(vertical_tile_4_31_to_tile_3_31_3),
		.out_wire_2_0(horizontal_tile_3_31_to_tile_3_30_0),
		.out_wire_2_1(horizontal_tile_3_31_to_tile_3_30_1),
		.out_wire_2_2(horizontal_tile_3_31_to_tile_3_30_2),
		.out_wire_2_3(horizontal_tile_3_31_to_tile_3_30_3),
		.in_wire_2_0(horizontal_tile_3_30_to_tile_3_31_0),
		.in_wire_2_1(horizontal_tile_3_30_to_tile_3_31_1),
		.in_wire_2_2(horizontal_tile_3_30_to_tile_3_31_2),
		.in_wire_2_3(horizontal_tile_3_30_to_tile_3_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(128)
	);

	pe_tile_left pe_tile_4_0(
		.out_wire_3_0(vertical_tile_4_0_to_tile_3_0_0),
		.out_wire_3_1(vertical_tile_4_0_to_tile_3_0_1),
		.out_wire_3_2(vertical_tile_4_0_to_tile_3_0_2),
		.out_wire_3_3(vertical_tile_4_0_to_tile_3_0_3),
		.in_wire_3_0(vertical_tile_3_0_to_tile_4_0_0),
		.in_wire_3_1(vertical_tile_3_0_to_tile_4_0_1),
		.in_wire_3_2(vertical_tile_3_0_to_tile_4_0_2),
		.in_wire_3_3(vertical_tile_3_0_to_tile_4_0_3),
		.out_wire_1_0(vertical_tile_4_0_to_tile_5_0_0),
		.out_wire_1_1(vertical_tile_4_0_to_tile_5_0_1),
		.out_wire_1_2(vertical_tile_4_0_to_tile_5_0_2),
		.out_wire_1_3(vertical_tile_4_0_to_tile_5_0_3),
		.in_wire_1_0(vertical_tile_5_0_to_tile_4_0_0),
		.in_wire_1_1(vertical_tile_5_0_to_tile_4_0_1),
		.in_wire_1_2(vertical_tile_5_0_to_tile_4_0_2),
		.in_wire_1_3(vertical_tile_5_0_to_tile_4_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_4_0_to_tile_4_1_0),
		.out_wire_0_1(horizontal_tile_4_0_to_tile_4_1_1),
		.out_wire_0_2(horizontal_tile_4_0_to_tile_4_1_2),
		.out_wire_0_3(horizontal_tile_4_0_to_tile_4_1_3),
		.in_wire_0_0(horizontal_tile_4_1_to_tile_4_0_0),
		.in_wire_0_1(horizontal_tile_4_1_to_tile_4_0_1),
		.in_wire_0_2(horizontal_tile_4_1_to_tile_4_0_2),
		.in_wire_0_3(horizontal_tile_4_1_to_tile_4_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(129)
	);

	pe_tile pe_tile_4_1(
		.out_wire_3_0(vertical_tile_4_1_to_tile_3_1_0),
		.out_wire_3_1(vertical_tile_4_1_to_tile_3_1_1),
		.out_wire_3_2(vertical_tile_4_1_to_tile_3_1_2),
		.out_wire_3_3(vertical_tile_4_1_to_tile_3_1_3),
		.in_wire_3_0(vertical_tile_3_1_to_tile_4_1_0),
		.in_wire_3_1(vertical_tile_3_1_to_tile_4_1_1),
		.in_wire_3_2(vertical_tile_3_1_to_tile_4_1_2),
		.in_wire_3_3(vertical_tile_3_1_to_tile_4_1_3),
		.out_wire_1_0(vertical_tile_4_1_to_tile_5_1_0),
		.out_wire_1_1(vertical_tile_4_1_to_tile_5_1_1),
		.out_wire_1_2(vertical_tile_4_1_to_tile_5_1_2),
		.out_wire_1_3(vertical_tile_4_1_to_tile_5_1_3),
		.in_wire_1_0(vertical_tile_5_1_to_tile_4_1_0),
		.in_wire_1_1(vertical_tile_5_1_to_tile_4_1_1),
		.in_wire_1_2(vertical_tile_5_1_to_tile_4_1_2),
		.in_wire_1_3(vertical_tile_5_1_to_tile_4_1_3),
		.out_wire_2_0(horizontal_tile_4_1_to_tile_4_0_0),
		.out_wire_2_1(horizontal_tile_4_1_to_tile_4_0_1),
		.out_wire_2_2(horizontal_tile_4_1_to_tile_4_0_2),
		.out_wire_2_3(horizontal_tile_4_1_to_tile_4_0_3),
		.in_wire_2_0(horizontal_tile_4_0_to_tile_4_1_0),
		.in_wire_2_1(horizontal_tile_4_0_to_tile_4_1_1),
		.in_wire_2_2(horizontal_tile_4_0_to_tile_4_1_2),
		.in_wire_2_3(horizontal_tile_4_0_to_tile_4_1_3),
		.out_wire_0_0(horizontal_tile_4_1_to_tile_4_2_0),
		.out_wire_0_1(horizontal_tile_4_1_to_tile_4_2_1),
		.out_wire_0_2(horizontal_tile_4_1_to_tile_4_2_2),
		.out_wire_0_3(horizontal_tile_4_1_to_tile_4_2_3),
		.in_wire_0_0(horizontal_tile_4_2_to_tile_4_1_0),
		.in_wire_0_1(horizontal_tile_4_2_to_tile_4_1_1),
		.in_wire_0_2(horizontal_tile_4_2_to_tile_4_1_2),
		.in_wire_0_3(horizontal_tile_4_2_to_tile_4_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(130)
	);

	pe_tile pe_tile_4_2(
		.out_wire_3_0(vertical_tile_4_2_to_tile_3_2_0),
		.out_wire_3_1(vertical_tile_4_2_to_tile_3_2_1),
		.out_wire_3_2(vertical_tile_4_2_to_tile_3_2_2),
		.out_wire_3_3(vertical_tile_4_2_to_tile_3_2_3),
		.in_wire_3_0(vertical_tile_3_2_to_tile_4_2_0),
		.in_wire_3_1(vertical_tile_3_2_to_tile_4_2_1),
		.in_wire_3_2(vertical_tile_3_2_to_tile_4_2_2),
		.in_wire_3_3(vertical_tile_3_2_to_tile_4_2_3),
		.out_wire_1_0(vertical_tile_4_2_to_tile_5_2_0),
		.out_wire_1_1(vertical_tile_4_2_to_tile_5_2_1),
		.out_wire_1_2(vertical_tile_4_2_to_tile_5_2_2),
		.out_wire_1_3(vertical_tile_4_2_to_tile_5_2_3),
		.in_wire_1_0(vertical_tile_5_2_to_tile_4_2_0),
		.in_wire_1_1(vertical_tile_5_2_to_tile_4_2_1),
		.in_wire_1_2(vertical_tile_5_2_to_tile_4_2_2),
		.in_wire_1_3(vertical_tile_5_2_to_tile_4_2_3),
		.out_wire_2_0(horizontal_tile_4_2_to_tile_4_1_0),
		.out_wire_2_1(horizontal_tile_4_2_to_tile_4_1_1),
		.out_wire_2_2(horizontal_tile_4_2_to_tile_4_1_2),
		.out_wire_2_3(horizontal_tile_4_2_to_tile_4_1_3),
		.in_wire_2_0(horizontal_tile_4_1_to_tile_4_2_0),
		.in_wire_2_1(horizontal_tile_4_1_to_tile_4_2_1),
		.in_wire_2_2(horizontal_tile_4_1_to_tile_4_2_2),
		.in_wire_2_3(horizontal_tile_4_1_to_tile_4_2_3),
		.out_wire_0_0(horizontal_tile_4_2_to_tile_4_3_0),
		.out_wire_0_1(horizontal_tile_4_2_to_tile_4_3_1),
		.out_wire_0_2(horizontal_tile_4_2_to_tile_4_3_2),
		.out_wire_0_3(horizontal_tile_4_2_to_tile_4_3_3),
		.in_wire_0_0(horizontal_tile_4_3_to_tile_4_2_0),
		.in_wire_0_1(horizontal_tile_4_3_to_tile_4_2_1),
		.in_wire_0_2(horizontal_tile_4_3_to_tile_4_2_2),
		.in_wire_0_3(horizontal_tile_4_3_to_tile_4_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(131)
	);

	pe_tile pe_tile_4_3(
		.out_wire_3_0(vertical_tile_4_3_to_tile_3_3_0),
		.out_wire_3_1(vertical_tile_4_3_to_tile_3_3_1),
		.out_wire_3_2(vertical_tile_4_3_to_tile_3_3_2),
		.out_wire_3_3(vertical_tile_4_3_to_tile_3_3_3),
		.in_wire_3_0(vertical_tile_3_3_to_tile_4_3_0),
		.in_wire_3_1(vertical_tile_3_3_to_tile_4_3_1),
		.in_wire_3_2(vertical_tile_3_3_to_tile_4_3_2),
		.in_wire_3_3(vertical_tile_3_3_to_tile_4_3_3),
		.out_wire_1_0(vertical_tile_4_3_to_tile_5_3_0),
		.out_wire_1_1(vertical_tile_4_3_to_tile_5_3_1),
		.out_wire_1_2(vertical_tile_4_3_to_tile_5_3_2),
		.out_wire_1_3(vertical_tile_4_3_to_tile_5_3_3),
		.in_wire_1_0(vertical_tile_5_3_to_tile_4_3_0),
		.in_wire_1_1(vertical_tile_5_3_to_tile_4_3_1),
		.in_wire_1_2(vertical_tile_5_3_to_tile_4_3_2),
		.in_wire_1_3(vertical_tile_5_3_to_tile_4_3_3),
		.out_wire_2_0(horizontal_tile_4_3_to_tile_4_2_0),
		.out_wire_2_1(horizontal_tile_4_3_to_tile_4_2_1),
		.out_wire_2_2(horizontal_tile_4_3_to_tile_4_2_2),
		.out_wire_2_3(horizontal_tile_4_3_to_tile_4_2_3),
		.in_wire_2_0(horizontal_tile_4_2_to_tile_4_3_0),
		.in_wire_2_1(horizontal_tile_4_2_to_tile_4_3_1),
		.in_wire_2_2(horizontal_tile_4_2_to_tile_4_3_2),
		.in_wire_2_3(horizontal_tile_4_2_to_tile_4_3_3),
		.out_wire_0_0(horizontal_tile_4_3_to_tile_4_4_0),
		.out_wire_0_1(horizontal_tile_4_3_to_tile_4_4_1),
		.out_wire_0_2(horizontal_tile_4_3_to_tile_4_4_2),
		.out_wire_0_3(horizontal_tile_4_3_to_tile_4_4_3),
		.in_wire_0_0(horizontal_tile_4_4_to_tile_4_3_0),
		.in_wire_0_1(horizontal_tile_4_4_to_tile_4_3_1),
		.in_wire_0_2(horizontal_tile_4_4_to_tile_4_3_2),
		.in_wire_0_3(horizontal_tile_4_4_to_tile_4_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(132)
	);

	pe_tile pe_tile_4_4(
		.out_wire_3_0(vertical_tile_4_4_to_tile_3_4_0),
		.out_wire_3_1(vertical_tile_4_4_to_tile_3_4_1),
		.out_wire_3_2(vertical_tile_4_4_to_tile_3_4_2),
		.out_wire_3_3(vertical_tile_4_4_to_tile_3_4_3),
		.in_wire_3_0(vertical_tile_3_4_to_tile_4_4_0),
		.in_wire_3_1(vertical_tile_3_4_to_tile_4_4_1),
		.in_wire_3_2(vertical_tile_3_4_to_tile_4_4_2),
		.in_wire_3_3(vertical_tile_3_4_to_tile_4_4_3),
		.out_wire_1_0(vertical_tile_4_4_to_tile_5_4_0),
		.out_wire_1_1(vertical_tile_4_4_to_tile_5_4_1),
		.out_wire_1_2(vertical_tile_4_4_to_tile_5_4_2),
		.out_wire_1_3(vertical_tile_4_4_to_tile_5_4_3),
		.in_wire_1_0(vertical_tile_5_4_to_tile_4_4_0),
		.in_wire_1_1(vertical_tile_5_4_to_tile_4_4_1),
		.in_wire_1_2(vertical_tile_5_4_to_tile_4_4_2),
		.in_wire_1_3(vertical_tile_5_4_to_tile_4_4_3),
		.out_wire_2_0(horizontal_tile_4_4_to_tile_4_3_0),
		.out_wire_2_1(horizontal_tile_4_4_to_tile_4_3_1),
		.out_wire_2_2(horizontal_tile_4_4_to_tile_4_3_2),
		.out_wire_2_3(horizontal_tile_4_4_to_tile_4_3_3),
		.in_wire_2_0(horizontal_tile_4_3_to_tile_4_4_0),
		.in_wire_2_1(horizontal_tile_4_3_to_tile_4_4_1),
		.in_wire_2_2(horizontal_tile_4_3_to_tile_4_4_2),
		.in_wire_2_3(horizontal_tile_4_3_to_tile_4_4_3),
		.out_wire_0_0(horizontal_tile_4_4_to_tile_4_5_0),
		.out_wire_0_1(horizontal_tile_4_4_to_tile_4_5_1),
		.out_wire_0_2(horizontal_tile_4_4_to_tile_4_5_2),
		.out_wire_0_3(horizontal_tile_4_4_to_tile_4_5_3),
		.in_wire_0_0(horizontal_tile_4_5_to_tile_4_4_0),
		.in_wire_0_1(horizontal_tile_4_5_to_tile_4_4_1),
		.in_wire_0_2(horizontal_tile_4_5_to_tile_4_4_2),
		.in_wire_0_3(horizontal_tile_4_5_to_tile_4_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(133)
	);

	pe_tile pe_tile_4_5(
		.out_wire_3_0(vertical_tile_4_5_to_tile_3_5_0),
		.out_wire_3_1(vertical_tile_4_5_to_tile_3_5_1),
		.out_wire_3_2(vertical_tile_4_5_to_tile_3_5_2),
		.out_wire_3_3(vertical_tile_4_5_to_tile_3_5_3),
		.in_wire_3_0(vertical_tile_3_5_to_tile_4_5_0),
		.in_wire_3_1(vertical_tile_3_5_to_tile_4_5_1),
		.in_wire_3_2(vertical_tile_3_5_to_tile_4_5_2),
		.in_wire_3_3(vertical_tile_3_5_to_tile_4_5_3),
		.out_wire_1_0(vertical_tile_4_5_to_tile_5_5_0),
		.out_wire_1_1(vertical_tile_4_5_to_tile_5_5_1),
		.out_wire_1_2(vertical_tile_4_5_to_tile_5_5_2),
		.out_wire_1_3(vertical_tile_4_5_to_tile_5_5_3),
		.in_wire_1_0(vertical_tile_5_5_to_tile_4_5_0),
		.in_wire_1_1(vertical_tile_5_5_to_tile_4_5_1),
		.in_wire_1_2(vertical_tile_5_5_to_tile_4_5_2),
		.in_wire_1_3(vertical_tile_5_5_to_tile_4_5_3),
		.out_wire_2_0(horizontal_tile_4_5_to_tile_4_4_0),
		.out_wire_2_1(horizontal_tile_4_5_to_tile_4_4_1),
		.out_wire_2_2(horizontal_tile_4_5_to_tile_4_4_2),
		.out_wire_2_3(horizontal_tile_4_5_to_tile_4_4_3),
		.in_wire_2_0(horizontal_tile_4_4_to_tile_4_5_0),
		.in_wire_2_1(horizontal_tile_4_4_to_tile_4_5_1),
		.in_wire_2_2(horizontal_tile_4_4_to_tile_4_5_2),
		.in_wire_2_3(horizontal_tile_4_4_to_tile_4_5_3),
		.out_wire_0_0(horizontal_tile_4_5_to_tile_4_6_0),
		.out_wire_0_1(horizontal_tile_4_5_to_tile_4_6_1),
		.out_wire_0_2(horizontal_tile_4_5_to_tile_4_6_2),
		.out_wire_0_3(horizontal_tile_4_5_to_tile_4_6_3),
		.in_wire_0_0(horizontal_tile_4_6_to_tile_4_5_0),
		.in_wire_0_1(horizontal_tile_4_6_to_tile_4_5_1),
		.in_wire_0_2(horizontal_tile_4_6_to_tile_4_5_2),
		.in_wire_0_3(horizontal_tile_4_6_to_tile_4_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(134)
	);

	pe_tile pe_tile_4_6(
		.out_wire_3_0(vertical_tile_4_6_to_tile_3_6_0),
		.out_wire_3_1(vertical_tile_4_6_to_tile_3_6_1),
		.out_wire_3_2(vertical_tile_4_6_to_tile_3_6_2),
		.out_wire_3_3(vertical_tile_4_6_to_tile_3_6_3),
		.in_wire_3_0(vertical_tile_3_6_to_tile_4_6_0),
		.in_wire_3_1(vertical_tile_3_6_to_tile_4_6_1),
		.in_wire_3_2(vertical_tile_3_6_to_tile_4_6_2),
		.in_wire_3_3(vertical_tile_3_6_to_tile_4_6_3),
		.out_wire_1_0(vertical_tile_4_6_to_tile_5_6_0),
		.out_wire_1_1(vertical_tile_4_6_to_tile_5_6_1),
		.out_wire_1_2(vertical_tile_4_6_to_tile_5_6_2),
		.out_wire_1_3(vertical_tile_4_6_to_tile_5_6_3),
		.in_wire_1_0(vertical_tile_5_6_to_tile_4_6_0),
		.in_wire_1_1(vertical_tile_5_6_to_tile_4_6_1),
		.in_wire_1_2(vertical_tile_5_6_to_tile_4_6_2),
		.in_wire_1_3(vertical_tile_5_6_to_tile_4_6_3),
		.out_wire_2_0(horizontal_tile_4_6_to_tile_4_5_0),
		.out_wire_2_1(horizontal_tile_4_6_to_tile_4_5_1),
		.out_wire_2_2(horizontal_tile_4_6_to_tile_4_5_2),
		.out_wire_2_3(horizontal_tile_4_6_to_tile_4_5_3),
		.in_wire_2_0(horizontal_tile_4_5_to_tile_4_6_0),
		.in_wire_2_1(horizontal_tile_4_5_to_tile_4_6_1),
		.in_wire_2_2(horizontal_tile_4_5_to_tile_4_6_2),
		.in_wire_2_3(horizontal_tile_4_5_to_tile_4_6_3),
		.out_wire_0_0(horizontal_tile_4_6_to_tile_4_7_0),
		.out_wire_0_1(horizontal_tile_4_6_to_tile_4_7_1),
		.out_wire_0_2(horizontal_tile_4_6_to_tile_4_7_2),
		.out_wire_0_3(horizontal_tile_4_6_to_tile_4_7_3),
		.in_wire_0_0(horizontal_tile_4_7_to_tile_4_6_0),
		.in_wire_0_1(horizontal_tile_4_7_to_tile_4_6_1),
		.in_wire_0_2(horizontal_tile_4_7_to_tile_4_6_2),
		.in_wire_0_3(horizontal_tile_4_7_to_tile_4_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(135)
	);

	pe_tile pe_tile_4_7(
		.out_wire_3_0(vertical_tile_4_7_to_tile_3_7_0),
		.out_wire_3_1(vertical_tile_4_7_to_tile_3_7_1),
		.out_wire_3_2(vertical_tile_4_7_to_tile_3_7_2),
		.out_wire_3_3(vertical_tile_4_7_to_tile_3_7_3),
		.in_wire_3_0(vertical_tile_3_7_to_tile_4_7_0),
		.in_wire_3_1(vertical_tile_3_7_to_tile_4_7_1),
		.in_wire_3_2(vertical_tile_3_7_to_tile_4_7_2),
		.in_wire_3_3(vertical_tile_3_7_to_tile_4_7_3),
		.out_wire_1_0(vertical_tile_4_7_to_tile_5_7_0),
		.out_wire_1_1(vertical_tile_4_7_to_tile_5_7_1),
		.out_wire_1_2(vertical_tile_4_7_to_tile_5_7_2),
		.out_wire_1_3(vertical_tile_4_7_to_tile_5_7_3),
		.in_wire_1_0(vertical_tile_5_7_to_tile_4_7_0),
		.in_wire_1_1(vertical_tile_5_7_to_tile_4_7_1),
		.in_wire_1_2(vertical_tile_5_7_to_tile_4_7_2),
		.in_wire_1_3(vertical_tile_5_7_to_tile_4_7_3),
		.out_wire_2_0(horizontal_tile_4_7_to_tile_4_6_0),
		.out_wire_2_1(horizontal_tile_4_7_to_tile_4_6_1),
		.out_wire_2_2(horizontal_tile_4_7_to_tile_4_6_2),
		.out_wire_2_3(horizontal_tile_4_7_to_tile_4_6_3),
		.in_wire_2_0(horizontal_tile_4_6_to_tile_4_7_0),
		.in_wire_2_1(horizontal_tile_4_6_to_tile_4_7_1),
		.in_wire_2_2(horizontal_tile_4_6_to_tile_4_7_2),
		.in_wire_2_3(horizontal_tile_4_6_to_tile_4_7_3),
		.out_wire_0_0(horizontal_tile_4_7_to_tile_4_8_0),
		.out_wire_0_1(horizontal_tile_4_7_to_tile_4_8_1),
		.out_wire_0_2(horizontal_tile_4_7_to_tile_4_8_2),
		.out_wire_0_3(horizontal_tile_4_7_to_tile_4_8_3),
		.in_wire_0_0(horizontal_tile_4_8_to_tile_4_7_0),
		.in_wire_0_1(horizontal_tile_4_8_to_tile_4_7_1),
		.in_wire_0_2(horizontal_tile_4_8_to_tile_4_7_2),
		.in_wire_0_3(horizontal_tile_4_8_to_tile_4_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(136)
	);

	pe_tile pe_tile_4_8(
		.out_wire_3_0(vertical_tile_4_8_to_tile_3_8_0),
		.out_wire_3_1(vertical_tile_4_8_to_tile_3_8_1),
		.out_wire_3_2(vertical_tile_4_8_to_tile_3_8_2),
		.out_wire_3_3(vertical_tile_4_8_to_tile_3_8_3),
		.in_wire_3_0(vertical_tile_3_8_to_tile_4_8_0),
		.in_wire_3_1(vertical_tile_3_8_to_tile_4_8_1),
		.in_wire_3_2(vertical_tile_3_8_to_tile_4_8_2),
		.in_wire_3_3(vertical_tile_3_8_to_tile_4_8_3),
		.out_wire_1_0(vertical_tile_4_8_to_tile_5_8_0),
		.out_wire_1_1(vertical_tile_4_8_to_tile_5_8_1),
		.out_wire_1_2(vertical_tile_4_8_to_tile_5_8_2),
		.out_wire_1_3(vertical_tile_4_8_to_tile_5_8_3),
		.in_wire_1_0(vertical_tile_5_8_to_tile_4_8_0),
		.in_wire_1_1(vertical_tile_5_8_to_tile_4_8_1),
		.in_wire_1_2(vertical_tile_5_8_to_tile_4_8_2),
		.in_wire_1_3(vertical_tile_5_8_to_tile_4_8_3),
		.out_wire_2_0(horizontal_tile_4_8_to_tile_4_7_0),
		.out_wire_2_1(horizontal_tile_4_8_to_tile_4_7_1),
		.out_wire_2_2(horizontal_tile_4_8_to_tile_4_7_2),
		.out_wire_2_3(horizontal_tile_4_8_to_tile_4_7_3),
		.in_wire_2_0(horizontal_tile_4_7_to_tile_4_8_0),
		.in_wire_2_1(horizontal_tile_4_7_to_tile_4_8_1),
		.in_wire_2_2(horizontal_tile_4_7_to_tile_4_8_2),
		.in_wire_2_3(horizontal_tile_4_7_to_tile_4_8_3),
		.out_wire_0_0(horizontal_tile_4_8_to_tile_4_9_0),
		.out_wire_0_1(horizontal_tile_4_8_to_tile_4_9_1),
		.out_wire_0_2(horizontal_tile_4_8_to_tile_4_9_2),
		.out_wire_0_3(horizontal_tile_4_8_to_tile_4_9_3),
		.in_wire_0_0(horizontal_tile_4_9_to_tile_4_8_0),
		.in_wire_0_1(horizontal_tile_4_9_to_tile_4_8_1),
		.in_wire_0_2(horizontal_tile_4_9_to_tile_4_8_2),
		.in_wire_0_3(horizontal_tile_4_9_to_tile_4_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(137)
	);

	pe_tile pe_tile_4_9(
		.out_wire_3_0(vertical_tile_4_9_to_tile_3_9_0),
		.out_wire_3_1(vertical_tile_4_9_to_tile_3_9_1),
		.out_wire_3_2(vertical_tile_4_9_to_tile_3_9_2),
		.out_wire_3_3(vertical_tile_4_9_to_tile_3_9_3),
		.in_wire_3_0(vertical_tile_3_9_to_tile_4_9_0),
		.in_wire_3_1(vertical_tile_3_9_to_tile_4_9_1),
		.in_wire_3_2(vertical_tile_3_9_to_tile_4_9_2),
		.in_wire_3_3(vertical_tile_3_9_to_tile_4_9_3),
		.out_wire_1_0(vertical_tile_4_9_to_tile_5_9_0),
		.out_wire_1_1(vertical_tile_4_9_to_tile_5_9_1),
		.out_wire_1_2(vertical_tile_4_9_to_tile_5_9_2),
		.out_wire_1_3(vertical_tile_4_9_to_tile_5_9_3),
		.in_wire_1_0(vertical_tile_5_9_to_tile_4_9_0),
		.in_wire_1_1(vertical_tile_5_9_to_tile_4_9_1),
		.in_wire_1_2(vertical_tile_5_9_to_tile_4_9_2),
		.in_wire_1_3(vertical_tile_5_9_to_tile_4_9_3),
		.out_wire_2_0(horizontal_tile_4_9_to_tile_4_8_0),
		.out_wire_2_1(horizontal_tile_4_9_to_tile_4_8_1),
		.out_wire_2_2(horizontal_tile_4_9_to_tile_4_8_2),
		.out_wire_2_3(horizontal_tile_4_9_to_tile_4_8_3),
		.in_wire_2_0(horizontal_tile_4_8_to_tile_4_9_0),
		.in_wire_2_1(horizontal_tile_4_8_to_tile_4_9_1),
		.in_wire_2_2(horizontal_tile_4_8_to_tile_4_9_2),
		.in_wire_2_3(horizontal_tile_4_8_to_tile_4_9_3),
		.out_wire_0_0(horizontal_tile_4_9_to_tile_4_10_0),
		.out_wire_0_1(horizontal_tile_4_9_to_tile_4_10_1),
		.out_wire_0_2(horizontal_tile_4_9_to_tile_4_10_2),
		.out_wire_0_3(horizontal_tile_4_9_to_tile_4_10_3),
		.in_wire_0_0(horizontal_tile_4_10_to_tile_4_9_0),
		.in_wire_0_1(horizontal_tile_4_10_to_tile_4_9_1),
		.in_wire_0_2(horizontal_tile_4_10_to_tile_4_9_2),
		.in_wire_0_3(horizontal_tile_4_10_to_tile_4_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(138)
	);

	pe_tile pe_tile_4_10(
		.out_wire_3_0(vertical_tile_4_10_to_tile_3_10_0),
		.out_wire_3_1(vertical_tile_4_10_to_tile_3_10_1),
		.out_wire_3_2(vertical_tile_4_10_to_tile_3_10_2),
		.out_wire_3_3(vertical_tile_4_10_to_tile_3_10_3),
		.in_wire_3_0(vertical_tile_3_10_to_tile_4_10_0),
		.in_wire_3_1(vertical_tile_3_10_to_tile_4_10_1),
		.in_wire_3_2(vertical_tile_3_10_to_tile_4_10_2),
		.in_wire_3_3(vertical_tile_3_10_to_tile_4_10_3),
		.out_wire_1_0(vertical_tile_4_10_to_tile_5_10_0),
		.out_wire_1_1(vertical_tile_4_10_to_tile_5_10_1),
		.out_wire_1_2(vertical_tile_4_10_to_tile_5_10_2),
		.out_wire_1_3(vertical_tile_4_10_to_tile_5_10_3),
		.in_wire_1_0(vertical_tile_5_10_to_tile_4_10_0),
		.in_wire_1_1(vertical_tile_5_10_to_tile_4_10_1),
		.in_wire_1_2(vertical_tile_5_10_to_tile_4_10_2),
		.in_wire_1_3(vertical_tile_5_10_to_tile_4_10_3),
		.out_wire_2_0(horizontal_tile_4_10_to_tile_4_9_0),
		.out_wire_2_1(horizontal_tile_4_10_to_tile_4_9_1),
		.out_wire_2_2(horizontal_tile_4_10_to_tile_4_9_2),
		.out_wire_2_3(horizontal_tile_4_10_to_tile_4_9_3),
		.in_wire_2_0(horizontal_tile_4_9_to_tile_4_10_0),
		.in_wire_2_1(horizontal_tile_4_9_to_tile_4_10_1),
		.in_wire_2_2(horizontal_tile_4_9_to_tile_4_10_2),
		.in_wire_2_3(horizontal_tile_4_9_to_tile_4_10_3),
		.out_wire_0_0(horizontal_tile_4_10_to_tile_4_11_0),
		.out_wire_0_1(horizontal_tile_4_10_to_tile_4_11_1),
		.out_wire_0_2(horizontal_tile_4_10_to_tile_4_11_2),
		.out_wire_0_3(horizontal_tile_4_10_to_tile_4_11_3),
		.in_wire_0_0(horizontal_tile_4_11_to_tile_4_10_0),
		.in_wire_0_1(horizontal_tile_4_11_to_tile_4_10_1),
		.in_wire_0_2(horizontal_tile_4_11_to_tile_4_10_2),
		.in_wire_0_3(horizontal_tile_4_11_to_tile_4_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(139)
	);

	pe_tile pe_tile_4_11(
		.out_wire_3_0(vertical_tile_4_11_to_tile_3_11_0),
		.out_wire_3_1(vertical_tile_4_11_to_tile_3_11_1),
		.out_wire_3_2(vertical_tile_4_11_to_tile_3_11_2),
		.out_wire_3_3(vertical_tile_4_11_to_tile_3_11_3),
		.in_wire_3_0(vertical_tile_3_11_to_tile_4_11_0),
		.in_wire_3_1(vertical_tile_3_11_to_tile_4_11_1),
		.in_wire_3_2(vertical_tile_3_11_to_tile_4_11_2),
		.in_wire_3_3(vertical_tile_3_11_to_tile_4_11_3),
		.out_wire_1_0(vertical_tile_4_11_to_tile_5_11_0),
		.out_wire_1_1(vertical_tile_4_11_to_tile_5_11_1),
		.out_wire_1_2(vertical_tile_4_11_to_tile_5_11_2),
		.out_wire_1_3(vertical_tile_4_11_to_tile_5_11_3),
		.in_wire_1_0(vertical_tile_5_11_to_tile_4_11_0),
		.in_wire_1_1(vertical_tile_5_11_to_tile_4_11_1),
		.in_wire_1_2(vertical_tile_5_11_to_tile_4_11_2),
		.in_wire_1_3(vertical_tile_5_11_to_tile_4_11_3),
		.out_wire_2_0(horizontal_tile_4_11_to_tile_4_10_0),
		.out_wire_2_1(horizontal_tile_4_11_to_tile_4_10_1),
		.out_wire_2_2(horizontal_tile_4_11_to_tile_4_10_2),
		.out_wire_2_3(horizontal_tile_4_11_to_tile_4_10_3),
		.in_wire_2_0(horizontal_tile_4_10_to_tile_4_11_0),
		.in_wire_2_1(horizontal_tile_4_10_to_tile_4_11_1),
		.in_wire_2_2(horizontal_tile_4_10_to_tile_4_11_2),
		.in_wire_2_3(horizontal_tile_4_10_to_tile_4_11_3),
		.out_wire_0_0(horizontal_tile_4_11_to_tile_4_12_0),
		.out_wire_0_1(horizontal_tile_4_11_to_tile_4_12_1),
		.out_wire_0_2(horizontal_tile_4_11_to_tile_4_12_2),
		.out_wire_0_3(horizontal_tile_4_11_to_tile_4_12_3),
		.in_wire_0_0(horizontal_tile_4_12_to_tile_4_11_0),
		.in_wire_0_1(horizontal_tile_4_12_to_tile_4_11_1),
		.in_wire_0_2(horizontal_tile_4_12_to_tile_4_11_2),
		.in_wire_0_3(horizontal_tile_4_12_to_tile_4_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(140)
	);

	pe_tile pe_tile_4_12(
		.out_wire_3_0(vertical_tile_4_12_to_tile_3_12_0),
		.out_wire_3_1(vertical_tile_4_12_to_tile_3_12_1),
		.out_wire_3_2(vertical_tile_4_12_to_tile_3_12_2),
		.out_wire_3_3(vertical_tile_4_12_to_tile_3_12_3),
		.in_wire_3_0(vertical_tile_3_12_to_tile_4_12_0),
		.in_wire_3_1(vertical_tile_3_12_to_tile_4_12_1),
		.in_wire_3_2(vertical_tile_3_12_to_tile_4_12_2),
		.in_wire_3_3(vertical_tile_3_12_to_tile_4_12_3),
		.out_wire_1_0(vertical_tile_4_12_to_tile_5_12_0),
		.out_wire_1_1(vertical_tile_4_12_to_tile_5_12_1),
		.out_wire_1_2(vertical_tile_4_12_to_tile_5_12_2),
		.out_wire_1_3(vertical_tile_4_12_to_tile_5_12_3),
		.in_wire_1_0(vertical_tile_5_12_to_tile_4_12_0),
		.in_wire_1_1(vertical_tile_5_12_to_tile_4_12_1),
		.in_wire_1_2(vertical_tile_5_12_to_tile_4_12_2),
		.in_wire_1_3(vertical_tile_5_12_to_tile_4_12_3),
		.out_wire_2_0(horizontal_tile_4_12_to_tile_4_11_0),
		.out_wire_2_1(horizontal_tile_4_12_to_tile_4_11_1),
		.out_wire_2_2(horizontal_tile_4_12_to_tile_4_11_2),
		.out_wire_2_3(horizontal_tile_4_12_to_tile_4_11_3),
		.in_wire_2_0(horizontal_tile_4_11_to_tile_4_12_0),
		.in_wire_2_1(horizontal_tile_4_11_to_tile_4_12_1),
		.in_wire_2_2(horizontal_tile_4_11_to_tile_4_12_2),
		.in_wire_2_3(horizontal_tile_4_11_to_tile_4_12_3),
		.out_wire_0_0(horizontal_tile_4_12_to_tile_4_13_0),
		.out_wire_0_1(horizontal_tile_4_12_to_tile_4_13_1),
		.out_wire_0_2(horizontal_tile_4_12_to_tile_4_13_2),
		.out_wire_0_3(horizontal_tile_4_12_to_tile_4_13_3),
		.in_wire_0_0(horizontal_tile_4_13_to_tile_4_12_0),
		.in_wire_0_1(horizontal_tile_4_13_to_tile_4_12_1),
		.in_wire_0_2(horizontal_tile_4_13_to_tile_4_12_2),
		.in_wire_0_3(horizontal_tile_4_13_to_tile_4_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(141)
	);

	pe_tile pe_tile_4_13(
		.out_wire_3_0(vertical_tile_4_13_to_tile_3_13_0),
		.out_wire_3_1(vertical_tile_4_13_to_tile_3_13_1),
		.out_wire_3_2(vertical_tile_4_13_to_tile_3_13_2),
		.out_wire_3_3(vertical_tile_4_13_to_tile_3_13_3),
		.in_wire_3_0(vertical_tile_3_13_to_tile_4_13_0),
		.in_wire_3_1(vertical_tile_3_13_to_tile_4_13_1),
		.in_wire_3_2(vertical_tile_3_13_to_tile_4_13_2),
		.in_wire_3_3(vertical_tile_3_13_to_tile_4_13_3),
		.out_wire_1_0(vertical_tile_4_13_to_tile_5_13_0),
		.out_wire_1_1(vertical_tile_4_13_to_tile_5_13_1),
		.out_wire_1_2(vertical_tile_4_13_to_tile_5_13_2),
		.out_wire_1_3(vertical_tile_4_13_to_tile_5_13_3),
		.in_wire_1_0(vertical_tile_5_13_to_tile_4_13_0),
		.in_wire_1_1(vertical_tile_5_13_to_tile_4_13_1),
		.in_wire_1_2(vertical_tile_5_13_to_tile_4_13_2),
		.in_wire_1_3(vertical_tile_5_13_to_tile_4_13_3),
		.out_wire_2_0(horizontal_tile_4_13_to_tile_4_12_0),
		.out_wire_2_1(horizontal_tile_4_13_to_tile_4_12_1),
		.out_wire_2_2(horizontal_tile_4_13_to_tile_4_12_2),
		.out_wire_2_3(horizontal_tile_4_13_to_tile_4_12_3),
		.in_wire_2_0(horizontal_tile_4_12_to_tile_4_13_0),
		.in_wire_2_1(horizontal_tile_4_12_to_tile_4_13_1),
		.in_wire_2_2(horizontal_tile_4_12_to_tile_4_13_2),
		.in_wire_2_3(horizontal_tile_4_12_to_tile_4_13_3),
		.out_wire_0_0(horizontal_tile_4_13_to_tile_4_14_0),
		.out_wire_0_1(horizontal_tile_4_13_to_tile_4_14_1),
		.out_wire_0_2(horizontal_tile_4_13_to_tile_4_14_2),
		.out_wire_0_3(horizontal_tile_4_13_to_tile_4_14_3),
		.in_wire_0_0(horizontal_tile_4_14_to_tile_4_13_0),
		.in_wire_0_1(horizontal_tile_4_14_to_tile_4_13_1),
		.in_wire_0_2(horizontal_tile_4_14_to_tile_4_13_2),
		.in_wire_0_3(horizontal_tile_4_14_to_tile_4_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(142)
	);

	pe_tile pe_tile_4_14(
		.out_wire_3_0(vertical_tile_4_14_to_tile_3_14_0),
		.out_wire_3_1(vertical_tile_4_14_to_tile_3_14_1),
		.out_wire_3_2(vertical_tile_4_14_to_tile_3_14_2),
		.out_wire_3_3(vertical_tile_4_14_to_tile_3_14_3),
		.in_wire_3_0(vertical_tile_3_14_to_tile_4_14_0),
		.in_wire_3_1(vertical_tile_3_14_to_tile_4_14_1),
		.in_wire_3_2(vertical_tile_3_14_to_tile_4_14_2),
		.in_wire_3_3(vertical_tile_3_14_to_tile_4_14_3),
		.out_wire_1_0(vertical_tile_4_14_to_tile_5_14_0),
		.out_wire_1_1(vertical_tile_4_14_to_tile_5_14_1),
		.out_wire_1_2(vertical_tile_4_14_to_tile_5_14_2),
		.out_wire_1_3(vertical_tile_4_14_to_tile_5_14_3),
		.in_wire_1_0(vertical_tile_5_14_to_tile_4_14_0),
		.in_wire_1_1(vertical_tile_5_14_to_tile_4_14_1),
		.in_wire_1_2(vertical_tile_5_14_to_tile_4_14_2),
		.in_wire_1_3(vertical_tile_5_14_to_tile_4_14_3),
		.out_wire_2_0(horizontal_tile_4_14_to_tile_4_13_0),
		.out_wire_2_1(horizontal_tile_4_14_to_tile_4_13_1),
		.out_wire_2_2(horizontal_tile_4_14_to_tile_4_13_2),
		.out_wire_2_3(horizontal_tile_4_14_to_tile_4_13_3),
		.in_wire_2_0(horizontal_tile_4_13_to_tile_4_14_0),
		.in_wire_2_1(horizontal_tile_4_13_to_tile_4_14_1),
		.in_wire_2_2(horizontal_tile_4_13_to_tile_4_14_2),
		.in_wire_2_3(horizontal_tile_4_13_to_tile_4_14_3),
		.out_wire_0_0(horizontal_tile_4_14_to_tile_4_15_0),
		.out_wire_0_1(horizontal_tile_4_14_to_tile_4_15_1),
		.out_wire_0_2(horizontal_tile_4_14_to_tile_4_15_2),
		.out_wire_0_3(horizontal_tile_4_14_to_tile_4_15_3),
		.in_wire_0_0(horizontal_tile_4_15_to_tile_4_14_0),
		.in_wire_0_1(horizontal_tile_4_15_to_tile_4_14_1),
		.in_wire_0_2(horizontal_tile_4_15_to_tile_4_14_2),
		.in_wire_0_3(horizontal_tile_4_15_to_tile_4_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(143)
	);

	pe_tile pe_tile_4_15(
		.out_wire_3_0(vertical_tile_4_15_to_tile_3_15_0),
		.out_wire_3_1(vertical_tile_4_15_to_tile_3_15_1),
		.out_wire_3_2(vertical_tile_4_15_to_tile_3_15_2),
		.out_wire_3_3(vertical_tile_4_15_to_tile_3_15_3),
		.in_wire_3_0(vertical_tile_3_15_to_tile_4_15_0),
		.in_wire_3_1(vertical_tile_3_15_to_tile_4_15_1),
		.in_wire_3_2(vertical_tile_3_15_to_tile_4_15_2),
		.in_wire_3_3(vertical_tile_3_15_to_tile_4_15_3),
		.out_wire_1_0(vertical_tile_4_15_to_tile_5_15_0),
		.out_wire_1_1(vertical_tile_4_15_to_tile_5_15_1),
		.out_wire_1_2(vertical_tile_4_15_to_tile_5_15_2),
		.out_wire_1_3(vertical_tile_4_15_to_tile_5_15_3),
		.in_wire_1_0(vertical_tile_5_15_to_tile_4_15_0),
		.in_wire_1_1(vertical_tile_5_15_to_tile_4_15_1),
		.in_wire_1_2(vertical_tile_5_15_to_tile_4_15_2),
		.in_wire_1_3(vertical_tile_5_15_to_tile_4_15_3),
		.out_wire_2_0(horizontal_tile_4_15_to_tile_4_14_0),
		.out_wire_2_1(horizontal_tile_4_15_to_tile_4_14_1),
		.out_wire_2_2(horizontal_tile_4_15_to_tile_4_14_2),
		.out_wire_2_3(horizontal_tile_4_15_to_tile_4_14_3),
		.in_wire_2_0(horizontal_tile_4_14_to_tile_4_15_0),
		.in_wire_2_1(horizontal_tile_4_14_to_tile_4_15_1),
		.in_wire_2_2(horizontal_tile_4_14_to_tile_4_15_2),
		.in_wire_2_3(horizontal_tile_4_14_to_tile_4_15_3),
		.out_wire_0_0(horizontal_tile_4_15_to_tile_4_16_0),
		.out_wire_0_1(horizontal_tile_4_15_to_tile_4_16_1),
		.out_wire_0_2(horizontal_tile_4_15_to_tile_4_16_2),
		.out_wire_0_3(horizontal_tile_4_15_to_tile_4_16_3),
		.in_wire_0_0(horizontal_tile_4_16_to_tile_4_15_0),
		.in_wire_0_1(horizontal_tile_4_16_to_tile_4_15_1),
		.in_wire_0_2(horizontal_tile_4_16_to_tile_4_15_2),
		.in_wire_0_3(horizontal_tile_4_16_to_tile_4_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(144)
	);

	pe_tile pe_tile_4_16(
		.out_wire_3_0(vertical_tile_4_16_to_tile_3_16_0),
		.out_wire_3_1(vertical_tile_4_16_to_tile_3_16_1),
		.out_wire_3_2(vertical_tile_4_16_to_tile_3_16_2),
		.out_wire_3_3(vertical_tile_4_16_to_tile_3_16_3),
		.in_wire_3_0(vertical_tile_3_16_to_tile_4_16_0),
		.in_wire_3_1(vertical_tile_3_16_to_tile_4_16_1),
		.in_wire_3_2(vertical_tile_3_16_to_tile_4_16_2),
		.in_wire_3_3(vertical_tile_3_16_to_tile_4_16_3),
		.out_wire_1_0(vertical_tile_4_16_to_tile_5_16_0),
		.out_wire_1_1(vertical_tile_4_16_to_tile_5_16_1),
		.out_wire_1_2(vertical_tile_4_16_to_tile_5_16_2),
		.out_wire_1_3(vertical_tile_4_16_to_tile_5_16_3),
		.in_wire_1_0(vertical_tile_5_16_to_tile_4_16_0),
		.in_wire_1_1(vertical_tile_5_16_to_tile_4_16_1),
		.in_wire_1_2(vertical_tile_5_16_to_tile_4_16_2),
		.in_wire_1_3(vertical_tile_5_16_to_tile_4_16_3),
		.out_wire_2_0(horizontal_tile_4_16_to_tile_4_15_0),
		.out_wire_2_1(horizontal_tile_4_16_to_tile_4_15_1),
		.out_wire_2_2(horizontal_tile_4_16_to_tile_4_15_2),
		.out_wire_2_3(horizontal_tile_4_16_to_tile_4_15_3),
		.in_wire_2_0(horizontal_tile_4_15_to_tile_4_16_0),
		.in_wire_2_1(horizontal_tile_4_15_to_tile_4_16_1),
		.in_wire_2_2(horizontal_tile_4_15_to_tile_4_16_2),
		.in_wire_2_3(horizontal_tile_4_15_to_tile_4_16_3),
		.out_wire_0_0(horizontal_tile_4_16_to_tile_4_17_0),
		.out_wire_0_1(horizontal_tile_4_16_to_tile_4_17_1),
		.out_wire_0_2(horizontal_tile_4_16_to_tile_4_17_2),
		.out_wire_0_3(horizontal_tile_4_16_to_tile_4_17_3),
		.in_wire_0_0(horizontal_tile_4_17_to_tile_4_16_0),
		.in_wire_0_1(horizontal_tile_4_17_to_tile_4_16_1),
		.in_wire_0_2(horizontal_tile_4_17_to_tile_4_16_2),
		.in_wire_0_3(horizontal_tile_4_17_to_tile_4_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(145)
	);

	pe_tile pe_tile_4_17(
		.out_wire_3_0(vertical_tile_4_17_to_tile_3_17_0),
		.out_wire_3_1(vertical_tile_4_17_to_tile_3_17_1),
		.out_wire_3_2(vertical_tile_4_17_to_tile_3_17_2),
		.out_wire_3_3(vertical_tile_4_17_to_tile_3_17_3),
		.in_wire_3_0(vertical_tile_3_17_to_tile_4_17_0),
		.in_wire_3_1(vertical_tile_3_17_to_tile_4_17_1),
		.in_wire_3_2(vertical_tile_3_17_to_tile_4_17_2),
		.in_wire_3_3(vertical_tile_3_17_to_tile_4_17_3),
		.out_wire_1_0(vertical_tile_4_17_to_tile_5_17_0),
		.out_wire_1_1(vertical_tile_4_17_to_tile_5_17_1),
		.out_wire_1_2(vertical_tile_4_17_to_tile_5_17_2),
		.out_wire_1_3(vertical_tile_4_17_to_tile_5_17_3),
		.in_wire_1_0(vertical_tile_5_17_to_tile_4_17_0),
		.in_wire_1_1(vertical_tile_5_17_to_tile_4_17_1),
		.in_wire_1_2(vertical_tile_5_17_to_tile_4_17_2),
		.in_wire_1_3(vertical_tile_5_17_to_tile_4_17_3),
		.out_wire_2_0(horizontal_tile_4_17_to_tile_4_16_0),
		.out_wire_2_1(horizontal_tile_4_17_to_tile_4_16_1),
		.out_wire_2_2(horizontal_tile_4_17_to_tile_4_16_2),
		.out_wire_2_3(horizontal_tile_4_17_to_tile_4_16_3),
		.in_wire_2_0(horizontal_tile_4_16_to_tile_4_17_0),
		.in_wire_2_1(horizontal_tile_4_16_to_tile_4_17_1),
		.in_wire_2_2(horizontal_tile_4_16_to_tile_4_17_2),
		.in_wire_2_3(horizontal_tile_4_16_to_tile_4_17_3),
		.out_wire_0_0(horizontal_tile_4_17_to_tile_4_18_0),
		.out_wire_0_1(horizontal_tile_4_17_to_tile_4_18_1),
		.out_wire_0_2(horizontal_tile_4_17_to_tile_4_18_2),
		.out_wire_0_3(horizontal_tile_4_17_to_tile_4_18_3),
		.in_wire_0_0(horizontal_tile_4_18_to_tile_4_17_0),
		.in_wire_0_1(horizontal_tile_4_18_to_tile_4_17_1),
		.in_wire_0_2(horizontal_tile_4_18_to_tile_4_17_2),
		.in_wire_0_3(horizontal_tile_4_18_to_tile_4_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(146)
	);

	pe_tile pe_tile_4_18(
		.out_wire_3_0(vertical_tile_4_18_to_tile_3_18_0),
		.out_wire_3_1(vertical_tile_4_18_to_tile_3_18_1),
		.out_wire_3_2(vertical_tile_4_18_to_tile_3_18_2),
		.out_wire_3_3(vertical_tile_4_18_to_tile_3_18_3),
		.in_wire_3_0(vertical_tile_3_18_to_tile_4_18_0),
		.in_wire_3_1(vertical_tile_3_18_to_tile_4_18_1),
		.in_wire_3_2(vertical_tile_3_18_to_tile_4_18_2),
		.in_wire_3_3(vertical_tile_3_18_to_tile_4_18_3),
		.out_wire_1_0(vertical_tile_4_18_to_tile_5_18_0),
		.out_wire_1_1(vertical_tile_4_18_to_tile_5_18_1),
		.out_wire_1_2(vertical_tile_4_18_to_tile_5_18_2),
		.out_wire_1_3(vertical_tile_4_18_to_tile_5_18_3),
		.in_wire_1_0(vertical_tile_5_18_to_tile_4_18_0),
		.in_wire_1_1(vertical_tile_5_18_to_tile_4_18_1),
		.in_wire_1_2(vertical_tile_5_18_to_tile_4_18_2),
		.in_wire_1_3(vertical_tile_5_18_to_tile_4_18_3),
		.out_wire_2_0(horizontal_tile_4_18_to_tile_4_17_0),
		.out_wire_2_1(horizontal_tile_4_18_to_tile_4_17_1),
		.out_wire_2_2(horizontal_tile_4_18_to_tile_4_17_2),
		.out_wire_2_3(horizontal_tile_4_18_to_tile_4_17_3),
		.in_wire_2_0(horizontal_tile_4_17_to_tile_4_18_0),
		.in_wire_2_1(horizontal_tile_4_17_to_tile_4_18_1),
		.in_wire_2_2(horizontal_tile_4_17_to_tile_4_18_2),
		.in_wire_2_3(horizontal_tile_4_17_to_tile_4_18_3),
		.out_wire_0_0(horizontal_tile_4_18_to_tile_4_19_0),
		.out_wire_0_1(horizontal_tile_4_18_to_tile_4_19_1),
		.out_wire_0_2(horizontal_tile_4_18_to_tile_4_19_2),
		.out_wire_0_3(horizontal_tile_4_18_to_tile_4_19_3),
		.in_wire_0_0(horizontal_tile_4_19_to_tile_4_18_0),
		.in_wire_0_1(horizontal_tile_4_19_to_tile_4_18_1),
		.in_wire_0_2(horizontal_tile_4_19_to_tile_4_18_2),
		.in_wire_0_3(horizontal_tile_4_19_to_tile_4_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(147)
	);

	pe_tile pe_tile_4_19(
		.out_wire_3_0(vertical_tile_4_19_to_tile_3_19_0),
		.out_wire_3_1(vertical_tile_4_19_to_tile_3_19_1),
		.out_wire_3_2(vertical_tile_4_19_to_tile_3_19_2),
		.out_wire_3_3(vertical_tile_4_19_to_tile_3_19_3),
		.in_wire_3_0(vertical_tile_3_19_to_tile_4_19_0),
		.in_wire_3_1(vertical_tile_3_19_to_tile_4_19_1),
		.in_wire_3_2(vertical_tile_3_19_to_tile_4_19_2),
		.in_wire_3_3(vertical_tile_3_19_to_tile_4_19_3),
		.out_wire_1_0(vertical_tile_4_19_to_tile_5_19_0),
		.out_wire_1_1(vertical_tile_4_19_to_tile_5_19_1),
		.out_wire_1_2(vertical_tile_4_19_to_tile_5_19_2),
		.out_wire_1_3(vertical_tile_4_19_to_tile_5_19_3),
		.in_wire_1_0(vertical_tile_5_19_to_tile_4_19_0),
		.in_wire_1_1(vertical_tile_5_19_to_tile_4_19_1),
		.in_wire_1_2(vertical_tile_5_19_to_tile_4_19_2),
		.in_wire_1_3(vertical_tile_5_19_to_tile_4_19_3),
		.out_wire_2_0(horizontal_tile_4_19_to_tile_4_18_0),
		.out_wire_2_1(horizontal_tile_4_19_to_tile_4_18_1),
		.out_wire_2_2(horizontal_tile_4_19_to_tile_4_18_2),
		.out_wire_2_3(horizontal_tile_4_19_to_tile_4_18_3),
		.in_wire_2_0(horizontal_tile_4_18_to_tile_4_19_0),
		.in_wire_2_1(horizontal_tile_4_18_to_tile_4_19_1),
		.in_wire_2_2(horizontal_tile_4_18_to_tile_4_19_2),
		.in_wire_2_3(horizontal_tile_4_18_to_tile_4_19_3),
		.out_wire_0_0(horizontal_tile_4_19_to_tile_4_20_0),
		.out_wire_0_1(horizontal_tile_4_19_to_tile_4_20_1),
		.out_wire_0_2(horizontal_tile_4_19_to_tile_4_20_2),
		.out_wire_0_3(horizontal_tile_4_19_to_tile_4_20_3),
		.in_wire_0_0(horizontal_tile_4_20_to_tile_4_19_0),
		.in_wire_0_1(horizontal_tile_4_20_to_tile_4_19_1),
		.in_wire_0_2(horizontal_tile_4_20_to_tile_4_19_2),
		.in_wire_0_3(horizontal_tile_4_20_to_tile_4_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(148)
	);

	pe_tile pe_tile_4_20(
		.out_wire_3_0(vertical_tile_4_20_to_tile_3_20_0),
		.out_wire_3_1(vertical_tile_4_20_to_tile_3_20_1),
		.out_wire_3_2(vertical_tile_4_20_to_tile_3_20_2),
		.out_wire_3_3(vertical_tile_4_20_to_tile_3_20_3),
		.in_wire_3_0(vertical_tile_3_20_to_tile_4_20_0),
		.in_wire_3_1(vertical_tile_3_20_to_tile_4_20_1),
		.in_wire_3_2(vertical_tile_3_20_to_tile_4_20_2),
		.in_wire_3_3(vertical_tile_3_20_to_tile_4_20_3),
		.out_wire_1_0(vertical_tile_4_20_to_tile_5_20_0),
		.out_wire_1_1(vertical_tile_4_20_to_tile_5_20_1),
		.out_wire_1_2(vertical_tile_4_20_to_tile_5_20_2),
		.out_wire_1_3(vertical_tile_4_20_to_tile_5_20_3),
		.in_wire_1_0(vertical_tile_5_20_to_tile_4_20_0),
		.in_wire_1_1(vertical_tile_5_20_to_tile_4_20_1),
		.in_wire_1_2(vertical_tile_5_20_to_tile_4_20_2),
		.in_wire_1_3(vertical_tile_5_20_to_tile_4_20_3),
		.out_wire_2_0(horizontal_tile_4_20_to_tile_4_19_0),
		.out_wire_2_1(horizontal_tile_4_20_to_tile_4_19_1),
		.out_wire_2_2(horizontal_tile_4_20_to_tile_4_19_2),
		.out_wire_2_3(horizontal_tile_4_20_to_tile_4_19_3),
		.in_wire_2_0(horizontal_tile_4_19_to_tile_4_20_0),
		.in_wire_2_1(horizontal_tile_4_19_to_tile_4_20_1),
		.in_wire_2_2(horizontal_tile_4_19_to_tile_4_20_2),
		.in_wire_2_3(horizontal_tile_4_19_to_tile_4_20_3),
		.out_wire_0_0(horizontal_tile_4_20_to_tile_4_21_0),
		.out_wire_0_1(horizontal_tile_4_20_to_tile_4_21_1),
		.out_wire_0_2(horizontal_tile_4_20_to_tile_4_21_2),
		.out_wire_0_3(horizontal_tile_4_20_to_tile_4_21_3),
		.in_wire_0_0(horizontal_tile_4_21_to_tile_4_20_0),
		.in_wire_0_1(horizontal_tile_4_21_to_tile_4_20_1),
		.in_wire_0_2(horizontal_tile_4_21_to_tile_4_20_2),
		.in_wire_0_3(horizontal_tile_4_21_to_tile_4_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(149)
	);

	pe_tile pe_tile_4_21(
		.out_wire_3_0(vertical_tile_4_21_to_tile_3_21_0),
		.out_wire_3_1(vertical_tile_4_21_to_tile_3_21_1),
		.out_wire_3_2(vertical_tile_4_21_to_tile_3_21_2),
		.out_wire_3_3(vertical_tile_4_21_to_tile_3_21_3),
		.in_wire_3_0(vertical_tile_3_21_to_tile_4_21_0),
		.in_wire_3_1(vertical_tile_3_21_to_tile_4_21_1),
		.in_wire_3_2(vertical_tile_3_21_to_tile_4_21_2),
		.in_wire_3_3(vertical_tile_3_21_to_tile_4_21_3),
		.out_wire_1_0(vertical_tile_4_21_to_tile_5_21_0),
		.out_wire_1_1(vertical_tile_4_21_to_tile_5_21_1),
		.out_wire_1_2(vertical_tile_4_21_to_tile_5_21_2),
		.out_wire_1_3(vertical_tile_4_21_to_tile_5_21_3),
		.in_wire_1_0(vertical_tile_5_21_to_tile_4_21_0),
		.in_wire_1_1(vertical_tile_5_21_to_tile_4_21_1),
		.in_wire_1_2(vertical_tile_5_21_to_tile_4_21_2),
		.in_wire_1_3(vertical_tile_5_21_to_tile_4_21_3),
		.out_wire_2_0(horizontal_tile_4_21_to_tile_4_20_0),
		.out_wire_2_1(horizontal_tile_4_21_to_tile_4_20_1),
		.out_wire_2_2(horizontal_tile_4_21_to_tile_4_20_2),
		.out_wire_2_3(horizontal_tile_4_21_to_tile_4_20_3),
		.in_wire_2_0(horizontal_tile_4_20_to_tile_4_21_0),
		.in_wire_2_1(horizontal_tile_4_20_to_tile_4_21_1),
		.in_wire_2_2(horizontal_tile_4_20_to_tile_4_21_2),
		.in_wire_2_3(horizontal_tile_4_20_to_tile_4_21_3),
		.out_wire_0_0(horizontal_tile_4_21_to_tile_4_22_0),
		.out_wire_0_1(horizontal_tile_4_21_to_tile_4_22_1),
		.out_wire_0_2(horizontal_tile_4_21_to_tile_4_22_2),
		.out_wire_0_3(horizontal_tile_4_21_to_tile_4_22_3),
		.in_wire_0_0(horizontal_tile_4_22_to_tile_4_21_0),
		.in_wire_0_1(horizontal_tile_4_22_to_tile_4_21_1),
		.in_wire_0_2(horizontal_tile_4_22_to_tile_4_21_2),
		.in_wire_0_3(horizontal_tile_4_22_to_tile_4_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(150)
	);

	pe_tile pe_tile_4_22(
		.out_wire_3_0(vertical_tile_4_22_to_tile_3_22_0),
		.out_wire_3_1(vertical_tile_4_22_to_tile_3_22_1),
		.out_wire_3_2(vertical_tile_4_22_to_tile_3_22_2),
		.out_wire_3_3(vertical_tile_4_22_to_tile_3_22_3),
		.in_wire_3_0(vertical_tile_3_22_to_tile_4_22_0),
		.in_wire_3_1(vertical_tile_3_22_to_tile_4_22_1),
		.in_wire_3_2(vertical_tile_3_22_to_tile_4_22_2),
		.in_wire_3_3(vertical_tile_3_22_to_tile_4_22_3),
		.out_wire_1_0(vertical_tile_4_22_to_tile_5_22_0),
		.out_wire_1_1(vertical_tile_4_22_to_tile_5_22_1),
		.out_wire_1_2(vertical_tile_4_22_to_tile_5_22_2),
		.out_wire_1_3(vertical_tile_4_22_to_tile_5_22_3),
		.in_wire_1_0(vertical_tile_5_22_to_tile_4_22_0),
		.in_wire_1_1(vertical_tile_5_22_to_tile_4_22_1),
		.in_wire_1_2(vertical_tile_5_22_to_tile_4_22_2),
		.in_wire_1_3(vertical_tile_5_22_to_tile_4_22_3),
		.out_wire_2_0(horizontal_tile_4_22_to_tile_4_21_0),
		.out_wire_2_1(horizontal_tile_4_22_to_tile_4_21_1),
		.out_wire_2_2(horizontal_tile_4_22_to_tile_4_21_2),
		.out_wire_2_3(horizontal_tile_4_22_to_tile_4_21_3),
		.in_wire_2_0(horizontal_tile_4_21_to_tile_4_22_0),
		.in_wire_2_1(horizontal_tile_4_21_to_tile_4_22_1),
		.in_wire_2_2(horizontal_tile_4_21_to_tile_4_22_2),
		.in_wire_2_3(horizontal_tile_4_21_to_tile_4_22_3),
		.out_wire_0_0(horizontal_tile_4_22_to_tile_4_23_0),
		.out_wire_0_1(horizontal_tile_4_22_to_tile_4_23_1),
		.out_wire_0_2(horizontal_tile_4_22_to_tile_4_23_2),
		.out_wire_0_3(horizontal_tile_4_22_to_tile_4_23_3),
		.in_wire_0_0(horizontal_tile_4_23_to_tile_4_22_0),
		.in_wire_0_1(horizontal_tile_4_23_to_tile_4_22_1),
		.in_wire_0_2(horizontal_tile_4_23_to_tile_4_22_2),
		.in_wire_0_3(horizontal_tile_4_23_to_tile_4_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(151)
	);

	pe_tile pe_tile_4_23(
		.out_wire_3_0(vertical_tile_4_23_to_tile_3_23_0),
		.out_wire_3_1(vertical_tile_4_23_to_tile_3_23_1),
		.out_wire_3_2(vertical_tile_4_23_to_tile_3_23_2),
		.out_wire_3_3(vertical_tile_4_23_to_tile_3_23_3),
		.in_wire_3_0(vertical_tile_3_23_to_tile_4_23_0),
		.in_wire_3_1(vertical_tile_3_23_to_tile_4_23_1),
		.in_wire_3_2(vertical_tile_3_23_to_tile_4_23_2),
		.in_wire_3_3(vertical_tile_3_23_to_tile_4_23_3),
		.out_wire_1_0(vertical_tile_4_23_to_tile_5_23_0),
		.out_wire_1_1(vertical_tile_4_23_to_tile_5_23_1),
		.out_wire_1_2(vertical_tile_4_23_to_tile_5_23_2),
		.out_wire_1_3(vertical_tile_4_23_to_tile_5_23_3),
		.in_wire_1_0(vertical_tile_5_23_to_tile_4_23_0),
		.in_wire_1_1(vertical_tile_5_23_to_tile_4_23_1),
		.in_wire_1_2(vertical_tile_5_23_to_tile_4_23_2),
		.in_wire_1_3(vertical_tile_5_23_to_tile_4_23_3),
		.out_wire_2_0(horizontal_tile_4_23_to_tile_4_22_0),
		.out_wire_2_1(horizontal_tile_4_23_to_tile_4_22_1),
		.out_wire_2_2(horizontal_tile_4_23_to_tile_4_22_2),
		.out_wire_2_3(horizontal_tile_4_23_to_tile_4_22_3),
		.in_wire_2_0(horizontal_tile_4_22_to_tile_4_23_0),
		.in_wire_2_1(horizontal_tile_4_22_to_tile_4_23_1),
		.in_wire_2_2(horizontal_tile_4_22_to_tile_4_23_2),
		.in_wire_2_3(horizontal_tile_4_22_to_tile_4_23_3),
		.out_wire_0_0(horizontal_tile_4_23_to_tile_4_24_0),
		.out_wire_0_1(horizontal_tile_4_23_to_tile_4_24_1),
		.out_wire_0_2(horizontal_tile_4_23_to_tile_4_24_2),
		.out_wire_0_3(horizontal_tile_4_23_to_tile_4_24_3),
		.in_wire_0_0(horizontal_tile_4_24_to_tile_4_23_0),
		.in_wire_0_1(horizontal_tile_4_24_to_tile_4_23_1),
		.in_wire_0_2(horizontal_tile_4_24_to_tile_4_23_2),
		.in_wire_0_3(horizontal_tile_4_24_to_tile_4_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(152)
	);

	pe_tile pe_tile_4_24(
		.out_wire_3_0(vertical_tile_4_24_to_tile_3_24_0),
		.out_wire_3_1(vertical_tile_4_24_to_tile_3_24_1),
		.out_wire_3_2(vertical_tile_4_24_to_tile_3_24_2),
		.out_wire_3_3(vertical_tile_4_24_to_tile_3_24_3),
		.in_wire_3_0(vertical_tile_3_24_to_tile_4_24_0),
		.in_wire_3_1(vertical_tile_3_24_to_tile_4_24_1),
		.in_wire_3_2(vertical_tile_3_24_to_tile_4_24_2),
		.in_wire_3_3(vertical_tile_3_24_to_tile_4_24_3),
		.out_wire_1_0(vertical_tile_4_24_to_tile_5_24_0),
		.out_wire_1_1(vertical_tile_4_24_to_tile_5_24_1),
		.out_wire_1_2(vertical_tile_4_24_to_tile_5_24_2),
		.out_wire_1_3(vertical_tile_4_24_to_tile_5_24_3),
		.in_wire_1_0(vertical_tile_5_24_to_tile_4_24_0),
		.in_wire_1_1(vertical_tile_5_24_to_tile_4_24_1),
		.in_wire_1_2(vertical_tile_5_24_to_tile_4_24_2),
		.in_wire_1_3(vertical_tile_5_24_to_tile_4_24_3),
		.out_wire_2_0(horizontal_tile_4_24_to_tile_4_23_0),
		.out_wire_2_1(horizontal_tile_4_24_to_tile_4_23_1),
		.out_wire_2_2(horizontal_tile_4_24_to_tile_4_23_2),
		.out_wire_2_3(horizontal_tile_4_24_to_tile_4_23_3),
		.in_wire_2_0(horizontal_tile_4_23_to_tile_4_24_0),
		.in_wire_2_1(horizontal_tile_4_23_to_tile_4_24_1),
		.in_wire_2_2(horizontal_tile_4_23_to_tile_4_24_2),
		.in_wire_2_3(horizontal_tile_4_23_to_tile_4_24_3),
		.out_wire_0_0(horizontal_tile_4_24_to_tile_4_25_0),
		.out_wire_0_1(horizontal_tile_4_24_to_tile_4_25_1),
		.out_wire_0_2(horizontal_tile_4_24_to_tile_4_25_2),
		.out_wire_0_3(horizontal_tile_4_24_to_tile_4_25_3),
		.in_wire_0_0(horizontal_tile_4_25_to_tile_4_24_0),
		.in_wire_0_1(horizontal_tile_4_25_to_tile_4_24_1),
		.in_wire_0_2(horizontal_tile_4_25_to_tile_4_24_2),
		.in_wire_0_3(horizontal_tile_4_25_to_tile_4_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(153)
	);

	pe_tile pe_tile_4_25(
		.out_wire_3_0(vertical_tile_4_25_to_tile_3_25_0),
		.out_wire_3_1(vertical_tile_4_25_to_tile_3_25_1),
		.out_wire_3_2(vertical_tile_4_25_to_tile_3_25_2),
		.out_wire_3_3(vertical_tile_4_25_to_tile_3_25_3),
		.in_wire_3_0(vertical_tile_3_25_to_tile_4_25_0),
		.in_wire_3_1(vertical_tile_3_25_to_tile_4_25_1),
		.in_wire_3_2(vertical_tile_3_25_to_tile_4_25_2),
		.in_wire_3_3(vertical_tile_3_25_to_tile_4_25_3),
		.out_wire_1_0(vertical_tile_4_25_to_tile_5_25_0),
		.out_wire_1_1(vertical_tile_4_25_to_tile_5_25_1),
		.out_wire_1_2(vertical_tile_4_25_to_tile_5_25_2),
		.out_wire_1_3(vertical_tile_4_25_to_tile_5_25_3),
		.in_wire_1_0(vertical_tile_5_25_to_tile_4_25_0),
		.in_wire_1_1(vertical_tile_5_25_to_tile_4_25_1),
		.in_wire_1_2(vertical_tile_5_25_to_tile_4_25_2),
		.in_wire_1_3(vertical_tile_5_25_to_tile_4_25_3),
		.out_wire_2_0(horizontal_tile_4_25_to_tile_4_24_0),
		.out_wire_2_1(horizontal_tile_4_25_to_tile_4_24_1),
		.out_wire_2_2(horizontal_tile_4_25_to_tile_4_24_2),
		.out_wire_2_3(horizontal_tile_4_25_to_tile_4_24_3),
		.in_wire_2_0(horizontal_tile_4_24_to_tile_4_25_0),
		.in_wire_2_1(horizontal_tile_4_24_to_tile_4_25_1),
		.in_wire_2_2(horizontal_tile_4_24_to_tile_4_25_2),
		.in_wire_2_3(horizontal_tile_4_24_to_tile_4_25_3),
		.out_wire_0_0(horizontal_tile_4_25_to_tile_4_26_0),
		.out_wire_0_1(horizontal_tile_4_25_to_tile_4_26_1),
		.out_wire_0_2(horizontal_tile_4_25_to_tile_4_26_2),
		.out_wire_0_3(horizontal_tile_4_25_to_tile_4_26_3),
		.in_wire_0_0(horizontal_tile_4_26_to_tile_4_25_0),
		.in_wire_0_1(horizontal_tile_4_26_to_tile_4_25_1),
		.in_wire_0_2(horizontal_tile_4_26_to_tile_4_25_2),
		.in_wire_0_3(horizontal_tile_4_26_to_tile_4_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(154)
	);

	pe_tile pe_tile_4_26(
		.out_wire_3_0(vertical_tile_4_26_to_tile_3_26_0),
		.out_wire_3_1(vertical_tile_4_26_to_tile_3_26_1),
		.out_wire_3_2(vertical_tile_4_26_to_tile_3_26_2),
		.out_wire_3_3(vertical_tile_4_26_to_tile_3_26_3),
		.in_wire_3_0(vertical_tile_3_26_to_tile_4_26_0),
		.in_wire_3_1(vertical_tile_3_26_to_tile_4_26_1),
		.in_wire_3_2(vertical_tile_3_26_to_tile_4_26_2),
		.in_wire_3_3(vertical_tile_3_26_to_tile_4_26_3),
		.out_wire_1_0(vertical_tile_4_26_to_tile_5_26_0),
		.out_wire_1_1(vertical_tile_4_26_to_tile_5_26_1),
		.out_wire_1_2(vertical_tile_4_26_to_tile_5_26_2),
		.out_wire_1_3(vertical_tile_4_26_to_tile_5_26_3),
		.in_wire_1_0(vertical_tile_5_26_to_tile_4_26_0),
		.in_wire_1_1(vertical_tile_5_26_to_tile_4_26_1),
		.in_wire_1_2(vertical_tile_5_26_to_tile_4_26_2),
		.in_wire_1_3(vertical_tile_5_26_to_tile_4_26_3),
		.out_wire_2_0(horizontal_tile_4_26_to_tile_4_25_0),
		.out_wire_2_1(horizontal_tile_4_26_to_tile_4_25_1),
		.out_wire_2_2(horizontal_tile_4_26_to_tile_4_25_2),
		.out_wire_2_3(horizontal_tile_4_26_to_tile_4_25_3),
		.in_wire_2_0(horizontal_tile_4_25_to_tile_4_26_0),
		.in_wire_2_1(horizontal_tile_4_25_to_tile_4_26_1),
		.in_wire_2_2(horizontal_tile_4_25_to_tile_4_26_2),
		.in_wire_2_3(horizontal_tile_4_25_to_tile_4_26_3),
		.out_wire_0_0(horizontal_tile_4_26_to_tile_4_27_0),
		.out_wire_0_1(horizontal_tile_4_26_to_tile_4_27_1),
		.out_wire_0_2(horizontal_tile_4_26_to_tile_4_27_2),
		.out_wire_0_3(horizontal_tile_4_26_to_tile_4_27_3),
		.in_wire_0_0(horizontal_tile_4_27_to_tile_4_26_0),
		.in_wire_0_1(horizontal_tile_4_27_to_tile_4_26_1),
		.in_wire_0_2(horizontal_tile_4_27_to_tile_4_26_2),
		.in_wire_0_3(horizontal_tile_4_27_to_tile_4_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(155)
	);

	pe_tile pe_tile_4_27(
		.out_wire_3_0(vertical_tile_4_27_to_tile_3_27_0),
		.out_wire_3_1(vertical_tile_4_27_to_tile_3_27_1),
		.out_wire_3_2(vertical_tile_4_27_to_tile_3_27_2),
		.out_wire_3_3(vertical_tile_4_27_to_tile_3_27_3),
		.in_wire_3_0(vertical_tile_3_27_to_tile_4_27_0),
		.in_wire_3_1(vertical_tile_3_27_to_tile_4_27_1),
		.in_wire_3_2(vertical_tile_3_27_to_tile_4_27_2),
		.in_wire_3_3(vertical_tile_3_27_to_tile_4_27_3),
		.out_wire_1_0(vertical_tile_4_27_to_tile_5_27_0),
		.out_wire_1_1(vertical_tile_4_27_to_tile_5_27_1),
		.out_wire_1_2(vertical_tile_4_27_to_tile_5_27_2),
		.out_wire_1_3(vertical_tile_4_27_to_tile_5_27_3),
		.in_wire_1_0(vertical_tile_5_27_to_tile_4_27_0),
		.in_wire_1_1(vertical_tile_5_27_to_tile_4_27_1),
		.in_wire_1_2(vertical_tile_5_27_to_tile_4_27_2),
		.in_wire_1_3(vertical_tile_5_27_to_tile_4_27_3),
		.out_wire_2_0(horizontal_tile_4_27_to_tile_4_26_0),
		.out_wire_2_1(horizontal_tile_4_27_to_tile_4_26_1),
		.out_wire_2_2(horizontal_tile_4_27_to_tile_4_26_2),
		.out_wire_2_3(horizontal_tile_4_27_to_tile_4_26_3),
		.in_wire_2_0(horizontal_tile_4_26_to_tile_4_27_0),
		.in_wire_2_1(horizontal_tile_4_26_to_tile_4_27_1),
		.in_wire_2_2(horizontal_tile_4_26_to_tile_4_27_2),
		.in_wire_2_3(horizontal_tile_4_26_to_tile_4_27_3),
		.out_wire_0_0(horizontal_tile_4_27_to_tile_4_28_0),
		.out_wire_0_1(horizontal_tile_4_27_to_tile_4_28_1),
		.out_wire_0_2(horizontal_tile_4_27_to_tile_4_28_2),
		.out_wire_0_3(horizontal_tile_4_27_to_tile_4_28_3),
		.in_wire_0_0(horizontal_tile_4_28_to_tile_4_27_0),
		.in_wire_0_1(horizontal_tile_4_28_to_tile_4_27_1),
		.in_wire_0_2(horizontal_tile_4_28_to_tile_4_27_2),
		.in_wire_0_3(horizontal_tile_4_28_to_tile_4_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(156)
	);

	pe_tile pe_tile_4_28(
		.out_wire_3_0(vertical_tile_4_28_to_tile_3_28_0),
		.out_wire_3_1(vertical_tile_4_28_to_tile_3_28_1),
		.out_wire_3_2(vertical_tile_4_28_to_tile_3_28_2),
		.out_wire_3_3(vertical_tile_4_28_to_tile_3_28_3),
		.in_wire_3_0(vertical_tile_3_28_to_tile_4_28_0),
		.in_wire_3_1(vertical_tile_3_28_to_tile_4_28_1),
		.in_wire_3_2(vertical_tile_3_28_to_tile_4_28_2),
		.in_wire_3_3(vertical_tile_3_28_to_tile_4_28_3),
		.out_wire_1_0(vertical_tile_4_28_to_tile_5_28_0),
		.out_wire_1_1(vertical_tile_4_28_to_tile_5_28_1),
		.out_wire_1_2(vertical_tile_4_28_to_tile_5_28_2),
		.out_wire_1_3(vertical_tile_4_28_to_tile_5_28_3),
		.in_wire_1_0(vertical_tile_5_28_to_tile_4_28_0),
		.in_wire_1_1(vertical_tile_5_28_to_tile_4_28_1),
		.in_wire_1_2(vertical_tile_5_28_to_tile_4_28_2),
		.in_wire_1_3(vertical_tile_5_28_to_tile_4_28_3),
		.out_wire_2_0(horizontal_tile_4_28_to_tile_4_27_0),
		.out_wire_2_1(horizontal_tile_4_28_to_tile_4_27_1),
		.out_wire_2_2(horizontal_tile_4_28_to_tile_4_27_2),
		.out_wire_2_3(horizontal_tile_4_28_to_tile_4_27_3),
		.in_wire_2_0(horizontal_tile_4_27_to_tile_4_28_0),
		.in_wire_2_1(horizontal_tile_4_27_to_tile_4_28_1),
		.in_wire_2_2(horizontal_tile_4_27_to_tile_4_28_2),
		.in_wire_2_3(horizontal_tile_4_27_to_tile_4_28_3),
		.out_wire_0_0(horizontal_tile_4_28_to_tile_4_29_0),
		.out_wire_0_1(horizontal_tile_4_28_to_tile_4_29_1),
		.out_wire_0_2(horizontal_tile_4_28_to_tile_4_29_2),
		.out_wire_0_3(horizontal_tile_4_28_to_tile_4_29_3),
		.in_wire_0_0(horizontal_tile_4_29_to_tile_4_28_0),
		.in_wire_0_1(horizontal_tile_4_29_to_tile_4_28_1),
		.in_wire_0_2(horizontal_tile_4_29_to_tile_4_28_2),
		.in_wire_0_3(horizontal_tile_4_29_to_tile_4_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(157)
	);

	pe_tile pe_tile_4_29(
		.out_wire_3_0(vertical_tile_4_29_to_tile_3_29_0),
		.out_wire_3_1(vertical_tile_4_29_to_tile_3_29_1),
		.out_wire_3_2(vertical_tile_4_29_to_tile_3_29_2),
		.out_wire_3_3(vertical_tile_4_29_to_tile_3_29_3),
		.in_wire_3_0(vertical_tile_3_29_to_tile_4_29_0),
		.in_wire_3_1(vertical_tile_3_29_to_tile_4_29_1),
		.in_wire_3_2(vertical_tile_3_29_to_tile_4_29_2),
		.in_wire_3_3(vertical_tile_3_29_to_tile_4_29_3),
		.out_wire_1_0(vertical_tile_4_29_to_tile_5_29_0),
		.out_wire_1_1(vertical_tile_4_29_to_tile_5_29_1),
		.out_wire_1_2(vertical_tile_4_29_to_tile_5_29_2),
		.out_wire_1_3(vertical_tile_4_29_to_tile_5_29_3),
		.in_wire_1_0(vertical_tile_5_29_to_tile_4_29_0),
		.in_wire_1_1(vertical_tile_5_29_to_tile_4_29_1),
		.in_wire_1_2(vertical_tile_5_29_to_tile_4_29_2),
		.in_wire_1_3(vertical_tile_5_29_to_tile_4_29_3),
		.out_wire_2_0(horizontal_tile_4_29_to_tile_4_28_0),
		.out_wire_2_1(horizontal_tile_4_29_to_tile_4_28_1),
		.out_wire_2_2(horizontal_tile_4_29_to_tile_4_28_2),
		.out_wire_2_3(horizontal_tile_4_29_to_tile_4_28_3),
		.in_wire_2_0(horizontal_tile_4_28_to_tile_4_29_0),
		.in_wire_2_1(horizontal_tile_4_28_to_tile_4_29_1),
		.in_wire_2_2(horizontal_tile_4_28_to_tile_4_29_2),
		.in_wire_2_3(horizontal_tile_4_28_to_tile_4_29_3),
		.out_wire_0_0(horizontal_tile_4_29_to_tile_4_30_0),
		.out_wire_0_1(horizontal_tile_4_29_to_tile_4_30_1),
		.out_wire_0_2(horizontal_tile_4_29_to_tile_4_30_2),
		.out_wire_0_3(horizontal_tile_4_29_to_tile_4_30_3),
		.in_wire_0_0(horizontal_tile_4_30_to_tile_4_29_0),
		.in_wire_0_1(horizontal_tile_4_30_to_tile_4_29_1),
		.in_wire_0_2(horizontal_tile_4_30_to_tile_4_29_2),
		.in_wire_0_3(horizontal_tile_4_30_to_tile_4_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(158)
	);

	pe_tile pe_tile_4_30(
		.out_wire_3_0(vertical_tile_4_30_to_tile_3_30_0),
		.out_wire_3_1(vertical_tile_4_30_to_tile_3_30_1),
		.out_wire_3_2(vertical_tile_4_30_to_tile_3_30_2),
		.out_wire_3_3(vertical_tile_4_30_to_tile_3_30_3),
		.in_wire_3_0(vertical_tile_3_30_to_tile_4_30_0),
		.in_wire_3_1(vertical_tile_3_30_to_tile_4_30_1),
		.in_wire_3_2(vertical_tile_3_30_to_tile_4_30_2),
		.in_wire_3_3(vertical_tile_3_30_to_tile_4_30_3),
		.out_wire_1_0(vertical_tile_4_30_to_tile_5_30_0),
		.out_wire_1_1(vertical_tile_4_30_to_tile_5_30_1),
		.out_wire_1_2(vertical_tile_4_30_to_tile_5_30_2),
		.out_wire_1_3(vertical_tile_4_30_to_tile_5_30_3),
		.in_wire_1_0(vertical_tile_5_30_to_tile_4_30_0),
		.in_wire_1_1(vertical_tile_5_30_to_tile_4_30_1),
		.in_wire_1_2(vertical_tile_5_30_to_tile_4_30_2),
		.in_wire_1_3(vertical_tile_5_30_to_tile_4_30_3),
		.out_wire_2_0(horizontal_tile_4_30_to_tile_4_29_0),
		.out_wire_2_1(horizontal_tile_4_30_to_tile_4_29_1),
		.out_wire_2_2(horizontal_tile_4_30_to_tile_4_29_2),
		.out_wire_2_3(horizontal_tile_4_30_to_tile_4_29_3),
		.in_wire_2_0(horizontal_tile_4_29_to_tile_4_30_0),
		.in_wire_2_1(horizontal_tile_4_29_to_tile_4_30_1),
		.in_wire_2_2(horizontal_tile_4_29_to_tile_4_30_2),
		.in_wire_2_3(horizontal_tile_4_29_to_tile_4_30_3),
		.out_wire_0_0(horizontal_tile_4_30_to_tile_4_31_0),
		.out_wire_0_1(horizontal_tile_4_30_to_tile_4_31_1),
		.out_wire_0_2(horizontal_tile_4_30_to_tile_4_31_2),
		.out_wire_0_3(horizontal_tile_4_30_to_tile_4_31_3),
		.in_wire_0_0(horizontal_tile_4_31_to_tile_4_30_0),
		.in_wire_0_1(horizontal_tile_4_31_to_tile_4_30_1),
		.in_wire_0_2(horizontal_tile_4_31_to_tile_4_30_2),
		.in_wire_0_3(horizontal_tile_4_31_to_tile_4_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(159)
	);

	pe_tile_right pe_tile_4_31(
		.out_wire_3_0(vertical_tile_4_31_to_tile_3_31_0),
		.out_wire_3_1(vertical_tile_4_31_to_tile_3_31_1),
		.out_wire_3_2(vertical_tile_4_31_to_tile_3_31_2),
		.out_wire_3_3(vertical_tile_4_31_to_tile_3_31_3),
		.in_wire_3_0(vertical_tile_3_31_to_tile_4_31_0),
		.in_wire_3_1(vertical_tile_3_31_to_tile_4_31_1),
		.in_wire_3_2(vertical_tile_3_31_to_tile_4_31_2),
		.in_wire_3_3(vertical_tile_3_31_to_tile_4_31_3),
		.out_wire_1_0(vertical_tile_4_31_to_tile_5_31_0),
		.out_wire_1_1(vertical_tile_4_31_to_tile_5_31_1),
		.out_wire_1_2(vertical_tile_4_31_to_tile_5_31_2),
		.out_wire_1_3(vertical_tile_4_31_to_tile_5_31_3),
		.in_wire_1_0(vertical_tile_5_31_to_tile_4_31_0),
		.in_wire_1_1(vertical_tile_5_31_to_tile_4_31_1),
		.in_wire_1_2(vertical_tile_5_31_to_tile_4_31_2),
		.in_wire_1_3(vertical_tile_5_31_to_tile_4_31_3),
		.out_wire_2_0(horizontal_tile_4_31_to_tile_4_30_0),
		.out_wire_2_1(horizontal_tile_4_31_to_tile_4_30_1),
		.out_wire_2_2(horizontal_tile_4_31_to_tile_4_30_2),
		.out_wire_2_3(horizontal_tile_4_31_to_tile_4_30_3),
		.in_wire_2_0(horizontal_tile_4_30_to_tile_4_31_0),
		.in_wire_2_1(horizontal_tile_4_30_to_tile_4_31_1),
		.in_wire_2_2(horizontal_tile_4_30_to_tile_4_31_2),
		.in_wire_2_3(horizontal_tile_4_30_to_tile_4_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(160)
	);

	pe_tile_left pe_tile_5_0(
		.out_wire_3_0(vertical_tile_5_0_to_tile_4_0_0),
		.out_wire_3_1(vertical_tile_5_0_to_tile_4_0_1),
		.out_wire_3_2(vertical_tile_5_0_to_tile_4_0_2),
		.out_wire_3_3(vertical_tile_5_0_to_tile_4_0_3),
		.in_wire_3_0(vertical_tile_4_0_to_tile_5_0_0),
		.in_wire_3_1(vertical_tile_4_0_to_tile_5_0_1),
		.in_wire_3_2(vertical_tile_4_0_to_tile_5_0_2),
		.in_wire_3_3(vertical_tile_4_0_to_tile_5_0_3),
		.out_wire_1_0(vertical_tile_5_0_to_tile_6_0_0),
		.out_wire_1_1(vertical_tile_5_0_to_tile_6_0_1),
		.out_wire_1_2(vertical_tile_5_0_to_tile_6_0_2),
		.out_wire_1_3(vertical_tile_5_0_to_tile_6_0_3),
		.in_wire_1_0(vertical_tile_6_0_to_tile_5_0_0),
		.in_wire_1_1(vertical_tile_6_0_to_tile_5_0_1),
		.in_wire_1_2(vertical_tile_6_0_to_tile_5_0_2),
		.in_wire_1_3(vertical_tile_6_0_to_tile_5_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_5_0_to_tile_5_1_0),
		.out_wire_0_1(horizontal_tile_5_0_to_tile_5_1_1),
		.out_wire_0_2(horizontal_tile_5_0_to_tile_5_1_2),
		.out_wire_0_3(horizontal_tile_5_0_to_tile_5_1_3),
		.in_wire_0_0(horizontal_tile_5_1_to_tile_5_0_0),
		.in_wire_0_1(horizontal_tile_5_1_to_tile_5_0_1),
		.in_wire_0_2(horizontal_tile_5_1_to_tile_5_0_2),
		.in_wire_0_3(horizontal_tile_5_1_to_tile_5_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(161)
	);

	pe_tile pe_tile_5_1(
		.out_wire_3_0(vertical_tile_5_1_to_tile_4_1_0),
		.out_wire_3_1(vertical_tile_5_1_to_tile_4_1_1),
		.out_wire_3_2(vertical_tile_5_1_to_tile_4_1_2),
		.out_wire_3_3(vertical_tile_5_1_to_tile_4_1_3),
		.in_wire_3_0(vertical_tile_4_1_to_tile_5_1_0),
		.in_wire_3_1(vertical_tile_4_1_to_tile_5_1_1),
		.in_wire_3_2(vertical_tile_4_1_to_tile_5_1_2),
		.in_wire_3_3(vertical_tile_4_1_to_tile_5_1_3),
		.out_wire_1_0(vertical_tile_5_1_to_tile_6_1_0),
		.out_wire_1_1(vertical_tile_5_1_to_tile_6_1_1),
		.out_wire_1_2(vertical_tile_5_1_to_tile_6_1_2),
		.out_wire_1_3(vertical_tile_5_1_to_tile_6_1_3),
		.in_wire_1_0(vertical_tile_6_1_to_tile_5_1_0),
		.in_wire_1_1(vertical_tile_6_1_to_tile_5_1_1),
		.in_wire_1_2(vertical_tile_6_1_to_tile_5_1_2),
		.in_wire_1_3(vertical_tile_6_1_to_tile_5_1_3),
		.out_wire_2_0(horizontal_tile_5_1_to_tile_5_0_0),
		.out_wire_2_1(horizontal_tile_5_1_to_tile_5_0_1),
		.out_wire_2_2(horizontal_tile_5_1_to_tile_5_0_2),
		.out_wire_2_3(horizontal_tile_5_1_to_tile_5_0_3),
		.in_wire_2_0(horizontal_tile_5_0_to_tile_5_1_0),
		.in_wire_2_1(horizontal_tile_5_0_to_tile_5_1_1),
		.in_wire_2_2(horizontal_tile_5_0_to_tile_5_1_2),
		.in_wire_2_3(horizontal_tile_5_0_to_tile_5_1_3),
		.out_wire_0_0(horizontal_tile_5_1_to_tile_5_2_0),
		.out_wire_0_1(horizontal_tile_5_1_to_tile_5_2_1),
		.out_wire_0_2(horizontal_tile_5_1_to_tile_5_2_2),
		.out_wire_0_3(horizontal_tile_5_1_to_tile_5_2_3),
		.in_wire_0_0(horizontal_tile_5_2_to_tile_5_1_0),
		.in_wire_0_1(horizontal_tile_5_2_to_tile_5_1_1),
		.in_wire_0_2(horizontal_tile_5_2_to_tile_5_1_2),
		.in_wire_0_3(horizontal_tile_5_2_to_tile_5_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(162)
	);

	pe_tile pe_tile_5_2(
		.out_wire_3_0(vertical_tile_5_2_to_tile_4_2_0),
		.out_wire_3_1(vertical_tile_5_2_to_tile_4_2_1),
		.out_wire_3_2(vertical_tile_5_2_to_tile_4_2_2),
		.out_wire_3_3(vertical_tile_5_2_to_tile_4_2_3),
		.in_wire_3_0(vertical_tile_4_2_to_tile_5_2_0),
		.in_wire_3_1(vertical_tile_4_2_to_tile_5_2_1),
		.in_wire_3_2(vertical_tile_4_2_to_tile_5_2_2),
		.in_wire_3_3(vertical_tile_4_2_to_tile_5_2_3),
		.out_wire_1_0(vertical_tile_5_2_to_tile_6_2_0),
		.out_wire_1_1(vertical_tile_5_2_to_tile_6_2_1),
		.out_wire_1_2(vertical_tile_5_2_to_tile_6_2_2),
		.out_wire_1_3(vertical_tile_5_2_to_tile_6_2_3),
		.in_wire_1_0(vertical_tile_6_2_to_tile_5_2_0),
		.in_wire_1_1(vertical_tile_6_2_to_tile_5_2_1),
		.in_wire_1_2(vertical_tile_6_2_to_tile_5_2_2),
		.in_wire_1_3(vertical_tile_6_2_to_tile_5_2_3),
		.out_wire_2_0(horizontal_tile_5_2_to_tile_5_1_0),
		.out_wire_2_1(horizontal_tile_5_2_to_tile_5_1_1),
		.out_wire_2_2(horizontal_tile_5_2_to_tile_5_1_2),
		.out_wire_2_3(horizontal_tile_5_2_to_tile_5_1_3),
		.in_wire_2_0(horizontal_tile_5_1_to_tile_5_2_0),
		.in_wire_2_1(horizontal_tile_5_1_to_tile_5_2_1),
		.in_wire_2_2(horizontal_tile_5_1_to_tile_5_2_2),
		.in_wire_2_3(horizontal_tile_5_1_to_tile_5_2_3),
		.out_wire_0_0(horizontal_tile_5_2_to_tile_5_3_0),
		.out_wire_0_1(horizontal_tile_5_2_to_tile_5_3_1),
		.out_wire_0_2(horizontal_tile_5_2_to_tile_5_3_2),
		.out_wire_0_3(horizontal_tile_5_2_to_tile_5_3_3),
		.in_wire_0_0(horizontal_tile_5_3_to_tile_5_2_0),
		.in_wire_0_1(horizontal_tile_5_3_to_tile_5_2_1),
		.in_wire_0_2(horizontal_tile_5_3_to_tile_5_2_2),
		.in_wire_0_3(horizontal_tile_5_3_to_tile_5_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(163)
	);

	pe_tile pe_tile_5_3(
		.out_wire_3_0(vertical_tile_5_3_to_tile_4_3_0),
		.out_wire_3_1(vertical_tile_5_3_to_tile_4_3_1),
		.out_wire_3_2(vertical_tile_5_3_to_tile_4_3_2),
		.out_wire_3_3(vertical_tile_5_3_to_tile_4_3_3),
		.in_wire_3_0(vertical_tile_4_3_to_tile_5_3_0),
		.in_wire_3_1(vertical_tile_4_3_to_tile_5_3_1),
		.in_wire_3_2(vertical_tile_4_3_to_tile_5_3_2),
		.in_wire_3_3(vertical_tile_4_3_to_tile_5_3_3),
		.out_wire_1_0(vertical_tile_5_3_to_tile_6_3_0),
		.out_wire_1_1(vertical_tile_5_3_to_tile_6_3_1),
		.out_wire_1_2(vertical_tile_5_3_to_tile_6_3_2),
		.out_wire_1_3(vertical_tile_5_3_to_tile_6_3_3),
		.in_wire_1_0(vertical_tile_6_3_to_tile_5_3_0),
		.in_wire_1_1(vertical_tile_6_3_to_tile_5_3_1),
		.in_wire_1_2(vertical_tile_6_3_to_tile_5_3_2),
		.in_wire_1_3(vertical_tile_6_3_to_tile_5_3_3),
		.out_wire_2_0(horizontal_tile_5_3_to_tile_5_2_0),
		.out_wire_2_1(horizontal_tile_5_3_to_tile_5_2_1),
		.out_wire_2_2(horizontal_tile_5_3_to_tile_5_2_2),
		.out_wire_2_3(horizontal_tile_5_3_to_tile_5_2_3),
		.in_wire_2_0(horizontal_tile_5_2_to_tile_5_3_0),
		.in_wire_2_1(horizontal_tile_5_2_to_tile_5_3_1),
		.in_wire_2_2(horizontal_tile_5_2_to_tile_5_3_2),
		.in_wire_2_3(horizontal_tile_5_2_to_tile_5_3_3),
		.out_wire_0_0(horizontal_tile_5_3_to_tile_5_4_0),
		.out_wire_0_1(horizontal_tile_5_3_to_tile_5_4_1),
		.out_wire_0_2(horizontal_tile_5_3_to_tile_5_4_2),
		.out_wire_0_3(horizontal_tile_5_3_to_tile_5_4_3),
		.in_wire_0_0(horizontal_tile_5_4_to_tile_5_3_0),
		.in_wire_0_1(horizontal_tile_5_4_to_tile_5_3_1),
		.in_wire_0_2(horizontal_tile_5_4_to_tile_5_3_2),
		.in_wire_0_3(horizontal_tile_5_4_to_tile_5_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(164)
	);

	pe_tile pe_tile_5_4(
		.out_wire_3_0(vertical_tile_5_4_to_tile_4_4_0),
		.out_wire_3_1(vertical_tile_5_4_to_tile_4_4_1),
		.out_wire_3_2(vertical_tile_5_4_to_tile_4_4_2),
		.out_wire_3_3(vertical_tile_5_4_to_tile_4_4_3),
		.in_wire_3_0(vertical_tile_4_4_to_tile_5_4_0),
		.in_wire_3_1(vertical_tile_4_4_to_tile_5_4_1),
		.in_wire_3_2(vertical_tile_4_4_to_tile_5_4_2),
		.in_wire_3_3(vertical_tile_4_4_to_tile_5_4_3),
		.out_wire_1_0(vertical_tile_5_4_to_tile_6_4_0),
		.out_wire_1_1(vertical_tile_5_4_to_tile_6_4_1),
		.out_wire_1_2(vertical_tile_5_4_to_tile_6_4_2),
		.out_wire_1_3(vertical_tile_5_4_to_tile_6_4_3),
		.in_wire_1_0(vertical_tile_6_4_to_tile_5_4_0),
		.in_wire_1_1(vertical_tile_6_4_to_tile_5_4_1),
		.in_wire_1_2(vertical_tile_6_4_to_tile_5_4_2),
		.in_wire_1_3(vertical_tile_6_4_to_tile_5_4_3),
		.out_wire_2_0(horizontal_tile_5_4_to_tile_5_3_0),
		.out_wire_2_1(horizontal_tile_5_4_to_tile_5_3_1),
		.out_wire_2_2(horizontal_tile_5_4_to_tile_5_3_2),
		.out_wire_2_3(horizontal_tile_5_4_to_tile_5_3_3),
		.in_wire_2_0(horizontal_tile_5_3_to_tile_5_4_0),
		.in_wire_2_1(horizontal_tile_5_3_to_tile_5_4_1),
		.in_wire_2_2(horizontal_tile_5_3_to_tile_5_4_2),
		.in_wire_2_3(horizontal_tile_5_3_to_tile_5_4_3),
		.out_wire_0_0(horizontal_tile_5_4_to_tile_5_5_0),
		.out_wire_0_1(horizontal_tile_5_4_to_tile_5_5_1),
		.out_wire_0_2(horizontal_tile_5_4_to_tile_5_5_2),
		.out_wire_0_3(horizontal_tile_5_4_to_tile_5_5_3),
		.in_wire_0_0(horizontal_tile_5_5_to_tile_5_4_0),
		.in_wire_0_1(horizontal_tile_5_5_to_tile_5_4_1),
		.in_wire_0_2(horizontal_tile_5_5_to_tile_5_4_2),
		.in_wire_0_3(horizontal_tile_5_5_to_tile_5_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(165)
	);

	pe_tile pe_tile_5_5(
		.out_wire_3_0(vertical_tile_5_5_to_tile_4_5_0),
		.out_wire_3_1(vertical_tile_5_5_to_tile_4_5_1),
		.out_wire_3_2(vertical_tile_5_5_to_tile_4_5_2),
		.out_wire_3_3(vertical_tile_5_5_to_tile_4_5_3),
		.in_wire_3_0(vertical_tile_4_5_to_tile_5_5_0),
		.in_wire_3_1(vertical_tile_4_5_to_tile_5_5_1),
		.in_wire_3_2(vertical_tile_4_5_to_tile_5_5_2),
		.in_wire_3_3(vertical_tile_4_5_to_tile_5_5_3),
		.out_wire_1_0(vertical_tile_5_5_to_tile_6_5_0),
		.out_wire_1_1(vertical_tile_5_5_to_tile_6_5_1),
		.out_wire_1_2(vertical_tile_5_5_to_tile_6_5_2),
		.out_wire_1_3(vertical_tile_5_5_to_tile_6_5_3),
		.in_wire_1_0(vertical_tile_6_5_to_tile_5_5_0),
		.in_wire_1_1(vertical_tile_6_5_to_tile_5_5_1),
		.in_wire_1_2(vertical_tile_6_5_to_tile_5_5_2),
		.in_wire_1_3(vertical_tile_6_5_to_tile_5_5_3),
		.out_wire_2_0(horizontal_tile_5_5_to_tile_5_4_0),
		.out_wire_2_1(horizontal_tile_5_5_to_tile_5_4_1),
		.out_wire_2_2(horizontal_tile_5_5_to_tile_5_4_2),
		.out_wire_2_3(horizontal_tile_5_5_to_tile_5_4_3),
		.in_wire_2_0(horizontal_tile_5_4_to_tile_5_5_0),
		.in_wire_2_1(horizontal_tile_5_4_to_tile_5_5_1),
		.in_wire_2_2(horizontal_tile_5_4_to_tile_5_5_2),
		.in_wire_2_3(horizontal_tile_5_4_to_tile_5_5_3),
		.out_wire_0_0(horizontal_tile_5_5_to_tile_5_6_0),
		.out_wire_0_1(horizontal_tile_5_5_to_tile_5_6_1),
		.out_wire_0_2(horizontal_tile_5_5_to_tile_5_6_2),
		.out_wire_0_3(horizontal_tile_5_5_to_tile_5_6_3),
		.in_wire_0_0(horizontal_tile_5_6_to_tile_5_5_0),
		.in_wire_0_1(horizontal_tile_5_6_to_tile_5_5_1),
		.in_wire_0_2(horizontal_tile_5_6_to_tile_5_5_2),
		.in_wire_0_3(horizontal_tile_5_6_to_tile_5_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(166)
	);

	pe_tile pe_tile_5_6(
		.out_wire_3_0(vertical_tile_5_6_to_tile_4_6_0),
		.out_wire_3_1(vertical_tile_5_6_to_tile_4_6_1),
		.out_wire_3_2(vertical_tile_5_6_to_tile_4_6_2),
		.out_wire_3_3(vertical_tile_5_6_to_tile_4_6_3),
		.in_wire_3_0(vertical_tile_4_6_to_tile_5_6_0),
		.in_wire_3_1(vertical_tile_4_6_to_tile_5_6_1),
		.in_wire_3_2(vertical_tile_4_6_to_tile_5_6_2),
		.in_wire_3_3(vertical_tile_4_6_to_tile_5_6_3),
		.out_wire_1_0(vertical_tile_5_6_to_tile_6_6_0),
		.out_wire_1_1(vertical_tile_5_6_to_tile_6_6_1),
		.out_wire_1_2(vertical_tile_5_6_to_tile_6_6_2),
		.out_wire_1_3(vertical_tile_5_6_to_tile_6_6_3),
		.in_wire_1_0(vertical_tile_6_6_to_tile_5_6_0),
		.in_wire_1_1(vertical_tile_6_6_to_tile_5_6_1),
		.in_wire_1_2(vertical_tile_6_6_to_tile_5_6_2),
		.in_wire_1_3(vertical_tile_6_6_to_tile_5_6_3),
		.out_wire_2_0(horizontal_tile_5_6_to_tile_5_5_0),
		.out_wire_2_1(horizontal_tile_5_6_to_tile_5_5_1),
		.out_wire_2_2(horizontal_tile_5_6_to_tile_5_5_2),
		.out_wire_2_3(horizontal_tile_5_6_to_tile_5_5_3),
		.in_wire_2_0(horizontal_tile_5_5_to_tile_5_6_0),
		.in_wire_2_1(horizontal_tile_5_5_to_tile_5_6_1),
		.in_wire_2_2(horizontal_tile_5_5_to_tile_5_6_2),
		.in_wire_2_3(horizontal_tile_5_5_to_tile_5_6_3),
		.out_wire_0_0(horizontal_tile_5_6_to_tile_5_7_0),
		.out_wire_0_1(horizontal_tile_5_6_to_tile_5_7_1),
		.out_wire_0_2(horizontal_tile_5_6_to_tile_5_7_2),
		.out_wire_0_3(horizontal_tile_5_6_to_tile_5_7_3),
		.in_wire_0_0(horizontal_tile_5_7_to_tile_5_6_0),
		.in_wire_0_1(horizontal_tile_5_7_to_tile_5_6_1),
		.in_wire_0_2(horizontal_tile_5_7_to_tile_5_6_2),
		.in_wire_0_3(horizontal_tile_5_7_to_tile_5_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(167)
	);

	pe_tile pe_tile_5_7(
		.out_wire_3_0(vertical_tile_5_7_to_tile_4_7_0),
		.out_wire_3_1(vertical_tile_5_7_to_tile_4_7_1),
		.out_wire_3_2(vertical_tile_5_7_to_tile_4_7_2),
		.out_wire_3_3(vertical_tile_5_7_to_tile_4_7_3),
		.in_wire_3_0(vertical_tile_4_7_to_tile_5_7_0),
		.in_wire_3_1(vertical_tile_4_7_to_tile_5_7_1),
		.in_wire_3_2(vertical_tile_4_7_to_tile_5_7_2),
		.in_wire_3_3(vertical_tile_4_7_to_tile_5_7_3),
		.out_wire_1_0(vertical_tile_5_7_to_tile_6_7_0),
		.out_wire_1_1(vertical_tile_5_7_to_tile_6_7_1),
		.out_wire_1_2(vertical_tile_5_7_to_tile_6_7_2),
		.out_wire_1_3(vertical_tile_5_7_to_tile_6_7_3),
		.in_wire_1_0(vertical_tile_6_7_to_tile_5_7_0),
		.in_wire_1_1(vertical_tile_6_7_to_tile_5_7_1),
		.in_wire_1_2(vertical_tile_6_7_to_tile_5_7_2),
		.in_wire_1_3(vertical_tile_6_7_to_tile_5_7_3),
		.out_wire_2_0(horizontal_tile_5_7_to_tile_5_6_0),
		.out_wire_2_1(horizontal_tile_5_7_to_tile_5_6_1),
		.out_wire_2_2(horizontal_tile_5_7_to_tile_5_6_2),
		.out_wire_2_3(horizontal_tile_5_7_to_tile_5_6_3),
		.in_wire_2_0(horizontal_tile_5_6_to_tile_5_7_0),
		.in_wire_2_1(horizontal_tile_5_6_to_tile_5_7_1),
		.in_wire_2_2(horizontal_tile_5_6_to_tile_5_7_2),
		.in_wire_2_3(horizontal_tile_5_6_to_tile_5_7_3),
		.out_wire_0_0(horizontal_tile_5_7_to_tile_5_8_0),
		.out_wire_0_1(horizontal_tile_5_7_to_tile_5_8_1),
		.out_wire_0_2(horizontal_tile_5_7_to_tile_5_8_2),
		.out_wire_0_3(horizontal_tile_5_7_to_tile_5_8_3),
		.in_wire_0_0(horizontal_tile_5_8_to_tile_5_7_0),
		.in_wire_0_1(horizontal_tile_5_8_to_tile_5_7_1),
		.in_wire_0_2(horizontal_tile_5_8_to_tile_5_7_2),
		.in_wire_0_3(horizontal_tile_5_8_to_tile_5_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(168)
	);

	pe_tile pe_tile_5_8(
		.out_wire_3_0(vertical_tile_5_8_to_tile_4_8_0),
		.out_wire_3_1(vertical_tile_5_8_to_tile_4_8_1),
		.out_wire_3_2(vertical_tile_5_8_to_tile_4_8_2),
		.out_wire_3_3(vertical_tile_5_8_to_tile_4_8_3),
		.in_wire_3_0(vertical_tile_4_8_to_tile_5_8_0),
		.in_wire_3_1(vertical_tile_4_8_to_tile_5_8_1),
		.in_wire_3_2(vertical_tile_4_8_to_tile_5_8_2),
		.in_wire_3_3(vertical_tile_4_8_to_tile_5_8_3),
		.out_wire_1_0(vertical_tile_5_8_to_tile_6_8_0),
		.out_wire_1_1(vertical_tile_5_8_to_tile_6_8_1),
		.out_wire_1_2(vertical_tile_5_8_to_tile_6_8_2),
		.out_wire_1_3(vertical_tile_5_8_to_tile_6_8_3),
		.in_wire_1_0(vertical_tile_6_8_to_tile_5_8_0),
		.in_wire_1_1(vertical_tile_6_8_to_tile_5_8_1),
		.in_wire_1_2(vertical_tile_6_8_to_tile_5_8_2),
		.in_wire_1_3(vertical_tile_6_8_to_tile_5_8_3),
		.out_wire_2_0(horizontal_tile_5_8_to_tile_5_7_0),
		.out_wire_2_1(horizontal_tile_5_8_to_tile_5_7_1),
		.out_wire_2_2(horizontal_tile_5_8_to_tile_5_7_2),
		.out_wire_2_3(horizontal_tile_5_8_to_tile_5_7_3),
		.in_wire_2_0(horizontal_tile_5_7_to_tile_5_8_0),
		.in_wire_2_1(horizontal_tile_5_7_to_tile_5_8_1),
		.in_wire_2_2(horizontal_tile_5_7_to_tile_5_8_2),
		.in_wire_2_3(horizontal_tile_5_7_to_tile_5_8_3),
		.out_wire_0_0(horizontal_tile_5_8_to_tile_5_9_0),
		.out_wire_0_1(horizontal_tile_5_8_to_tile_5_9_1),
		.out_wire_0_2(horizontal_tile_5_8_to_tile_5_9_2),
		.out_wire_0_3(horizontal_tile_5_8_to_tile_5_9_3),
		.in_wire_0_0(horizontal_tile_5_9_to_tile_5_8_0),
		.in_wire_0_1(horizontal_tile_5_9_to_tile_5_8_1),
		.in_wire_0_2(horizontal_tile_5_9_to_tile_5_8_2),
		.in_wire_0_3(horizontal_tile_5_9_to_tile_5_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(169)
	);

	pe_tile pe_tile_5_9(
		.out_wire_3_0(vertical_tile_5_9_to_tile_4_9_0),
		.out_wire_3_1(vertical_tile_5_9_to_tile_4_9_1),
		.out_wire_3_2(vertical_tile_5_9_to_tile_4_9_2),
		.out_wire_3_3(vertical_tile_5_9_to_tile_4_9_3),
		.in_wire_3_0(vertical_tile_4_9_to_tile_5_9_0),
		.in_wire_3_1(vertical_tile_4_9_to_tile_5_9_1),
		.in_wire_3_2(vertical_tile_4_9_to_tile_5_9_2),
		.in_wire_3_3(vertical_tile_4_9_to_tile_5_9_3),
		.out_wire_1_0(vertical_tile_5_9_to_tile_6_9_0),
		.out_wire_1_1(vertical_tile_5_9_to_tile_6_9_1),
		.out_wire_1_2(vertical_tile_5_9_to_tile_6_9_2),
		.out_wire_1_3(vertical_tile_5_9_to_tile_6_9_3),
		.in_wire_1_0(vertical_tile_6_9_to_tile_5_9_0),
		.in_wire_1_1(vertical_tile_6_9_to_tile_5_9_1),
		.in_wire_1_2(vertical_tile_6_9_to_tile_5_9_2),
		.in_wire_1_3(vertical_tile_6_9_to_tile_5_9_3),
		.out_wire_2_0(horizontal_tile_5_9_to_tile_5_8_0),
		.out_wire_2_1(horizontal_tile_5_9_to_tile_5_8_1),
		.out_wire_2_2(horizontal_tile_5_9_to_tile_5_8_2),
		.out_wire_2_3(horizontal_tile_5_9_to_tile_5_8_3),
		.in_wire_2_0(horizontal_tile_5_8_to_tile_5_9_0),
		.in_wire_2_1(horizontal_tile_5_8_to_tile_5_9_1),
		.in_wire_2_2(horizontal_tile_5_8_to_tile_5_9_2),
		.in_wire_2_3(horizontal_tile_5_8_to_tile_5_9_3),
		.out_wire_0_0(horizontal_tile_5_9_to_tile_5_10_0),
		.out_wire_0_1(horizontal_tile_5_9_to_tile_5_10_1),
		.out_wire_0_2(horizontal_tile_5_9_to_tile_5_10_2),
		.out_wire_0_3(horizontal_tile_5_9_to_tile_5_10_3),
		.in_wire_0_0(horizontal_tile_5_10_to_tile_5_9_0),
		.in_wire_0_1(horizontal_tile_5_10_to_tile_5_9_1),
		.in_wire_0_2(horizontal_tile_5_10_to_tile_5_9_2),
		.in_wire_0_3(horizontal_tile_5_10_to_tile_5_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(170)
	);

	pe_tile pe_tile_5_10(
		.out_wire_3_0(vertical_tile_5_10_to_tile_4_10_0),
		.out_wire_3_1(vertical_tile_5_10_to_tile_4_10_1),
		.out_wire_3_2(vertical_tile_5_10_to_tile_4_10_2),
		.out_wire_3_3(vertical_tile_5_10_to_tile_4_10_3),
		.in_wire_3_0(vertical_tile_4_10_to_tile_5_10_0),
		.in_wire_3_1(vertical_tile_4_10_to_tile_5_10_1),
		.in_wire_3_2(vertical_tile_4_10_to_tile_5_10_2),
		.in_wire_3_3(vertical_tile_4_10_to_tile_5_10_3),
		.out_wire_1_0(vertical_tile_5_10_to_tile_6_10_0),
		.out_wire_1_1(vertical_tile_5_10_to_tile_6_10_1),
		.out_wire_1_2(vertical_tile_5_10_to_tile_6_10_2),
		.out_wire_1_3(vertical_tile_5_10_to_tile_6_10_3),
		.in_wire_1_0(vertical_tile_6_10_to_tile_5_10_0),
		.in_wire_1_1(vertical_tile_6_10_to_tile_5_10_1),
		.in_wire_1_2(vertical_tile_6_10_to_tile_5_10_2),
		.in_wire_1_3(vertical_tile_6_10_to_tile_5_10_3),
		.out_wire_2_0(horizontal_tile_5_10_to_tile_5_9_0),
		.out_wire_2_1(horizontal_tile_5_10_to_tile_5_9_1),
		.out_wire_2_2(horizontal_tile_5_10_to_tile_5_9_2),
		.out_wire_2_3(horizontal_tile_5_10_to_tile_5_9_3),
		.in_wire_2_0(horizontal_tile_5_9_to_tile_5_10_0),
		.in_wire_2_1(horizontal_tile_5_9_to_tile_5_10_1),
		.in_wire_2_2(horizontal_tile_5_9_to_tile_5_10_2),
		.in_wire_2_3(horizontal_tile_5_9_to_tile_5_10_3),
		.out_wire_0_0(horizontal_tile_5_10_to_tile_5_11_0),
		.out_wire_0_1(horizontal_tile_5_10_to_tile_5_11_1),
		.out_wire_0_2(horizontal_tile_5_10_to_tile_5_11_2),
		.out_wire_0_3(horizontal_tile_5_10_to_tile_5_11_3),
		.in_wire_0_0(horizontal_tile_5_11_to_tile_5_10_0),
		.in_wire_0_1(horizontal_tile_5_11_to_tile_5_10_1),
		.in_wire_0_2(horizontal_tile_5_11_to_tile_5_10_2),
		.in_wire_0_3(horizontal_tile_5_11_to_tile_5_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(171)
	);

	pe_tile pe_tile_5_11(
		.out_wire_3_0(vertical_tile_5_11_to_tile_4_11_0),
		.out_wire_3_1(vertical_tile_5_11_to_tile_4_11_1),
		.out_wire_3_2(vertical_tile_5_11_to_tile_4_11_2),
		.out_wire_3_3(vertical_tile_5_11_to_tile_4_11_3),
		.in_wire_3_0(vertical_tile_4_11_to_tile_5_11_0),
		.in_wire_3_1(vertical_tile_4_11_to_tile_5_11_1),
		.in_wire_3_2(vertical_tile_4_11_to_tile_5_11_2),
		.in_wire_3_3(vertical_tile_4_11_to_tile_5_11_3),
		.out_wire_1_0(vertical_tile_5_11_to_tile_6_11_0),
		.out_wire_1_1(vertical_tile_5_11_to_tile_6_11_1),
		.out_wire_1_2(vertical_tile_5_11_to_tile_6_11_2),
		.out_wire_1_3(vertical_tile_5_11_to_tile_6_11_3),
		.in_wire_1_0(vertical_tile_6_11_to_tile_5_11_0),
		.in_wire_1_1(vertical_tile_6_11_to_tile_5_11_1),
		.in_wire_1_2(vertical_tile_6_11_to_tile_5_11_2),
		.in_wire_1_3(vertical_tile_6_11_to_tile_5_11_3),
		.out_wire_2_0(horizontal_tile_5_11_to_tile_5_10_0),
		.out_wire_2_1(horizontal_tile_5_11_to_tile_5_10_1),
		.out_wire_2_2(horizontal_tile_5_11_to_tile_5_10_2),
		.out_wire_2_3(horizontal_tile_5_11_to_tile_5_10_3),
		.in_wire_2_0(horizontal_tile_5_10_to_tile_5_11_0),
		.in_wire_2_1(horizontal_tile_5_10_to_tile_5_11_1),
		.in_wire_2_2(horizontal_tile_5_10_to_tile_5_11_2),
		.in_wire_2_3(horizontal_tile_5_10_to_tile_5_11_3),
		.out_wire_0_0(horizontal_tile_5_11_to_tile_5_12_0),
		.out_wire_0_1(horizontal_tile_5_11_to_tile_5_12_1),
		.out_wire_0_2(horizontal_tile_5_11_to_tile_5_12_2),
		.out_wire_0_3(horizontal_tile_5_11_to_tile_5_12_3),
		.in_wire_0_0(horizontal_tile_5_12_to_tile_5_11_0),
		.in_wire_0_1(horizontal_tile_5_12_to_tile_5_11_1),
		.in_wire_0_2(horizontal_tile_5_12_to_tile_5_11_2),
		.in_wire_0_3(horizontal_tile_5_12_to_tile_5_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(172)
	);

	pe_tile pe_tile_5_12(
		.out_wire_3_0(vertical_tile_5_12_to_tile_4_12_0),
		.out_wire_3_1(vertical_tile_5_12_to_tile_4_12_1),
		.out_wire_3_2(vertical_tile_5_12_to_tile_4_12_2),
		.out_wire_3_3(vertical_tile_5_12_to_tile_4_12_3),
		.in_wire_3_0(vertical_tile_4_12_to_tile_5_12_0),
		.in_wire_3_1(vertical_tile_4_12_to_tile_5_12_1),
		.in_wire_3_2(vertical_tile_4_12_to_tile_5_12_2),
		.in_wire_3_3(vertical_tile_4_12_to_tile_5_12_3),
		.out_wire_1_0(vertical_tile_5_12_to_tile_6_12_0),
		.out_wire_1_1(vertical_tile_5_12_to_tile_6_12_1),
		.out_wire_1_2(vertical_tile_5_12_to_tile_6_12_2),
		.out_wire_1_3(vertical_tile_5_12_to_tile_6_12_3),
		.in_wire_1_0(vertical_tile_6_12_to_tile_5_12_0),
		.in_wire_1_1(vertical_tile_6_12_to_tile_5_12_1),
		.in_wire_1_2(vertical_tile_6_12_to_tile_5_12_2),
		.in_wire_1_3(vertical_tile_6_12_to_tile_5_12_3),
		.out_wire_2_0(horizontal_tile_5_12_to_tile_5_11_0),
		.out_wire_2_1(horizontal_tile_5_12_to_tile_5_11_1),
		.out_wire_2_2(horizontal_tile_5_12_to_tile_5_11_2),
		.out_wire_2_3(horizontal_tile_5_12_to_tile_5_11_3),
		.in_wire_2_0(horizontal_tile_5_11_to_tile_5_12_0),
		.in_wire_2_1(horizontal_tile_5_11_to_tile_5_12_1),
		.in_wire_2_2(horizontal_tile_5_11_to_tile_5_12_2),
		.in_wire_2_3(horizontal_tile_5_11_to_tile_5_12_3),
		.out_wire_0_0(horizontal_tile_5_12_to_tile_5_13_0),
		.out_wire_0_1(horizontal_tile_5_12_to_tile_5_13_1),
		.out_wire_0_2(horizontal_tile_5_12_to_tile_5_13_2),
		.out_wire_0_3(horizontal_tile_5_12_to_tile_5_13_3),
		.in_wire_0_0(horizontal_tile_5_13_to_tile_5_12_0),
		.in_wire_0_1(horizontal_tile_5_13_to_tile_5_12_1),
		.in_wire_0_2(horizontal_tile_5_13_to_tile_5_12_2),
		.in_wire_0_3(horizontal_tile_5_13_to_tile_5_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(173)
	);

	pe_tile pe_tile_5_13(
		.out_wire_3_0(vertical_tile_5_13_to_tile_4_13_0),
		.out_wire_3_1(vertical_tile_5_13_to_tile_4_13_1),
		.out_wire_3_2(vertical_tile_5_13_to_tile_4_13_2),
		.out_wire_3_3(vertical_tile_5_13_to_tile_4_13_3),
		.in_wire_3_0(vertical_tile_4_13_to_tile_5_13_0),
		.in_wire_3_1(vertical_tile_4_13_to_tile_5_13_1),
		.in_wire_3_2(vertical_tile_4_13_to_tile_5_13_2),
		.in_wire_3_3(vertical_tile_4_13_to_tile_5_13_3),
		.out_wire_1_0(vertical_tile_5_13_to_tile_6_13_0),
		.out_wire_1_1(vertical_tile_5_13_to_tile_6_13_1),
		.out_wire_1_2(vertical_tile_5_13_to_tile_6_13_2),
		.out_wire_1_3(vertical_tile_5_13_to_tile_6_13_3),
		.in_wire_1_0(vertical_tile_6_13_to_tile_5_13_0),
		.in_wire_1_1(vertical_tile_6_13_to_tile_5_13_1),
		.in_wire_1_2(vertical_tile_6_13_to_tile_5_13_2),
		.in_wire_1_3(vertical_tile_6_13_to_tile_5_13_3),
		.out_wire_2_0(horizontal_tile_5_13_to_tile_5_12_0),
		.out_wire_2_1(horizontal_tile_5_13_to_tile_5_12_1),
		.out_wire_2_2(horizontal_tile_5_13_to_tile_5_12_2),
		.out_wire_2_3(horizontal_tile_5_13_to_tile_5_12_3),
		.in_wire_2_0(horizontal_tile_5_12_to_tile_5_13_0),
		.in_wire_2_1(horizontal_tile_5_12_to_tile_5_13_1),
		.in_wire_2_2(horizontal_tile_5_12_to_tile_5_13_2),
		.in_wire_2_3(horizontal_tile_5_12_to_tile_5_13_3),
		.out_wire_0_0(horizontal_tile_5_13_to_tile_5_14_0),
		.out_wire_0_1(horizontal_tile_5_13_to_tile_5_14_1),
		.out_wire_0_2(horizontal_tile_5_13_to_tile_5_14_2),
		.out_wire_0_3(horizontal_tile_5_13_to_tile_5_14_3),
		.in_wire_0_0(horizontal_tile_5_14_to_tile_5_13_0),
		.in_wire_0_1(horizontal_tile_5_14_to_tile_5_13_1),
		.in_wire_0_2(horizontal_tile_5_14_to_tile_5_13_2),
		.in_wire_0_3(horizontal_tile_5_14_to_tile_5_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(174)
	);

	pe_tile pe_tile_5_14(
		.out_wire_3_0(vertical_tile_5_14_to_tile_4_14_0),
		.out_wire_3_1(vertical_tile_5_14_to_tile_4_14_1),
		.out_wire_3_2(vertical_tile_5_14_to_tile_4_14_2),
		.out_wire_3_3(vertical_tile_5_14_to_tile_4_14_3),
		.in_wire_3_0(vertical_tile_4_14_to_tile_5_14_0),
		.in_wire_3_1(vertical_tile_4_14_to_tile_5_14_1),
		.in_wire_3_2(vertical_tile_4_14_to_tile_5_14_2),
		.in_wire_3_3(vertical_tile_4_14_to_tile_5_14_3),
		.out_wire_1_0(vertical_tile_5_14_to_tile_6_14_0),
		.out_wire_1_1(vertical_tile_5_14_to_tile_6_14_1),
		.out_wire_1_2(vertical_tile_5_14_to_tile_6_14_2),
		.out_wire_1_3(vertical_tile_5_14_to_tile_6_14_3),
		.in_wire_1_0(vertical_tile_6_14_to_tile_5_14_0),
		.in_wire_1_1(vertical_tile_6_14_to_tile_5_14_1),
		.in_wire_1_2(vertical_tile_6_14_to_tile_5_14_2),
		.in_wire_1_3(vertical_tile_6_14_to_tile_5_14_3),
		.out_wire_2_0(horizontal_tile_5_14_to_tile_5_13_0),
		.out_wire_2_1(horizontal_tile_5_14_to_tile_5_13_1),
		.out_wire_2_2(horizontal_tile_5_14_to_tile_5_13_2),
		.out_wire_2_3(horizontal_tile_5_14_to_tile_5_13_3),
		.in_wire_2_0(horizontal_tile_5_13_to_tile_5_14_0),
		.in_wire_2_1(horizontal_tile_5_13_to_tile_5_14_1),
		.in_wire_2_2(horizontal_tile_5_13_to_tile_5_14_2),
		.in_wire_2_3(horizontal_tile_5_13_to_tile_5_14_3),
		.out_wire_0_0(horizontal_tile_5_14_to_tile_5_15_0),
		.out_wire_0_1(horizontal_tile_5_14_to_tile_5_15_1),
		.out_wire_0_2(horizontal_tile_5_14_to_tile_5_15_2),
		.out_wire_0_3(horizontal_tile_5_14_to_tile_5_15_3),
		.in_wire_0_0(horizontal_tile_5_15_to_tile_5_14_0),
		.in_wire_0_1(horizontal_tile_5_15_to_tile_5_14_1),
		.in_wire_0_2(horizontal_tile_5_15_to_tile_5_14_2),
		.in_wire_0_3(horizontal_tile_5_15_to_tile_5_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(175)
	);

	pe_tile pe_tile_5_15(
		.out_wire_3_0(vertical_tile_5_15_to_tile_4_15_0),
		.out_wire_3_1(vertical_tile_5_15_to_tile_4_15_1),
		.out_wire_3_2(vertical_tile_5_15_to_tile_4_15_2),
		.out_wire_3_3(vertical_tile_5_15_to_tile_4_15_3),
		.in_wire_3_0(vertical_tile_4_15_to_tile_5_15_0),
		.in_wire_3_1(vertical_tile_4_15_to_tile_5_15_1),
		.in_wire_3_2(vertical_tile_4_15_to_tile_5_15_2),
		.in_wire_3_3(vertical_tile_4_15_to_tile_5_15_3),
		.out_wire_1_0(vertical_tile_5_15_to_tile_6_15_0),
		.out_wire_1_1(vertical_tile_5_15_to_tile_6_15_1),
		.out_wire_1_2(vertical_tile_5_15_to_tile_6_15_2),
		.out_wire_1_3(vertical_tile_5_15_to_tile_6_15_3),
		.in_wire_1_0(vertical_tile_6_15_to_tile_5_15_0),
		.in_wire_1_1(vertical_tile_6_15_to_tile_5_15_1),
		.in_wire_1_2(vertical_tile_6_15_to_tile_5_15_2),
		.in_wire_1_3(vertical_tile_6_15_to_tile_5_15_3),
		.out_wire_2_0(horizontal_tile_5_15_to_tile_5_14_0),
		.out_wire_2_1(horizontal_tile_5_15_to_tile_5_14_1),
		.out_wire_2_2(horizontal_tile_5_15_to_tile_5_14_2),
		.out_wire_2_3(horizontal_tile_5_15_to_tile_5_14_3),
		.in_wire_2_0(horizontal_tile_5_14_to_tile_5_15_0),
		.in_wire_2_1(horizontal_tile_5_14_to_tile_5_15_1),
		.in_wire_2_2(horizontal_tile_5_14_to_tile_5_15_2),
		.in_wire_2_3(horizontal_tile_5_14_to_tile_5_15_3),
		.out_wire_0_0(horizontal_tile_5_15_to_tile_5_16_0),
		.out_wire_0_1(horizontal_tile_5_15_to_tile_5_16_1),
		.out_wire_0_2(horizontal_tile_5_15_to_tile_5_16_2),
		.out_wire_0_3(horizontal_tile_5_15_to_tile_5_16_3),
		.in_wire_0_0(horizontal_tile_5_16_to_tile_5_15_0),
		.in_wire_0_1(horizontal_tile_5_16_to_tile_5_15_1),
		.in_wire_0_2(horizontal_tile_5_16_to_tile_5_15_2),
		.in_wire_0_3(horizontal_tile_5_16_to_tile_5_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(176)
	);

	pe_tile pe_tile_5_16(
		.out_wire_3_0(vertical_tile_5_16_to_tile_4_16_0),
		.out_wire_3_1(vertical_tile_5_16_to_tile_4_16_1),
		.out_wire_3_2(vertical_tile_5_16_to_tile_4_16_2),
		.out_wire_3_3(vertical_tile_5_16_to_tile_4_16_3),
		.in_wire_3_0(vertical_tile_4_16_to_tile_5_16_0),
		.in_wire_3_1(vertical_tile_4_16_to_tile_5_16_1),
		.in_wire_3_2(vertical_tile_4_16_to_tile_5_16_2),
		.in_wire_3_3(vertical_tile_4_16_to_tile_5_16_3),
		.out_wire_1_0(vertical_tile_5_16_to_tile_6_16_0),
		.out_wire_1_1(vertical_tile_5_16_to_tile_6_16_1),
		.out_wire_1_2(vertical_tile_5_16_to_tile_6_16_2),
		.out_wire_1_3(vertical_tile_5_16_to_tile_6_16_3),
		.in_wire_1_0(vertical_tile_6_16_to_tile_5_16_0),
		.in_wire_1_1(vertical_tile_6_16_to_tile_5_16_1),
		.in_wire_1_2(vertical_tile_6_16_to_tile_5_16_2),
		.in_wire_1_3(vertical_tile_6_16_to_tile_5_16_3),
		.out_wire_2_0(horizontal_tile_5_16_to_tile_5_15_0),
		.out_wire_2_1(horizontal_tile_5_16_to_tile_5_15_1),
		.out_wire_2_2(horizontal_tile_5_16_to_tile_5_15_2),
		.out_wire_2_3(horizontal_tile_5_16_to_tile_5_15_3),
		.in_wire_2_0(horizontal_tile_5_15_to_tile_5_16_0),
		.in_wire_2_1(horizontal_tile_5_15_to_tile_5_16_1),
		.in_wire_2_2(horizontal_tile_5_15_to_tile_5_16_2),
		.in_wire_2_3(horizontal_tile_5_15_to_tile_5_16_3),
		.out_wire_0_0(horizontal_tile_5_16_to_tile_5_17_0),
		.out_wire_0_1(horizontal_tile_5_16_to_tile_5_17_1),
		.out_wire_0_2(horizontal_tile_5_16_to_tile_5_17_2),
		.out_wire_0_3(horizontal_tile_5_16_to_tile_5_17_3),
		.in_wire_0_0(horizontal_tile_5_17_to_tile_5_16_0),
		.in_wire_0_1(horizontal_tile_5_17_to_tile_5_16_1),
		.in_wire_0_2(horizontal_tile_5_17_to_tile_5_16_2),
		.in_wire_0_3(horizontal_tile_5_17_to_tile_5_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(177)
	);

	pe_tile pe_tile_5_17(
		.out_wire_3_0(vertical_tile_5_17_to_tile_4_17_0),
		.out_wire_3_1(vertical_tile_5_17_to_tile_4_17_1),
		.out_wire_3_2(vertical_tile_5_17_to_tile_4_17_2),
		.out_wire_3_3(vertical_tile_5_17_to_tile_4_17_3),
		.in_wire_3_0(vertical_tile_4_17_to_tile_5_17_0),
		.in_wire_3_1(vertical_tile_4_17_to_tile_5_17_1),
		.in_wire_3_2(vertical_tile_4_17_to_tile_5_17_2),
		.in_wire_3_3(vertical_tile_4_17_to_tile_5_17_3),
		.out_wire_1_0(vertical_tile_5_17_to_tile_6_17_0),
		.out_wire_1_1(vertical_tile_5_17_to_tile_6_17_1),
		.out_wire_1_2(vertical_tile_5_17_to_tile_6_17_2),
		.out_wire_1_3(vertical_tile_5_17_to_tile_6_17_3),
		.in_wire_1_0(vertical_tile_6_17_to_tile_5_17_0),
		.in_wire_1_1(vertical_tile_6_17_to_tile_5_17_1),
		.in_wire_1_2(vertical_tile_6_17_to_tile_5_17_2),
		.in_wire_1_3(vertical_tile_6_17_to_tile_5_17_3),
		.out_wire_2_0(horizontal_tile_5_17_to_tile_5_16_0),
		.out_wire_2_1(horizontal_tile_5_17_to_tile_5_16_1),
		.out_wire_2_2(horizontal_tile_5_17_to_tile_5_16_2),
		.out_wire_2_3(horizontal_tile_5_17_to_tile_5_16_3),
		.in_wire_2_0(horizontal_tile_5_16_to_tile_5_17_0),
		.in_wire_2_1(horizontal_tile_5_16_to_tile_5_17_1),
		.in_wire_2_2(horizontal_tile_5_16_to_tile_5_17_2),
		.in_wire_2_3(horizontal_tile_5_16_to_tile_5_17_3),
		.out_wire_0_0(horizontal_tile_5_17_to_tile_5_18_0),
		.out_wire_0_1(horizontal_tile_5_17_to_tile_5_18_1),
		.out_wire_0_2(horizontal_tile_5_17_to_tile_5_18_2),
		.out_wire_0_3(horizontal_tile_5_17_to_tile_5_18_3),
		.in_wire_0_0(horizontal_tile_5_18_to_tile_5_17_0),
		.in_wire_0_1(horizontal_tile_5_18_to_tile_5_17_1),
		.in_wire_0_2(horizontal_tile_5_18_to_tile_5_17_2),
		.in_wire_0_3(horizontal_tile_5_18_to_tile_5_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(178)
	);

	pe_tile pe_tile_5_18(
		.out_wire_3_0(vertical_tile_5_18_to_tile_4_18_0),
		.out_wire_3_1(vertical_tile_5_18_to_tile_4_18_1),
		.out_wire_3_2(vertical_tile_5_18_to_tile_4_18_2),
		.out_wire_3_3(vertical_tile_5_18_to_tile_4_18_3),
		.in_wire_3_0(vertical_tile_4_18_to_tile_5_18_0),
		.in_wire_3_1(vertical_tile_4_18_to_tile_5_18_1),
		.in_wire_3_2(vertical_tile_4_18_to_tile_5_18_2),
		.in_wire_3_3(vertical_tile_4_18_to_tile_5_18_3),
		.out_wire_1_0(vertical_tile_5_18_to_tile_6_18_0),
		.out_wire_1_1(vertical_tile_5_18_to_tile_6_18_1),
		.out_wire_1_2(vertical_tile_5_18_to_tile_6_18_2),
		.out_wire_1_3(vertical_tile_5_18_to_tile_6_18_3),
		.in_wire_1_0(vertical_tile_6_18_to_tile_5_18_0),
		.in_wire_1_1(vertical_tile_6_18_to_tile_5_18_1),
		.in_wire_1_2(vertical_tile_6_18_to_tile_5_18_2),
		.in_wire_1_3(vertical_tile_6_18_to_tile_5_18_3),
		.out_wire_2_0(horizontal_tile_5_18_to_tile_5_17_0),
		.out_wire_2_1(horizontal_tile_5_18_to_tile_5_17_1),
		.out_wire_2_2(horizontal_tile_5_18_to_tile_5_17_2),
		.out_wire_2_3(horizontal_tile_5_18_to_tile_5_17_3),
		.in_wire_2_0(horizontal_tile_5_17_to_tile_5_18_0),
		.in_wire_2_1(horizontal_tile_5_17_to_tile_5_18_1),
		.in_wire_2_2(horizontal_tile_5_17_to_tile_5_18_2),
		.in_wire_2_3(horizontal_tile_5_17_to_tile_5_18_3),
		.out_wire_0_0(horizontal_tile_5_18_to_tile_5_19_0),
		.out_wire_0_1(horizontal_tile_5_18_to_tile_5_19_1),
		.out_wire_0_2(horizontal_tile_5_18_to_tile_5_19_2),
		.out_wire_0_3(horizontal_tile_5_18_to_tile_5_19_3),
		.in_wire_0_0(horizontal_tile_5_19_to_tile_5_18_0),
		.in_wire_0_1(horizontal_tile_5_19_to_tile_5_18_1),
		.in_wire_0_2(horizontal_tile_5_19_to_tile_5_18_2),
		.in_wire_0_3(horizontal_tile_5_19_to_tile_5_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(179)
	);

	pe_tile pe_tile_5_19(
		.out_wire_3_0(vertical_tile_5_19_to_tile_4_19_0),
		.out_wire_3_1(vertical_tile_5_19_to_tile_4_19_1),
		.out_wire_3_2(vertical_tile_5_19_to_tile_4_19_2),
		.out_wire_3_3(vertical_tile_5_19_to_tile_4_19_3),
		.in_wire_3_0(vertical_tile_4_19_to_tile_5_19_0),
		.in_wire_3_1(vertical_tile_4_19_to_tile_5_19_1),
		.in_wire_3_2(vertical_tile_4_19_to_tile_5_19_2),
		.in_wire_3_3(vertical_tile_4_19_to_tile_5_19_3),
		.out_wire_1_0(vertical_tile_5_19_to_tile_6_19_0),
		.out_wire_1_1(vertical_tile_5_19_to_tile_6_19_1),
		.out_wire_1_2(vertical_tile_5_19_to_tile_6_19_2),
		.out_wire_1_3(vertical_tile_5_19_to_tile_6_19_3),
		.in_wire_1_0(vertical_tile_6_19_to_tile_5_19_0),
		.in_wire_1_1(vertical_tile_6_19_to_tile_5_19_1),
		.in_wire_1_2(vertical_tile_6_19_to_tile_5_19_2),
		.in_wire_1_3(vertical_tile_6_19_to_tile_5_19_3),
		.out_wire_2_0(horizontal_tile_5_19_to_tile_5_18_0),
		.out_wire_2_1(horizontal_tile_5_19_to_tile_5_18_1),
		.out_wire_2_2(horizontal_tile_5_19_to_tile_5_18_2),
		.out_wire_2_3(horizontal_tile_5_19_to_tile_5_18_3),
		.in_wire_2_0(horizontal_tile_5_18_to_tile_5_19_0),
		.in_wire_2_1(horizontal_tile_5_18_to_tile_5_19_1),
		.in_wire_2_2(horizontal_tile_5_18_to_tile_5_19_2),
		.in_wire_2_3(horizontal_tile_5_18_to_tile_5_19_3),
		.out_wire_0_0(horizontal_tile_5_19_to_tile_5_20_0),
		.out_wire_0_1(horizontal_tile_5_19_to_tile_5_20_1),
		.out_wire_0_2(horizontal_tile_5_19_to_tile_5_20_2),
		.out_wire_0_3(horizontal_tile_5_19_to_tile_5_20_3),
		.in_wire_0_0(horizontal_tile_5_20_to_tile_5_19_0),
		.in_wire_0_1(horizontal_tile_5_20_to_tile_5_19_1),
		.in_wire_0_2(horizontal_tile_5_20_to_tile_5_19_2),
		.in_wire_0_3(horizontal_tile_5_20_to_tile_5_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(180)
	);

	pe_tile pe_tile_5_20(
		.out_wire_3_0(vertical_tile_5_20_to_tile_4_20_0),
		.out_wire_3_1(vertical_tile_5_20_to_tile_4_20_1),
		.out_wire_3_2(vertical_tile_5_20_to_tile_4_20_2),
		.out_wire_3_3(vertical_tile_5_20_to_tile_4_20_3),
		.in_wire_3_0(vertical_tile_4_20_to_tile_5_20_0),
		.in_wire_3_1(vertical_tile_4_20_to_tile_5_20_1),
		.in_wire_3_2(vertical_tile_4_20_to_tile_5_20_2),
		.in_wire_3_3(vertical_tile_4_20_to_tile_5_20_3),
		.out_wire_1_0(vertical_tile_5_20_to_tile_6_20_0),
		.out_wire_1_1(vertical_tile_5_20_to_tile_6_20_1),
		.out_wire_1_2(vertical_tile_5_20_to_tile_6_20_2),
		.out_wire_1_3(vertical_tile_5_20_to_tile_6_20_3),
		.in_wire_1_0(vertical_tile_6_20_to_tile_5_20_0),
		.in_wire_1_1(vertical_tile_6_20_to_tile_5_20_1),
		.in_wire_1_2(vertical_tile_6_20_to_tile_5_20_2),
		.in_wire_1_3(vertical_tile_6_20_to_tile_5_20_3),
		.out_wire_2_0(horizontal_tile_5_20_to_tile_5_19_0),
		.out_wire_2_1(horizontal_tile_5_20_to_tile_5_19_1),
		.out_wire_2_2(horizontal_tile_5_20_to_tile_5_19_2),
		.out_wire_2_3(horizontal_tile_5_20_to_tile_5_19_3),
		.in_wire_2_0(horizontal_tile_5_19_to_tile_5_20_0),
		.in_wire_2_1(horizontal_tile_5_19_to_tile_5_20_1),
		.in_wire_2_2(horizontal_tile_5_19_to_tile_5_20_2),
		.in_wire_2_3(horizontal_tile_5_19_to_tile_5_20_3),
		.out_wire_0_0(horizontal_tile_5_20_to_tile_5_21_0),
		.out_wire_0_1(horizontal_tile_5_20_to_tile_5_21_1),
		.out_wire_0_2(horizontal_tile_5_20_to_tile_5_21_2),
		.out_wire_0_3(horizontal_tile_5_20_to_tile_5_21_3),
		.in_wire_0_0(horizontal_tile_5_21_to_tile_5_20_0),
		.in_wire_0_1(horizontal_tile_5_21_to_tile_5_20_1),
		.in_wire_0_2(horizontal_tile_5_21_to_tile_5_20_2),
		.in_wire_0_3(horizontal_tile_5_21_to_tile_5_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(181)
	);

	pe_tile pe_tile_5_21(
		.out_wire_3_0(vertical_tile_5_21_to_tile_4_21_0),
		.out_wire_3_1(vertical_tile_5_21_to_tile_4_21_1),
		.out_wire_3_2(vertical_tile_5_21_to_tile_4_21_2),
		.out_wire_3_3(vertical_tile_5_21_to_tile_4_21_3),
		.in_wire_3_0(vertical_tile_4_21_to_tile_5_21_0),
		.in_wire_3_1(vertical_tile_4_21_to_tile_5_21_1),
		.in_wire_3_2(vertical_tile_4_21_to_tile_5_21_2),
		.in_wire_3_3(vertical_tile_4_21_to_tile_5_21_3),
		.out_wire_1_0(vertical_tile_5_21_to_tile_6_21_0),
		.out_wire_1_1(vertical_tile_5_21_to_tile_6_21_1),
		.out_wire_1_2(vertical_tile_5_21_to_tile_6_21_2),
		.out_wire_1_3(vertical_tile_5_21_to_tile_6_21_3),
		.in_wire_1_0(vertical_tile_6_21_to_tile_5_21_0),
		.in_wire_1_1(vertical_tile_6_21_to_tile_5_21_1),
		.in_wire_1_2(vertical_tile_6_21_to_tile_5_21_2),
		.in_wire_1_3(vertical_tile_6_21_to_tile_5_21_3),
		.out_wire_2_0(horizontal_tile_5_21_to_tile_5_20_0),
		.out_wire_2_1(horizontal_tile_5_21_to_tile_5_20_1),
		.out_wire_2_2(horizontal_tile_5_21_to_tile_5_20_2),
		.out_wire_2_3(horizontal_tile_5_21_to_tile_5_20_3),
		.in_wire_2_0(horizontal_tile_5_20_to_tile_5_21_0),
		.in_wire_2_1(horizontal_tile_5_20_to_tile_5_21_1),
		.in_wire_2_2(horizontal_tile_5_20_to_tile_5_21_2),
		.in_wire_2_3(horizontal_tile_5_20_to_tile_5_21_3),
		.out_wire_0_0(horizontal_tile_5_21_to_tile_5_22_0),
		.out_wire_0_1(horizontal_tile_5_21_to_tile_5_22_1),
		.out_wire_0_2(horizontal_tile_5_21_to_tile_5_22_2),
		.out_wire_0_3(horizontal_tile_5_21_to_tile_5_22_3),
		.in_wire_0_0(horizontal_tile_5_22_to_tile_5_21_0),
		.in_wire_0_1(horizontal_tile_5_22_to_tile_5_21_1),
		.in_wire_0_2(horizontal_tile_5_22_to_tile_5_21_2),
		.in_wire_0_3(horizontal_tile_5_22_to_tile_5_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(182)
	);

	pe_tile pe_tile_5_22(
		.out_wire_3_0(vertical_tile_5_22_to_tile_4_22_0),
		.out_wire_3_1(vertical_tile_5_22_to_tile_4_22_1),
		.out_wire_3_2(vertical_tile_5_22_to_tile_4_22_2),
		.out_wire_3_3(vertical_tile_5_22_to_tile_4_22_3),
		.in_wire_3_0(vertical_tile_4_22_to_tile_5_22_0),
		.in_wire_3_1(vertical_tile_4_22_to_tile_5_22_1),
		.in_wire_3_2(vertical_tile_4_22_to_tile_5_22_2),
		.in_wire_3_3(vertical_tile_4_22_to_tile_5_22_3),
		.out_wire_1_0(vertical_tile_5_22_to_tile_6_22_0),
		.out_wire_1_1(vertical_tile_5_22_to_tile_6_22_1),
		.out_wire_1_2(vertical_tile_5_22_to_tile_6_22_2),
		.out_wire_1_3(vertical_tile_5_22_to_tile_6_22_3),
		.in_wire_1_0(vertical_tile_6_22_to_tile_5_22_0),
		.in_wire_1_1(vertical_tile_6_22_to_tile_5_22_1),
		.in_wire_1_2(vertical_tile_6_22_to_tile_5_22_2),
		.in_wire_1_3(vertical_tile_6_22_to_tile_5_22_3),
		.out_wire_2_0(horizontal_tile_5_22_to_tile_5_21_0),
		.out_wire_2_1(horizontal_tile_5_22_to_tile_5_21_1),
		.out_wire_2_2(horizontal_tile_5_22_to_tile_5_21_2),
		.out_wire_2_3(horizontal_tile_5_22_to_tile_5_21_3),
		.in_wire_2_0(horizontal_tile_5_21_to_tile_5_22_0),
		.in_wire_2_1(horizontal_tile_5_21_to_tile_5_22_1),
		.in_wire_2_2(horizontal_tile_5_21_to_tile_5_22_2),
		.in_wire_2_3(horizontal_tile_5_21_to_tile_5_22_3),
		.out_wire_0_0(horizontal_tile_5_22_to_tile_5_23_0),
		.out_wire_0_1(horizontal_tile_5_22_to_tile_5_23_1),
		.out_wire_0_2(horizontal_tile_5_22_to_tile_5_23_2),
		.out_wire_0_3(horizontal_tile_5_22_to_tile_5_23_3),
		.in_wire_0_0(horizontal_tile_5_23_to_tile_5_22_0),
		.in_wire_0_1(horizontal_tile_5_23_to_tile_5_22_1),
		.in_wire_0_2(horizontal_tile_5_23_to_tile_5_22_2),
		.in_wire_0_3(horizontal_tile_5_23_to_tile_5_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(183)
	);

	pe_tile pe_tile_5_23(
		.out_wire_3_0(vertical_tile_5_23_to_tile_4_23_0),
		.out_wire_3_1(vertical_tile_5_23_to_tile_4_23_1),
		.out_wire_3_2(vertical_tile_5_23_to_tile_4_23_2),
		.out_wire_3_3(vertical_tile_5_23_to_tile_4_23_3),
		.in_wire_3_0(vertical_tile_4_23_to_tile_5_23_0),
		.in_wire_3_1(vertical_tile_4_23_to_tile_5_23_1),
		.in_wire_3_2(vertical_tile_4_23_to_tile_5_23_2),
		.in_wire_3_3(vertical_tile_4_23_to_tile_5_23_3),
		.out_wire_1_0(vertical_tile_5_23_to_tile_6_23_0),
		.out_wire_1_1(vertical_tile_5_23_to_tile_6_23_1),
		.out_wire_1_2(vertical_tile_5_23_to_tile_6_23_2),
		.out_wire_1_3(vertical_tile_5_23_to_tile_6_23_3),
		.in_wire_1_0(vertical_tile_6_23_to_tile_5_23_0),
		.in_wire_1_1(vertical_tile_6_23_to_tile_5_23_1),
		.in_wire_1_2(vertical_tile_6_23_to_tile_5_23_2),
		.in_wire_1_3(vertical_tile_6_23_to_tile_5_23_3),
		.out_wire_2_0(horizontal_tile_5_23_to_tile_5_22_0),
		.out_wire_2_1(horizontal_tile_5_23_to_tile_5_22_1),
		.out_wire_2_2(horizontal_tile_5_23_to_tile_5_22_2),
		.out_wire_2_3(horizontal_tile_5_23_to_tile_5_22_3),
		.in_wire_2_0(horizontal_tile_5_22_to_tile_5_23_0),
		.in_wire_2_1(horizontal_tile_5_22_to_tile_5_23_1),
		.in_wire_2_2(horizontal_tile_5_22_to_tile_5_23_2),
		.in_wire_2_3(horizontal_tile_5_22_to_tile_5_23_3),
		.out_wire_0_0(horizontal_tile_5_23_to_tile_5_24_0),
		.out_wire_0_1(horizontal_tile_5_23_to_tile_5_24_1),
		.out_wire_0_2(horizontal_tile_5_23_to_tile_5_24_2),
		.out_wire_0_3(horizontal_tile_5_23_to_tile_5_24_3),
		.in_wire_0_0(horizontal_tile_5_24_to_tile_5_23_0),
		.in_wire_0_1(horizontal_tile_5_24_to_tile_5_23_1),
		.in_wire_0_2(horizontal_tile_5_24_to_tile_5_23_2),
		.in_wire_0_3(horizontal_tile_5_24_to_tile_5_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(184)
	);

	pe_tile pe_tile_5_24(
		.out_wire_3_0(vertical_tile_5_24_to_tile_4_24_0),
		.out_wire_3_1(vertical_tile_5_24_to_tile_4_24_1),
		.out_wire_3_2(vertical_tile_5_24_to_tile_4_24_2),
		.out_wire_3_3(vertical_tile_5_24_to_tile_4_24_3),
		.in_wire_3_0(vertical_tile_4_24_to_tile_5_24_0),
		.in_wire_3_1(vertical_tile_4_24_to_tile_5_24_1),
		.in_wire_3_2(vertical_tile_4_24_to_tile_5_24_2),
		.in_wire_3_3(vertical_tile_4_24_to_tile_5_24_3),
		.out_wire_1_0(vertical_tile_5_24_to_tile_6_24_0),
		.out_wire_1_1(vertical_tile_5_24_to_tile_6_24_1),
		.out_wire_1_2(vertical_tile_5_24_to_tile_6_24_2),
		.out_wire_1_3(vertical_tile_5_24_to_tile_6_24_3),
		.in_wire_1_0(vertical_tile_6_24_to_tile_5_24_0),
		.in_wire_1_1(vertical_tile_6_24_to_tile_5_24_1),
		.in_wire_1_2(vertical_tile_6_24_to_tile_5_24_2),
		.in_wire_1_3(vertical_tile_6_24_to_tile_5_24_3),
		.out_wire_2_0(horizontal_tile_5_24_to_tile_5_23_0),
		.out_wire_2_1(horizontal_tile_5_24_to_tile_5_23_1),
		.out_wire_2_2(horizontal_tile_5_24_to_tile_5_23_2),
		.out_wire_2_3(horizontal_tile_5_24_to_tile_5_23_3),
		.in_wire_2_0(horizontal_tile_5_23_to_tile_5_24_0),
		.in_wire_2_1(horizontal_tile_5_23_to_tile_5_24_1),
		.in_wire_2_2(horizontal_tile_5_23_to_tile_5_24_2),
		.in_wire_2_3(horizontal_tile_5_23_to_tile_5_24_3),
		.out_wire_0_0(horizontal_tile_5_24_to_tile_5_25_0),
		.out_wire_0_1(horizontal_tile_5_24_to_tile_5_25_1),
		.out_wire_0_2(horizontal_tile_5_24_to_tile_5_25_2),
		.out_wire_0_3(horizontal_tile_5_24_to_tile_5_25_3),
		.in_wire_0_0(horizontal_tile_5_25_to_tile_5_24_0),
		.in_wire_0_1(horizontal_tile_5_25_to_tile_5_24_1),
		.in_wire_0_2(horizontal_tile_5_25_to_tile_5_24_2),
		.in_wire_0_3(horizontal_tile_5_25_to_tile_5_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(185)
	);

	pe_tile pe_tile_5_25(
		.out_wire_3_0(vertical_tile_5_25_to_tile_4_25_0),
		.out_wire_3_1(vertical_tile_5_25_to_tile_4_25_1),
		.out_wire_3_2(vertical_tile_5_25_to_tile_4_25_2),
		.out_wire_3_3(vertical_tile_5_25_to_tile_4_25_3),
		.in_wire_3_0(vertical_tile_4_25_to_tile_5_25_0),
		.in_wire_3_1(vertical_tile_4_25_to_tile_5_25_1),
		.in_wire_3_2(vertical_tile_4_25_to_tile_5_25_2),
		.in_wire_3_3(vertical_tile_4_25_to_tile_5_25_3),
		.out_wire_1_0(vertical_tile_5_25_to_tile_6_25_0),
		.out_wire_1_1(vertical_tile_5_25_to_tile_6_25_1),
		.out_wire_1_2(vertical_tile_5_25_to_tile_6_25_2),
		.out_wire_1_3(vertical_tile_5_25_to_tile_6_25_3),
		.in_wire_1_0(vertical_tile_6_25_to_tile_5_25_0),
		.in_wire_1_1(vertical_tile_6_25_to_tile_5_25_1),
		.in_wire_1_2(vertical_tile_6_25_to_tile_5_25_2),
		.in_wire_1_3(vertical_tile_6_25_to_tile_5_25_3),
		.out_wire_2_0(horizontal_tile_5_25_to_tile_5_24_0),
		.out_wire_2_1(horizontal_tile_5_25_to_tile_5_24_1),
		.out_wire_2_2(horizontal_tile_5_25_to_tile_5_24_2),
		.out_wire_2_3(horizontal_tile_5_25_to_tile_5_24_3),
		.in_wire_2_0(horizontal_tile_5_24_to_tile_5_25_0),
		.in_wire_2_1(horizontal_tile_5_24_to_tile_5_25_1),
		.in_wire_2_2(horizontal_tile_5_24_to_tile_5_25_2),
		.in_wire_2_3(horizontal_tile_5_24_to_tile_5_25_3),
		.out_wire_0_0(horizontal_tile_5_25_to_tile_5_26_0),
		.out_wire_0_1(horizontal_tile_5_25_to_tile_5_26_1),
		.out_wire_0_2(horizontal_tile_5_25_to_tile_5_26_2),
		.out_wire_0_3(horizontal_tile_5_25_to_tile_5_26_3),
		.in_wire_0_0(horizontal_tile_5_26_to_tile_5_25_0),
		.in_wire_0_1(horizontal_tile_5_26_to_tile_5_25_1),
		.in_wire_0_2(horizontal_tile_5_26_to_tile_5_25_2),
		.in_wire_0_3(horizontal_tile_5_26_to_tile_5_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(186)
	);

	pe_tile pe_tile_5_26(
		.out_wire_3_0(vertical_tile_5_26_to_tile_4_26_0),
		.out_wire_3_1(vertical_tile_5_26_to_tile_4_26_1),
		.out_wire_3_2(vertical_tile_5_26_to_tile_4_26_2),
		.out_wire_3_3(vertical_tile_5_26_to_tile_4_26_3),
		.in_wire_3_0(vertical_tile_4_26_to_tile_5_26_0),
		.in_wire_3_1(vertical_tile_4_26_to_tile_5_26_1),
		.in_wire_3_2(vertical_tile_4_26_to_tile_5_26_2),
		.in_wire_3_3(vertical_tile_4_26_to_tile_5_26_3),
		.out_wire_1_0(vertical_tile_5_26_to_tile_6_26_0),
		.out_wire_1_1(vertical_tile_5_26_to_tile_6_26_1),
		.out_wire_1_2(vertical_tile_5_26_to_tile_6_26_2),
		.out_wire_1_3(vertical_tile_5_26_to_tile_6_26_3),
		.in_wire_1_0(vertical_tile_6_26_to_tile_5_26_0),
		.in_wire_1_1(vertical_tile_6_26_to_tile_5_26_1),
		.in_wire_1_2(vertical_tile_6_26_to_tile_5_26_2),
		.in_wire_1_3(vertical_tile_6_26_to_tile_5_26_3),
		.out_wire_2_0(horizontal_tile_5_26_to_tile_5_25_0),
		.out_wire_2_1(horizontal_tile_5_26_to_tile_5_25_1),
		.out_wire_2_2(horizontal_tile_5_26_to_tile_5_25_2),
		.out_wire_2_3(horizontal_tile_5_26_to_tile_5_25_3),
		.in_wire_2_0(horizontal_tile_5_25_to_tile_5_26_0),
		.in_wire_2_1(horizontal_tile_5_25_to_tile_5_26_1),
		.in_wire_2_2(horizontal_tile_5_25_to_tile_5_26_2),
		.in_wire_2_3(horizontal_tile_5_25_to_tile_5_26_3),
		.out_wire_0_0(horizontal_tile_5_26_to_tile_5_27_0),
		.out_wire_0_1(horizontal_tile_5_26_to_tile_5_27_1),
		.out_wire_0_2(horizontal_tile_5_26_to_tile_5_27_2),
		.out_wire_0_3(horizontal_tile_5_26_to_tile_5_27_3),
		.in_wire_0_0(horizontal_tile_5_27_to_tile_5_26_0),
		.in_wire_0_1(horizontal_tile_5_27_to_tile_5_26_1),
		.in_wire_0_2(horizontal_tile_5_27_to_tile_5_26_2),
		.in_wire_0_3(horizontal_tile_5_27_to_tile_5_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(187)
	);

	pe_tile pe_tile_5_27(
		.out_wire_3_0(vertical_tile_5_27_to_tile_4_27_0),
		.out_wire_3_1(vertical_tile_5_27_to_tile_4_27_1),
		.out_wire_3_2(vertical_tile_5_27_to_tile_4_27_2),
		.out_wire_3_3(vertical_tile_5_27_to_tile_4_27_3),
		.in_wire_3_0(vertical_tile_4_27_to_tile_5_27_0),
		.in_wire_3_1(vertical_tile_4_27_to_tile_5_27_1),
		.in_wire_3_2(vertical_tile_4_27_to_tile_5_27_2),
		.in_wire_3_3(vertical_tile_4_27_to_tile_5_27_3),
		.out_wire_1_0(vertical_tile_5_27_to_tile_6_27_0),
		.out_wire_1_1(vertical_tile_5_27_to_tile_6_27_1),
		.out_wire_1_2(vertical_tile_5_27_to_tile_6_27_2),
		.out_wire_1_3(vertical_tile_5_27_to_tile_6_27_3),
		.in_wire_1_0(vertical_tile_6_27_to_tile_5_27_0),
		.in_wire_1_1(vertical_tile_6_27_to_tile_5_27_1),
		.in_wire_1_2(vertical_tile_6_27_to_tile_5_27_2),
		.in_wire_1_3(vertical_tile_6_27_to_tile_5_27_3),
		.out_wire_2_0(horizontal_tile_5_27_to_tile_5_26_0),
		.out_wire_2_1(horizontal_tile_5_27_to_tile_5_26_1),
		.out_wire_2_2(horizontal_tile_5_27_to_tile_5_26_2),
		.out_wire_2_3(horizontal_tile_5_27_to_tile_5_26_3),
		.in_wire_2_0(horizontal_tile_5_26_to_tile_5_27_0),
		.in_wire_2_1(horizontal_tile_5_26_to_tile_5_27_1),
		.in_wire_2_2(horizontal_tile_5_26_to_tile_5_27_2),
		.in_wire_2_3(horizontal_tile_5_26_to_tile_5_27_3),
		.out_wire_0_0(horizontal_tile_5_27_to_tile_5_28_0),
		.out_wire_0_1(horizontal_tile_5_27_to_tile_5_28_1),
		.out_wire_0_2(horizontal_tile_5_27_to_tile_5_28_2),
		.out_wire_0_3(horizontal_tile_5_27_to_tile_5_28_3),
		.in_wire_0_0(horizontal_tile_5_28_to_tile_5_27_0),
		.in_wire_0_1(horizontal_tile_5_28_to_tile_5_27_1),
		.in_wire_0_2(horizontal_tile_5_28_to_tile_5_27_2),
		.in_wire_0_3(horizontal_tile_5_28_to_tile_5_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(188)
	);

	pe_tile pe_tile_5_28(
		.out_wire_3_0(vertical_tile_5_28_to_tile_4_28_0),
		.out_wire_3_1(vertical_tile_5_28_to_tile_4_28_1),
		.out_wire_3_2(vertical_tile_5_28_to_tile_4_28_2),
		.out_wire_3_3(vertical_tile_5_28_to_tile_4_28_3),
		.in_wire_3_0(vertical_tile_4_28_to_tile_5_28_0),
		.in_wire_3_1(vertical_tile_4_28_to_tile_5_28_1),
		.in_wire_3_2(vertical_tile_4_28_to_tile_5_28_2),
		.in_wire_3_3(vertical_tile_4_28_to_tile_5_28_3),
		.out_wire_1_0(vertical_tile_5_28_to_tile_6_28_0),
		.out_wire_1_1(vertical_tile_5_28_to_tile_6_28_1),
		.out_wire_1_2(vertical_tile_5_28_to_tile_6_28_2),
		.out_wire_1_3(vertical_tile_5_28_to_tile_6_28_3),
		.in_wire_1_0(vertical_tile_6_28_to_tile_5_28_0),
		.in_wire_1_1(vertical_tile_6_28_to_tile_5_28_1),
		.in_wire_1_2(vertical_tile_6_28_to_tile_5_28_2),
		.in_wire_1_3(vertical_tile_6_28_to_tile_5_28_3),
		.out_wire_2_0(horizontal_tile_5_28_to_tile_5_27_0),
		.out_wire_2_1(horizontal_tile_5_28_to_tile_5_27_1),
		.out_wire_2_2(horizontal_tile_5_28_to_tile_5_27_2),
		.out_wire_2_3(horizontal_tile_5_28_to_tile_5_27_3),
		.in_wire_2_0(horizontal_tile_5_27_to_tile_5_28_0),
		.in_wire_2_1(horizontal_tile_5_27_to_tile_5_28_1),
		.in_wire_2_2(horizontal_tile_5_27_to_tile_5_28_2),
		.in_wire_2_3(horizontal_tile_5_27_to_tile_5_28_3),
		.out_wire_0_0(horizontal_tile_5_28_to_tile_5_29_0),
		.out_wire_0_1(horizontal_tile_5_28_to_tile_5_29_1),
		.out_wire_0_2(horizontal_tile_5_28_to_tile_5_29_2),
		.out_wire_0_3(horizontal_tile_5_28_to_tile_5_29_3),
		.in_wire_0_0(horizontal_tile_5_29_to_tile_5_28_0),
		.in_wire_0_1(horizontal_tile_5_29_to_tile_5_28_1),
		.in_wire_0_2(horizontal_tile_5_29_to_tile_5_28_2),
		.in_wire_0_3(horizontal_tile_5_29_to_tile_5_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(189)
	);

	pe_tile pe_tile_5_29(
		.out_wire_3_0(vertical_tile_5_29_to_tile_4_29_0),
		.out_wire_3_1(vertical_tile_5_29_to_tile_4_29_1),
		.out_wire_3_2(vertical_tile_5_29_to_tile_4_29_2),
		.out_wire_3_3(vertical_tile_5_29_to_tile_4_29_3),
		.in_wire_3_0(vertical_tile_4_29_to_tile_5_29_0),
		.in_wire_3_1(vertical_tile_4_29_to_tile_5_29_1),
		.in_wire_3_2(vertical_tile_4_29_to_tile_5_29_2),
		.in_wire_3_3(vertical_tile_4_29_to_tile_5_29_3),
		.out_wire_1_0(vertical_tile_5_29_to_tile_6_29_0),
		.out_wire_1_1(vertical_tile_5_29_to_tile_6_29_1),
		.out_wire_1_2(vertical_tile_5_29_to_tile_6_29_2),
		.out_wire_1_3(vertical_tile_5_29_to_tile_6_29_3),
		.in_wire_1_0(vertical_tile_6_29_to_tile_5_29_0),
		.in_wire_1_1(vertical_tile_6_29_to_tile_5_29_1),
		.in_wire_1_2(vertical_tile_6_29_to_tile_5_29_2),
		.in_wire_1_3(vertical_tile_6_29_to_tile_5_29_3),
		.out_wire_2_0(horizontal_tile_5_29_to_tile_5_28_0),
		.out_wire_2_1(horizontal_tile_5_29_to_tile_5_28_1),
		.out_wire_2_2(horizontal_tile_5_29_to_tile_5_28_2),
		.out_wire_2_3(horizontal_tile_5_29_to_tile_5_28_3),
		.in_wire_2_0(horizontal_tile_5_28_to_tile_5_29_0),
		.in_wire_2_1(horizontal_tile_5_28_to_tile_5_29_1),
		.in_wire_2_2(horizontal_tile_5_28_to_tile_5_29_2),
		.in_wire_2_3(horizontal_tile_5_28_to_tile_5_29_3),
		.out_wire_0_0(horizontal_tile_5_29_to_tile_5_30_0),
		.out_wire_0_1(horizontal_tile_5_29_to_tile_5_30_1),
		.out_wire_0_2(horizontal_tile_5_29_to_tile_5_30_2),
		.out_wire_0_3(horizontal_tile_5_29_to_tile_5_30_3),
		.in_wire_0_0(horizontal_tile_5_30_to_tile_5_29_0),
		.in_wire_0_1(horizontal_tile_5_30_to_tile_5_29_1),
		.in_wire_0_2(horizontal_tile_5_30_to_tile_5_29_2),
		.in_wire_0_3(horizontal_tile_5_30_to_tile_5_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(190)
	);

	pe_tile pe_tile_5_30(
		.out_wire_3_0(vertical_tile_5_30_to_tile_4_30_0),
		.out_wire_3_1(vertical_tile_5_30_to_tile_4_30_1),
		.out_wire_3_2(vertical_tile_5_30_to_tile_4_30_2),
		.out_wire_3_3(vertical_tile_5_30_to_tile_4_30_3),
		.in_wire_3_0(vertical_tile_4_30_to_tile_5_30_0),
		.in_wire_3_1(vertical_tile_4_30_to_tile_5_30_1),
		.in_wire_3_2(vertical_tile_4_30_to_tile_5_30_2),
		.in_wire_3_3(vertical_tile_4_30_to_tile_5_30_3),
		.out_wire_1_0(vertical_tile_5_30_to_tile_6_30_0),
		.out_wire_1_1(vertical_tile_5_30_to_tile_6_30_1),
		.out_wire_1_2(vertical_tile_5_30_to_tile_6_30_2),
		.out_wire_1_3(vertical_tile_5_30_to_tile_6_30_3),
		.in_wire_1_0(vertical_tile_6_30_to_tile_5_30_0),
		.in_wire_1_1(vertical_tile_6_30_to_tile_5_30_1),
		.in_wire_1_2(vertical_tile_6_30_to_tile_5_30_2),
		.in_wire_1_3(vertical_tile_6_30_to_tile_5_30_3),
		.out_wire_2_0(horizontal_tile_5_30_to_tile_5_29_0),
		.out_wire_2_1(horizontal_tile_5_30_to_tile_5_29_1),
		.out_wire_2_2(horizontal_tile_5_30_to_tile_5_29_2),
		.out_wire_2_3(horizontal_tile_5_30_to_tile_5_29_3),
		.in_wire_2_0(horizontal_tile_5_29_to_tile_5_30_0),
		.in_wire_2_1(horizontal_tile_5_29_to_tile_5_30_1),
		.in_wire_2_2(horizontal_tile_5_29_to_tile_5_30_2),
		.in_wire_2_3(horizontal_tile_5_29_to_tile_5_30_3),
		.out_wire_0_0(horizontal_tile_5_30_to_tile_5_31_0),
		.out_wire_0_1(horizontal_tile_5_30_to_tile_5_31_1),
		.out_wire_0_2(horizontal_tile_5_30_to_tile_5_31_2),
		.out_wire_0_3(horizontal_tile_5_30_to_tile_5_31_3),
		.in_wire_0_0(horizontal_tile_5_31_to_tile_5_30_0),
		.in_wire_0_1(horizontal_tile_5_31_to_tile_5_30_1),
		.in_wire_0_2(horizontal_tile_5_31_to_tile_5_30_2),
		.in_wire_0_3(horizontal_tile_5_31_to_tile_5_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(191)
	);

	pe_tile_right pe_tile_5_31(
		.out_wire_3_0(vertical_tile_5_31_to_tile_4_31_0),
		.out_wire_3_1(vertical_tile_5_31_to_tile_4_31_1),
		.out_wire_3_2(vertical_tile_5_31_to_tile_4_31_2),
		.out_wire_3_3(vertical_tile_5_31_to_tile_4_31_3),
		.in_wire_3_0(vertical_tile_4_31_to_tile_5_31_0),
		.in_wire_3_1(vertical_tile_4_31_to_tile_5_31_1),
		.in_wire_3_2(vertical_tile_4_31_to_tile_5_31_2),
		.in_wire_3_3(vertical_tile_4_31_to_tile_5_31_3),
		.out_wire_1_0(vertical_tile_5_31_to_tile_6_31_0),
		.out_wire_1_1(vertical_tile_5_31_to_tile_6_31_1),
		.out_wire_1_2(vertical_tile_5_31_to_tile_6_31_2),
		.out_wire_1_3(vertical_tile_5_31_to_tile_6_31_3),
		.in_wire_1_0(vertical_tile_6_31_to_tile_5_31_0),
		.in_wire_1_1(vertical_tile_6_31_to_tile_5_31_1),
		.in_wire_1_2(vertical_tile_6_31_to_tile_5_31_2),
		.in_wire_1_3(vertical_tile_6_31_to_tile_5_31_3),
		.out_wire_2_0(horizontal_tile_5_31_to_tile_5_30_0),
		.out_wire_2_1(horizontal_tile_5_31_to_tile_5_30_1),
		.out_wire_2_2(horizontal_tile_5_31_to_tile_5_30_2),
		.out_wire_2_3(horizontal_tile_5_31_to_tile_5_30_3),
		.in_wire_2_0(horizontal_tile_5_30_to_tile_5_31_0),
		.in_wire_2_1(horizontal_tile_5_30_to_tile_5_31_1),
		.in_wire_2_2(horizontal_tile_5_30_to_tile_5_31_2),
		.in_wire_2_3(horizontal_tile_5_30_to_tile_5_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(192)
	);

	pe_tile_left pe_tile_6_0(
		.out_wire_3_0(vertical_tile_6_0_to_tile_5_0_0),
		.out_wire_3_1(vertical_tile_6_0_to_tile_5_0_1),
		.out_wire_3_2(vertical_tile_6_0_to_tile_5_0_2),
		.out_wire_3_3(vertical_tile_6_0_to_tile_5_0_3),
		.in_wire_3_0(vertical_tile_5_0_to_tile_6_0_0),
		.in_wire_3_1(vertical_tile_5_0_to_tile_6_0_1),
		.in_wire_3_2(vertical_tile_5_0_to_tile_6_0_2),
		.in_wire_3_3(vertical_tile_5_0_to_tile_6_0_3),
		.out_wire_1_0(vertical_tile_6_0_to_tile_7_0_0),
		.out_wire_1_1(vertical_tile_6_0_to_tile_7_0_1),
		.out_wire_1_2(vertical_tile_6_0_to_tile_7_0_2),
		.out_wire_1_3(vertical_tile_6_0_to_tile_7_0_3),
		.in_wire_1_0(vertical_tile_7_0_to_tile_6_0_0),
		.in_wire_1_1(vertical_tile_7_0_to_tile_6_0_1),
		.in_wire_1_2(vertical_tile_7_0_to_tile_6_0_2),
		.in_wire_1_3(vertical_tile_7_0_to_tile_6_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_6_0_to_tile_6_1_0),
		.out_wire_0_1(horizontal_tile_6_0_to_tile_6_1_1),
		.out_wire_0_2(horizontal_tile_6_0_to_tile_6_1_2),
		.out_wire_0_3(horizontal_tile_6_0_to_tile_6_1_3),
		.in_wire_0_0(horizontal_tile_6_1_to_tile_6_0_0),
		.in_wire_0_1(horizontal_tile_6_1_to_tile_6_0_1),
		.in_wire_0_2(horizontal_tile_6_1_to_tile_6_0_2),
		.in_wire_0_3(horizontal_tile_6_1_to_tile_6_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(193)
	);

	pe_tile pe_tile_6_1(
		.out_wire_3_0(vertical_tile_6_1_to_tile_5_1_0),
		.out_wire_3_1(vertical_tile_6_1_to_tile_5_1_1),
		.out_wire_3_2(vertical_tile_6_1_to_tile_5_1_2),
		.out_wire_3_3(vertical_tile_6_1_to_tile_5_1_3),
		.in_wire_3_0(vertical_tile_5_1_to_tile_6_1_0),
		.in_wire_3_1(vertical_tile_5_1_to_tile_6_1_1),
		.in_wire_3_2(vertical_tile_5_1_to_tile_6_1_2),
		.in_wire_3_3(vertical_tile_5_1_to_tile_6_1_3),
		.out_wire_1_0(vertical_tile_6_1_to_tile_7_1_0),
		.out_wire_1_1(vertical_tile_6_1_to_tile_7_1_1),
		.out_wire_1_2(vertical_tile_6_1_to_tile_7_1_2),
		.out_wire_1_3(vertical_tile_6_1_to_tile_7_1_3),
		.in_wire_1_0(vertical_tile_7_1_to_tile_6_1_0),
		.in_wire_1_1(vertical_tile_7_1_to_tile_6_1_1),
		.in_wire_1_2(vertical_tile_7_1_to_tile_6_1_2),
		.in_wire_1_3(vertical_tile_7_1_to_tile_6_1_3),
		.out_wire_2_0(horizontal_tile_6_1_to_tile_6_0_0),
		.out_wire_2_1(horizontal_tile_6_1_to_tile_6_0_1),
		.out_wire_2_2(horizontal_tile_6_1_to_tile_6_0_2),
		.out_wire_2_3(horizontal_tile_6_1_to_tile_6_0_3),
		.in_wire_2_0(horizontal_tile_6_0_to_tile_6_1_0),
		.in_wire_2_1(horizontal_tile_6_0_to_tile_6_1_1),
		.in_wire_2_2(horizontal_tile_6_0_to_tile_6_1_2),
		.in_wire_2_3(horizontal_tile_6_0_to_tile_6_1_3),
		.out_wire_0_0(horizontal_tile_6_1_to_tile_6_2_0),
		.out_wire_0_1(horizontal_tile_6_1_to_tile_6_2_1),
		.out_wire_0_2(horizontal_tile_6_1_to_tile_6_2_2),
		.out_wire_0_3(horizontal_tile_6_1_to_tile_6_2_3),
		.in_wire_0_0(horizontal_tile_6_2_to_tile_6_1_0),
		.in_wire_0_1(horizontal_tile_6_2_to_tile_6_1_1),
		.in_wire_0_2(horizontal_tile_6_2_to_tile_6_1_2),
		.in_wire_0_3(horizontal_tile_6_2_to_tile_6_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(194)
	);

	pe_tile pe_tile_6_2(
		.out_wire_3_0(vertical_tile_6_2_to_tile_5_2_0),
		.out_wire_3_1(vertical_tile_6_2_to_tile_5_2_1),
		.out_wire_3_2(vertical_tile_6_2_to_tile_5_2_2),
		.out_wire_3_3(vertical_tile_6_2_to_tile_5_2_3),
		.in_wire_3_0(vertical_tile_5_2_to_tile_6_2_0),
		.in_wire_3_1(vertical_tile_5_2_to_tile_6_2_1),
		.in_wire_3_2(vertical_tile_5_2_to_tile_6_2_2),
		.in_wire_3_3(vertical_tile_5_2_to_tile_6_2_3),
		.out_wire_1_0(vertical_tile_6_2_to_tile_7_2_0),
		.out_wire_1_1(vertical_tile_6_2_to_tile_7_2_1),
		.out_wire_1_2(vertical_tile_6_2_to_tile_7_2_2),
		.out_wire_1_3(vertical_tile_6_2_to_tile_7_2_3),
		.in_wire_1_0(vertical_tile_7_2_to_tile_6_2_0),
		.in_wire_1_1(vertical_tile_7_2_to_tile_6_2_1),
		.in_wire_1_2(vertical_tile_7_2_to_tile_6_2_2),
		.in_wire_1_3(vertical_tile_7_2_to_tile_6_2_3),
		.out_wire_2_0(horizontal_tile_6_2_to_tile_6_1_0),
		.out_wire_2_1(horizontal_tile_6_2_to_tile_6_1_1),
		.out_wire_2_2(horizontal_tile_6_2_to_tile_6_1_2),
		.out_wire_2_3(horizontal_tile_6_2_to_tile_6_1_3),
		.in_wire_2_0(horizontal_tile_6_1_to_tile_6_2_0),
		.in_wire_2_1(horizontal_tile_6_1_to_tile_6_2_1),
		.in_wire_2_2(horizontal_tile_6_1_to_tile_6_2_2),
		.in_wire_2_3(horizontal_tile_6_1_to_tile_6_2_3),
		.out_wire_0_0(horizontal_tile_6_2_to_tile_6_3_0),
		.out_wire_0_1(horizontal_tile_6_2_to_tile_6_3_1),
		.out_wire_0_2(horizontal_tile_6_2_to_tile_6_3_2),
		.out_wire_0_3(horizontal_tile_6_2_to_tile_6_3_3),
		.in_wire_0_0(horizontal_tile_6_3_to_tile_6_2_0),
		.in_wire_0_1(horizontal_tile_6_3_to_tile_6_2_1),
		.in_wire_0_2(horizontal_tile_6_3_to_tile_6_2_2),
		.in_wire_0_3(horizontal_tile_6_3_to_tile_6_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(195)
	);

	pe_tile pe_tile_6_3(
		.out_wire_3_0(vertical_tile_6_3_to_tile_5_3_0),
		.out_wire_3_1(vertical_tile_6_3_to_tile_5_3_1),
		.out_wire_3_2(vertical_tile_6_3_to_tile_5_3_2),
		.out_wire_3_3(vertical_tile_6_3_to_tile_5_3_3),
		.in_wire_3_0(vertical_tile_5_3_to_tile_6_3_0),
		.in_wire_3_1(vertical_tile_5_3_to_tile_6_3_1),
		.in_wire_3_2(vertical_tile_5_3_to_tile_6_3_2),
		.in_wire_3_3(vertical_tile_5_3_to_tile_6_3_3),
		.out_wire_1_0(vertical_tile_6_3_to_tile_7_3_0),
		.out_wire_1_1(vertical_tile_6_3_to_tile_7_3_1),
		.out_wire_1_2(vertical_tile_6_3_to_tile_7_3_2),
		.out_wire_1_3(vertical_tile_6_3_to_tile_7_3_3),
		.in_wire_1_0(vertical_tile_7_3_to_tile_6_3_0),
		.in_wire_1_1(vertical_tile_7_3_to_tile_6_3_1),
		.in_wire_1_2(vertical_tile_7_3_to_tile_6_3_2),
		.in_wire_1_3(vertical_tile_7_3_to_tile_6_3_3),
		.out_wire_2_0(horizontal_tile_6_3_to_tile_6_2_0),
		.out_wire_2_1(horizontal_tile_6_3_to_tile_6_2_1),
		.out_wire_2_2(horizontal_tile_6_3_to_tile_6_2_2),
		.out_wire_2_3(horizontal_tile_6_3_to_tile_6_2_3),
		.in_wire_2_0(horizontal_tile_6_2_to_tile_6_3_0),
		.in_wire_2_1(horizontal_tile_6_2_to_tile_6_3_1),
		.in_wire_2_2(horizontal_tile_6_2_to_tile_6_3_2),
		.in_wire_2_3(horizontal_tile_6_2_to_tile_6_3_3),
		.out_wire_0_0(horizontal_tile_6_3_to_tile_6_4_0),
		.out_wire_0_1(horizontal_tile_6_3_to_tile_6_4_1),
		.out_wire_0_2(horizontal_tile_6_3_to_tile_6_4_2),
		.out_wire_0_3(horizontal_tile_6_3_to_tile_6_4_3),
		.in_wire_0_0(horizontal_tile_6_4_to_tile_6_3_0),
		.in_wire_0_1(horizontal_tile_6_4_to_tile_6_3_1),
		.in_wire_0_2(horizontal_tile_6_4_to_tile_6_3_2),
		.in_wire_0_3(horizontal_tile_6_4_to_tile_6_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(196)
	);

	pe_tile pe_tile_6_4(
		.out_wire_3_0(vertical_tile_6_4_to_tile_5_4_0),
		.out_wire_3_1(vertical_tile_6_4_to_tile_5_4_1),
		.out_wire_3_2(vertical_tile_6_4_to_tile_5_4_2),
		.out_wire_3_3(vertical_tile_6_4_to_tile_5_4_3),
		.in_wire_3_0(vertical_tile_5_4_to_tile_6_4_0),
		.in_wire_3_1(vertical_tile_5_4_to_tile_6_4_1),
		.in_wire_3_2(vertical_tile_5_4_to_tile_6_4_2),
		.in_wire_3_3(vertical_tile_5_4_to_tile_6_4_3),
		.out_wire_1_0(vertical_tile_6_4_to_tile_7_4_0),
		.out_wire_1_1(vertical_tile_6_4_to_tile_7_4_1),
		.out_wire_1_2(vertical_tile_6_4_to_tile_7_4_2),
		.out_wire_1_3(vertical_tile_6_4_to_tile_7_4_3),
		.in_wire_1_0(vertical_tile_7_4_to_tile_6_4_0),
		.in_wire_1_1(vertical_tile_7_4_to_tile_6_4_1),
		.in_wire_1_2(vertical_tile_7_4_to_tile_6_4_2),
		.in_wire_1_3(vertical_tile_7_4_to_tile_6_4_3),
		.out_wire_2_0(horizontal_tile_6_4_to_tile_6_3_0),
		.out_wire_2_1(horizontal_tile_6_4_to_tile_6_3_1),
		.out_wire_2_2(horizontal_tile_6_4_to_tile_6_3_2),
		.out_wire_2_3(horizontal_tile_6_4_to_tile_6_3_3),
		.in_wire_2_0(horizontal_tile_6_3_to_tile_6_4_0),
		.in_wire_2_1(horizontal_tile_6_3_to_tile_6_4_1),
		.in_wire_2_2(horizontal_tile_6_3_to_tile_6_4_2),
		.in_wire_2_3(horizontal_tile_6_3_to_tile_6_4_3),
		.out_wire_0_0(horizontal_tile_6_4_to_tile_6_5_0),
		.out_wire_0_1(horizontal_tile_6_4_to_tile_6_5_1),
		.out_wire_0_2(horizontal_tile_6_4_to_tile_6_5_2),
		.out_wire_0_3(horizontal_tile_6_4_to_tile_6_5_3),
		.in_wire_0_0(horizontal_tile_6_5_to_tile_6_4_0),
		.in_wire_0_1(horizontal_tile_6_5_to_tile_6_4_1),
		.in_wire_0_2(horizontal_tile_6_5_to_tile_6_4_2),
		.in_wire_0_3(horizontal_tile_6_5_to_tile_6_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(197)
	);

	pe_tile pe_tile_6_5(
		.out_wire_3_0(vertical_tile_6_5_to_tile_5_5_0),
		.out_wire_3_1(vertical_tile_6_5_to_tile_5_5_1),
		.out_wire_3_2(vertical_tile_6_5_to_tile_5_5_2),
		.out_wire_3_3(vertical_tile_6_5_to_tile_5_5_3),
		.in_wire_3_0(vertical_tile_5_5_to_tile_6_5_0),
		.in_wire_3_1(vertical_tile_5_5_to_tile_6_5_1),
		.in_wire_3_2(vertical_tile_5_5_to_tile_6_5_2),
		.in_wire_3_3(vertical_tile_5_5_to_tile_6_5_3),
		.out_wire_1_0(vertical_tile_6_5_to_tile_7_5_0),
		.out_wire_1_1(vertical_tile_6_5_to_tile_7_5_1),
		.out_wire_1_2(vertical_tile_6_5_to_tile_7_5_2),
		.out_wire_1_3(vertical_tile_6_5_to_tile_7_5_3),
		.in_wire_1_0(vertical_tile_7_5_to_tile_6_5_0),
		.in_wire_1_1(vertical_tile_7_5_to_tile_6_5_1),
		.in_wire_1_2(vertical_tile_7_5_to_tile_6_5_2),
		.in_wire_1_3(vertical_tile_7_5_to_tile_6_5_3),
		.out_wire_2_0(horizontal_tile_6_5_to_tile_6_4_0),
		.out_wire_2_1(horizontal_tile_6_5_to_tile_6_4_1),
		.out_wire_2_2(horizontal_tile_6_5_to_tile_6_4_2),
		.out_wire_2_3(horizontal_tile_6_5_to_tile_6_4_3),
		.in_wire_2_0(horizontal_tile_6_4_to_tile_6_5_0),
		.in_wire_2_1(horizontal_tile_6_4_to_tile_6_5_1),
		.in_wire_2_2(horizontal_tile_6_4_to_tile_6_5_2),
		.in_wire_2_3(horizontal_tile_6_4_to_tile_6_5_3),
		.out_wire_0_0(horizontal_tile_6_5_to_tile_6_6_0),
		.out_wire_0_1(horizontal_tile_6_5_to_tile_6_6_1),
		.out_wire_0_2(horizontal_tile_6_5_to_tile_6_6_2),
		.out_wire_0_3(horizontal_tile_6_5_to_tile_6_6_3),
		.in_wire_0_0(horizontal_tile_6_6_to_tile_6_5_0),
		.in_wire_0_1(horizontal_tile_6_6_to_tile_6_5_1),
		.in_wire_0_2(horizontal_tile_6_6_to_tile_6_5_2),
		.in_wire_0_3(horizontal_tile_6_6_to_tile_6_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(198)
	);

	pe_tile pe_tile_6_6(
		.out_wire_3_0(vertical_tile_6_6_to_tile_5_6_0),
		.out_wire_3_1(vertical_tile_6_6_to_tile_5_6_1),
		.out_wire_3_2(vertical_tile_6_6_to_tile_5_6_2),
		.out_wire_3_3(vertical_tile_6_6_to_tile_5_6_3),
		.in_wire_3_0(vertical_tile_5_6_to_tile_6_6_0),
		.in_wire_3_1(vertical_tile_5_6_to_tile_6_6_1),
		.in_wire_3_2(vertical_tile_5_6_to_tile_6_6_2),
		.in_wire_3_3(vertical_tile_5_6_to_tile_6_6_3),
		.out_wire_1_0(vertical_tile_6_6_to_tile_7_6_0),
		.out_wire_1_1(vertical_tile_6_6_to_tile_7_6_1),
		.out_wire_1_2(vertical_tile_6_6_to_tile_7_6_2),
		.out_wire_1_3(vertical_tile_6_6_to_tile_7_6_3),
		.in_wire_1_0(vertical_tile_7_6_to_tile_6_6_0),
		.in_wire_1_1(vertical_tile_7_6_to_tile_6_6_1),
		.in_wire_1_2(vertical_tile_7_6_to_tile_6_6_2),
		.in_wire_1_3(vertical_tile_7_6_to_tile_6_6_3),
		.out_wire_2_0(horizontal_tile_6_6_to_tile_6_5_0),
		.out_wire_2_1(horizontal_tile_6_6_to_tile_6_5_1),
		.out_wire_2_2(horizontal_tile_6_6_to_tile_6_5_2),
		.out_wire_2_3(horizontal_tile_6_6_to_tile_6_5_3),
		.in_wire_2_0(horizontal_tile_6_5_to_tile_6_6_0),
		.in_wire_2_1(horizontal_tile_6_5_to_tile_6_6_1),
		.in_wire_2_2(horizontal_tile_6_5_to_tile_6_6_2),
		.in_wire_2_3(horizontal_tile_6_5_to_tile_6_6_3),
		.out_wire_0_0(horizontal_tile_6_6_to_tile_6_7_0),
		.out_wire_0_1(horizontal_tile_6_6_to_tile_6_7_1),
		.out_wire_0_2(horizontal_tile_6_6_to_tile_6_7_2),
		.out_wire_0_3(horizontal_tile_6_6_to_tile_6_7_3),
		.in_wire_0_0(horizontal_tile_6_7_to_tile_6_6_0),
		.in_wire_0_1(horizontal_tile_6_7_to_tile_6_6_1),
		.in_wire_0_2(horizontal_tile_6_7_to_tile_6_6_2),
		.in_wire_0_3(horizontal_tile_6_7_to_tile_6_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(199)
	);

	pe_tile pe_tile_6_7(
		.out_wire_3_0(vertical_tile_6_7_to_tile_5_7_0),
		.out_wire_3_1(vertical_tile_6_7_to_tile_5_7_1),
		.out_wire_3_2(vertical_tile_6_7_to_tile_5_7_2),
		.out_wire_3_3(vertical_tile_6_7_to_tile_5_7_3),
		.in_wire_3_0(vertical_tile_5_7_to_tile_6_7_0),
		.in_wire_3_1(vertical_tile_5_7_to_tile_6_7_1),
		.in_wire_3_2(vertical_tile_5_7_to_tile_6_7_2),
		.in_wire_3_3(vertical_tile_5_7_to_tile_6_7_3),
		.out_wire_1_0(vertical_tile_6_7_to_tile_7_7_0),
		.out_wire_1_1(vertical_tile_6_7_to_tile_7_7_1),
		.out_wire_1_2(vertical_tile_6_7_to_tile_7_7_2),
		.out_wire_1_3(vertical_tile_6_7_to_tile_7_7_3),
		.in_wire_1_0(vertical_tile_7_7_to_tile_6_7_0),
		.in_wire_1_1(vertical_tile_7_7_to_tile_6_7_1),
		.in_wire_1_2(vertical_tile_7_7_to_tile_6_7_2),
		.in_wire_1_3(vertical_tile_7_7_to_tile_6_7_3),
		.out_wire_2_0(horizontal_tile_6_7_to_tile_6_6_0),
		.out_wire_2_1(horizontal_tile_6_7_to_tile_6_6_1),
		.out_wire_2_2(horizontal_tile_6_7_to_tile_6_6_2),
		.out_wire_2_3(horizontal_tile_6_7_to_tile_6_6_3),
		.in_wire_2_0(horizontal_tile_6_6_to_tile_6_7_0),
		.in_wire_2_1(horizontal_tile_6_6_to_tile_6_7_1),
		.in_wire_2_2(horizontal_tile_6_6_to_tile_6_7_2),
		.in_wire_2_3(horizontal_tile_6_6_to_tile_6_7_3),
		.out_wire_0_0(horizontal_tile_6_7_to_tile_6_8_0),
		.out_wire_0_1(horizontal_tile_6_7_to_tile_6_8_1),
		.out_wire_0_2(horizontal_tile_6_7_to_tile_6_8_2),
		.out_wire_0_3(horizontal_tile_6_7_to_tile_6_8_3),
		.in_wire_0_0(horizontal_tile_6_8_to_tile_6_7_0),
		.in_wire_0_1(horizontal_tile_6_8_to_tile_6_7_1),
		.in_wire_0_2(horizontal_tile_6_8_to_tile_6_7_2),
		.in_wire_0_3(horizontal_tile_6_8_to_tile_6_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(200)
	);

	pe_tile pe_tile_6_8(
		.out_wire_3_0(vertical_tile_6_8_to_tile_5_8_0),
		.out_wire_3_1(vertical_tile_6_8_to_tile_5_8_1),
		.out_wire_3_2(vertical_tile_6_8_to_tile_5_8_2),
		.out_wire_3_3(vertical_tile_6_8_to_tile_5_8_3),
		.in_wire_3_0(vertical_tile_5_8_to_tile_6_8_0),
		.in_wire_3_1(vertical_tile_5_8_to_tile_6_8_1),
		.in_wire_3_2(vertical_tile_5_8_to_tile_6_8_2),
		.in_wire_3_3(vertical_tile_5_8_to_tile_6_8_3),
		.out_wire_1_0(vertical_tile_6_8_to_tile_7_8_0),
		.out_wire_1_1(vertical_tile_6_8_to_tile_7_8_1),
		.out_wire_1_2(vertical_tile_6_8_to_tile_7_8_2),
		.out_wire_1_3(vertical_tile_6_8_to_tile_7_8_3),
		.in_wire_1_0(vertical_tile_7_8_to_tile_6_8_0),
		.in_wire_1_1(vertical_tile_7_8_to_tile_6_8_1),
		.in_wire_1_2(vertical_tile_7_8_to_tile_6_8_2),
		.in_wire_1_3(vertical_tile_7_8_to_tile_6_8_3),
		.out_wire_2_0(horizontal_tile_6_8_to_tile_6_7_0),
		.out_wire_2_1(horizontal_tile_6_8_to_tile_6_7_1),
		.out_wire_2_2(horizontal_tile_6_8_to_tile_6_7_2),
		.out_wire_2_3(horizontal_tile_6_8_to_tile_6_7_3),
		.in_wire_2_0(horizontal_tile_6_7_to_tile_6_8_0),
		.in_wire_2_1(horizontal_tile_6_7_to_tile_6_8_1),
		.in_wire_2_2(horizontal_tile_6_7_to_tile_6_8_2),
		.in_wire_2_3(horizontal_tile_6_7_to_tile_6_8_3),
		.out_wire_0_0(horizontal_tile_6_8_to_tile_6_9_0),
		.out_wire_0_1(horizontal_tile_6_8_to_tile_6_9_1),
		.out_wire_0_2(horizontal_tile_6_8_to_tile_6_9_2),
		.out_wire_0_3(horizontal_tile_6_8_to_tile_6_9_3),
		.in_wire_0_0(horizontal_tile_6_9_to_tile_6_8_0),
		.in_wire_0_1(horizontal_tile_6_9_to_tile_6_8_1),
		.in_wire_0_2(horizontal_tile_6_9_to_tile_6_8_2),
		.in_wire_0_3(horizontal_tile_6_9_to_tile_6_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(201)
	);

	pe_tile pe_tile_6_9(
		.out_wire_3_0(vertical_tile_6_9_to_tile_5_9_0),
		.out_wire_3_1(vertical_tile_6_9_to_tile_5_9_1),
		.out_wire_3_2(vertical_tile_6_9_to_tile_5_9_2),
		.out_wire_3_3(vertical_tile_6_9_to_tile_5_9_3),
		.in_wire_3_0(vertical_tile_5_9_to_tile_6_9_0),
		.in_wire_3_1(vertical_tile_5_9_to_tile_6_9_1),
		.in_wire_3_2(vertical_tile_5_9_to_tile_6_9_2),
		.in_wire_3_3(vertical_tile_5_9_to_tile_6_9_3),
		.out_wire_1_0(vertical_tile_6_9_to_tile_7_9_0),
		.out_wire_1_1(vertical_tile_6_9_to_tile_7_9_1),
		.out_wire_1_2(vertical_tile_6_9_to_tile_7_9_2),
		.out_wire_1_3(vertical_tile_6_9_to_tile_7_9_3),
		.in_wire_1_0(vertical_tile_7_9_to_tile_6_9_0),
		.in_wire_1_1(vertical_tile_7_9_to_tile_6_9_1),
		.in_wire_1_2(vertical_tile_7_9_to_tile_6_9_2),
		.in_wire_1_3(vertical_tile_7_9_to_tile_6_9_3),
		.out_wire_2_0(horizontal_tile_6_9_to_tile_6_8_0),
		.out_wire_2_1(horizontal_tile_6_9_to_tile_6_8_1),
		.out_wire_2_2(horizontal_tile_6_9_to_tile_6_8_2),
		.out_wire_2_3(horizontal_tile_6_9_to_tile_6_8_3),
		.in_wire_2_0(horizontal_tile_6_8_to_tile_6_9_0),
		.in_wire_2_1(horizontal_tile_6_8_to_tile_6_9_1),
		.in_wire_2_2(horizontal_tile_6_8_to_tile_6_9_2),
		.in_wire_2_3(horizontal_tile_6_8_to_tile_6_9_3),
		.out_wire_0_0(horizontal_tile_6_9_to_tile_6_10_0),
		.out_wire_0_1(horizontal_tile_6_9_to_tile_6_10_1),
		.out_wire_0_2(horizontal_tile_6_9_to_tile_6_10_2),
		.out_wire_0_3(horizontal_tile_6_9_to_tile_6_10_3),
		.in_wire_0_0(horizontal_tile_6_10_to_tile_6_9_0),
		.in_wire_0_1(horizontal_tile_6_10_to_tile_6_9_1),
		.in_wire_0_2(horizontal_tile_6_10_to_tile_6_9_2),
		.in_wire_0_3(horizontal_tile_6_10_to_tile_6_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(202)
	);

	pe_tile pe_tile_6_10(
		.out_wire_3_0(vertical_tile_6_10_to_tile_5_10_0),
		.out_wire_3_1(vertical_tile_6_10_to_tile_5_10_1),
		.out_wire_3_2(vertical_tile_6_10_to_tile_5_10_2),
		.out_wire_3_3(vertical_tile_6_10_to_tile_5_10_3),
		.in_wire_3_0(vertical_tile_5_10_to_tile_6_10_0),
		.in_wire_3_1(vertical_tile_5_10_to_tile_6_10_1),
		.in_wire_3_2(vertical_tile_5_10_to_tile_6_10_2),
		.in_wire_3_3(vertical_tile_5_10_to_tile_6_10_3),
		.out_wire_1_0(vertical_tile_6_10_to_tile_7_10_0),
		.out_wire_1_1(vertical_tile_6_10_to_tile_7_10_1),
		.out_wire_1_2(vertical_tile_6_10_to_tile_7_10_2),
		.out_wire_1_3(vertical_tile_6_10_to_tile_7_10_3),
		.in_wire_1_0(vertical_tile_7_10_to_tile_6_10_0),
		.in_wire_1_1(vertical_tile_7_10_to_tile_6_10_1),
		.in_wire_1_2(vertical_tile_7_10_to_tile_6_10_2),
		.in_wire_1_3(vertical_tile_7_10_to_tile_6_10_3),
		.out_wire_2_0(horizontal_tile_6_10_to_tile_6_9_0),
		.out_wire_2_1(horizontal_tile_6_10_to_tile_6_9_1),
		.out_wire_2_2(horizontal_tile_6_10_to_tile_6_9_2),
		.out_wire_2_3(horizontal_tile_6_10_to_tile_6_9_3),
		.in_wire_2_0(horizontal_tile_6_9_to_tile_6_10_0),
		.in_wire_2_1(horizontal_tile_6_9_to_tile_6_10_1),
		.in_wire_2_2(horizontal_tile_6_9_to_tile_6_10_2),
		.in_wire_2_3(horizontal_tile_6_9_to_tile_6_10_3),
		.out_wire_0_0(horizontal_tile_6_10_to_tile_6_11_0),
		.out_wire_0_1(horizontal_tile_6_10_to_tile_6_11_1),
		.out_wire_0_2(horizontal_tile_6_10_to_tile_6_11_2),
		.out_wire_0_3(horizontal_tile_6_10_to_tile_6_11_3),
		.in_wire_0_0(horizontal_tile_6_11_to_tile_6_10_0),
		.in_wire_0_1(horizontal_tile_6_11_to_tile_6_10_1),
		.in_wire_0_2(horizontal_tile_6_11_to_tile_6_10_2),
		.in_wire_0_3(horizontal_tile_6_11_to_tile_6_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(203)
	);

	pe_tile pe_tile_6_11(
		.out_wire_3_0(vertical_tile_6_11_to_tile_5_11_0),
		.out_wire_3_1(vertical_tile_6_11_to_tile_5_11_1),
		.out_wire_3_2(vertical_tile_6_11_to_tile_5_11_2),
		.out_wire_3_3(vertical_tile_6_11_to_tile_5_11_3),
		.in_wire_3_0(vertical_tile_5_11_to_tile_6_11_0),
		.in_wire_3_1(vertical_tile_5_11_to_tile_6_11_1),
		.in_wire_3_2(vertical_tile_5_11_to_tile_6_11_2),
		.in_wire_3_3(vertical_tile_5_11_to_tile_6_11_3),
		.out_wire_1_0(vertical_tile_6_11_to_tile_7_11_0),
		.out_wire_1_1(vertical_tile_6_11_to_tile_7_11_1),
		.out_wire_1_2(vertical_tile_6_11_to_tile_7_11_2),
		.out_wire_1_3(vertical_tile_6_11_to_tile_7_11_3),
		.in_wire_1_0(vertical_tile_7_11_to_tile_6_11_0),
		.in_wire_1_1(vertical_tile_7_11_to_tile_6_11_1),
		.in_wire_1_2(vertical_tile_7_11_to_tile_6_11_2),
		.in_wire_1_3(vertical_tile_7_11_to_tile_6_11_3),
		.out_wire_2_0(horizontal_tile_6_11_to_tile_6_10_0),
		.out_wire_2_1(horizontal_tile_6_11_to_tile_6_10_1),
		.out_wire_2_2(horizontal_tile_6_11_to_tile_6_10_2),
		.out_wire_2_3(horizontal_tile_6_11_to_tile_6_10_3),
		.in_wire_2_0(horizontal_tile_6_10_to_tile_6_11_0),
		.in_wire_2_1(horizontal_tile_6_10_to_tile_6_11_1),
		.in_wire_2_2(horizontal_tile_6_10_to_tile_6_11_2),
		.in_wire_2_3(horizontal_tile_6_10_to_tile_6_11_3),
		.out_wire_0_0(horizontal_tile_6_11_to_tile_6_12_0),
		.out_wire_0_1(horizontal_tile_6_11_to_tile_6_12_1),
		.out_wire_0_2(horizontal_tile_6_11_to_tile_6_12_2),
		.out_wire_0_3(horizontal_tile_6_11_to_tile_6_12_3),
		.in_wire_0_0(horizontal_tile_6_12_to_tile_6_11_0),
		.in_wire_0_1(horizontal_tile_6_12_to_tile_6_11_1),
		.in_wire_0_2(horizontal_tile_6_12_to_tile_6_11_2),
		.in_wire_0_3(horizontal_tile_6_12_to_tile_6_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(204)
	);

	pe_tile pe_tile_6_12(
		.out_wire_3_0(vertical_tile_6_12_to_tile_5_12_0),
		.out_wire_3_1(vertical_tile_6_12_to_tile_5_12_1),
		.out_wire_3_2(vertical_tile_6_12_to_tile_5_12_2),
		.out_wire_3_3(vertical_tile_6_12_to_tile_5_12_3),
		.in_wire_3_0(vertical_tile_5_12_to_tile_6_12_0),
		.in_wire_3_1(vertical_tile_5_12_to_tile_6_12_1),
		.in_wire_3_2(vertical_tile_5_12_to_tile_6_12_2),
		.in_wire_3_3(vertical_tile_5_12_to_tile_6_12_3),
		.out_wire_1_0(vertical_tile_6_12_to_tile_7_12_0),
		.out_wire_1_1(vertical_tile_6_12_to_tile_7_12_1),
		.out_wire_1_2(vertical_tile_6_12_to_tile_7_12_2),
		.out_wire_1_3(vertical_tile_6_12_to_tile_7_12_3),
		.in_wire_1_0(vertical_tile_7_12_to_tile_6_12_0),
		.in_wire_1_1(vertical_tile_7_12_to_tile_6_12_1),
		.in_wire_1_2(vertical_tile_7_12_to_tile_6_12_2),
		.in_wire_1_3(vertical_tile_7_12_to_tile_6_12_3),
		.out_wire_2_0(horizontal_tile_6_12_to_tile_6_11_0),
		.out_wire_2_1(horizontal_tile_6_12_to_tile_6_11_1),
		.out_wire_2_2(horizontal_tile_6_12_to_tile_6_11_2),
		.out_wire_2_3(horizontal_tile_6_12_to_tile_6_11_3),
		.in_wire_2_0(horizontal_tile_6_11_to_tile_6_12_0),
		.in_wire_2_1(horizontal_tile_6_11_to_tile_6_12_1),
		.in_wire_2_2(horizontal_tile_6_11_to_tile_6_12_2),
		.in_wire_2_3(horizontal_tile_6_11_to_tile_6_12_3),
		.out_wire_0_0(horizontal_tile_6_12_to_tile_6_13_0),
		.out_wire_0_1(horizontal_tile_6_12_to_tile_6_13_1),
		.out_wire_0_2(horizontal_tile_6_12_to_tile_6_13_2),
		.out_wire_0_3(horizontal_tile_6_12_to_tile_6_13_3),
		.in_wire_0_0(horizontal_tile_6_13_to_tile_6_12_0),
		.in_wire_0_1(horizontal_tile_6_13_to_tile_6_12_1),
		.in_wire_0_2(horizontal_tile_6_13_to_tile_6_12_2),
		.in_wire_0_3(horizontal_tile_6_13_to_tile_6_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(205)
	);

	pe_tile pe_tile_6_13(
		.out_wire_3_0(vertical_tile_6_13_to_tile_5_13_0),
		.out_wire_3_1(vertical_tile_6_13_to_tile_5_13_1),
		.out_wire_3_2(vertical_tile_6_13_to_tile_5_13_2),
		.out_wire_3_3(vertical_tile_6_13_to_tile_5_13_3),
		.in_wire_3_0(vertical_tile_5_13_to_tile_6_13_0),
		.in_wire_3_1(vertical_tile_5_13_to_tile_6_13_1),
		.in_wire_3_2(vertical_tile_5_13_to_tile_6_13_2),
		.in_wire_3_3(vertical_tile_5_13_to_tile_6_13_3),
		.out_wire_1_0(vertical_tile_6_13_to_tile_7_13_0),
		.out_wire_1_1(vertical_tile_6_13_to_tile_7_13_1),
		.out_wire_1_2(vertical_tile_6_13_to_tile_7_13_2),
		.out_wire_1_3(vertical_tile_6_13_to_tile_7_13_3),
		.in_wire_1_0(vertical_tile_7_13_to_tile_6_13_0),
		.in_wire_1_1(vertical_tile_7_13_to_tile_6_13_1),
		.in_wire_1_2(vertical_tile_7_13_to_tile_6_13_2),
		.in_wire_1_3(vertical_tile_7_13_to_tile_6_13_3),
		.out_wire_2_0(horizontal_tile_6_13_to_tile_6_12_0),
		.out_wire_2_1(horizontal_tile_6_13_to_tile_6_12_1),
		.out_wire_2_2(horizontal_tile_6_13_to_tile_6_12_2),
		.out_wire_2_3(horizontal_tile_6_13_to_tile_6_12_3),
		.in_wire_2_0(horizontal_tile_6_12_to_tile_6_13_0),
		.in_wire_2_1(horizontal_tile_6_12_to_tile_6_13_1),
		.in_wire_2_2(horizontal_tile_6_12_to_tile_6_13_2),
		.in_wire_2_3(horizontal_tile_6_12_to_tile_6_13_3),
		.out_wire_0_0(horizontal_tile_6_13_to_tile_6_14_0),
		.out_wire_0_1(horizontal_tile_6_13_to_tile_6_14_1),
		.out_wire_0_2(horizontal_tile_6_13_to_tile_6_14_2),
		.out_wire_0_3(horizontal_tile_6_13_to_tile_6_14_3),
		.in_wire_0_0(horizontal_tile_6_14_to_tile_6_13_0),
		.in_wire_0_1(horizontal_tile_6_14_to_tile_6_13_1),
		.in_wire_0_2(horizontal_tile_6_14_to_tile_6_13_2),
		.in_wire_0_3(horizontal_tile_6_14_to_tile_6_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(206)
	);

	pe_tile pe_tile_6_14(
		.out_wire_3_0(vertical_tile_6_14_to_tile_5_14_0),
		.out_wire_3_1(vertical_tile_6_14_to_tile_5_14_1),
		.out_wire_3_2(vertical_tile_6_14_to_tile_5_14_2),
		.out_wire_3_3(vertical_tile_6_14_to_tile_5_14_3),
		.in_wire_3_0(vertical_tile_5_14_to_tile_6_14_0),
		.in_wire_3_1(vertical_tile_5_14_to_tile_6_14_1),
		.in_wire_3_2(vertical_tile_5_14_to_tile_6_14_2),
		.in_wire_3_3(vertical_tile_5_14_to_tile_6_14_3),
		.out_wire_1_0(vertical_tile_6_14_to_tile_7_14_0),
		.out_wire_1_1(vertical_tile_6_14_to_tile_7_14_1),
		.out_wire_1_2(vertical_tile_6_14_to_tile_7_14_2),
		.out_wire_1_3(vertical_tile_6_14_to_tile_7_14_3),
		.in_wire_1_0(vertical_tile_7_14_to_tile_6_14_0),
		.in_wire_1_1(vertical_tile_7_14_to_tile_6_14_1),
		.in_wire_1_2(vertical_tile_7_14_to_tile_6_14_2),
		.in_wire_1_3(vertical_tile_7_14_to_tile_6_14_3),
		.out_wire_2_0(horizontal_tile_6_14_to_tile_6_13_0),
		.out_wire_2_1(horizontal_tile_6_14_to_tile_6_13_1),
		.out_wire_2_2(horizontal_tile_6_14_to_tile_6_13_2),
		.out_wire_2_3(horizontal_tile_6_14_to_tile_6_13_3),
		.in_wire_2_0(horizontal_tile_6_13_to_tile_6_14_0),
		.in_wire_2_1(horizontal_tile_6_13_to_tile_6_14_1),
		.in_wire_2_2(horizontal_tile_6_13_to_tile_6_14_2),
		.in_wire_2_3(horizontal_tile_6_13_to_tile_6_14_3),
		.out_wire_0_0(horizontal_tile_6_14_to_tile_6_15_0),
		.out_wire_0_1(horizontal_tile_6_14_to_tile_6_15_1),
		.out_wire_0_2(horizontal_tile_6_14_to_tile_6_15_2),
		.out_wire_0_3(horizontal_tile_6_14_to_tile_6_15_3),
		.in_wire_0_0(horizontal_tile_6_15_to_tile_6_14_0),
		.in_wire_0_1(horizontal_tile_6_15_to_tile_6_14_1),
		.in_wire_0_2(horizontal_tile_6_15_to_tile_6_14_2),
		.in_wire_0_3(horizontal_tile_6_15_to_tile_6_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(207)
	);

	pe_tile pe_tile_6_15(
		.out_wire_3_0(vertical_tile_6_15_to_tile_5_15_0),
		.out_wire_3_1(vertical_tile_6_15_to_tile_5_15_1),
		.out_wire_3_2(vertical_tile_6_15_to_tile_5_15_2),
		.out_wire_3_3(vertical_tile_6_15_to_tile_5_15_3),
		.in_wire_3_0(vertical_tile_5_15_to_tile_6_15_0),
		.in_wire_3_1(vertical_tile_5_15_to_tile_6_15_1),
		.in_wire_3_2(vertical_tile_5_15_to_tile_6_15_2),
		.in_wire_3_3(vertical_tile_5_15_to_tile_6_15_3),
		.out_wire_1_0(vertical_tile_6_15_to_tile_7_15_0),
		.out_wire_1_1(vertical_tile_6_15_to_tile_7_15_1),
		.out_wire_1_2(vertical_tile_6_15_to_tile_7_15_2),
		.out_wire_1_3(vertical_tile_6_15_to_tile_7_15_3),
		.in_wire_1_0(vertical_tile_7_15_to_tile_6_15_0),
		.in_wire_1_1(vertical_tile_7_15_to_tile_6_15_1),
		.in_wire_1_2(vertical_tile_7_15_to_tile_6_15_2),
		.in_wire_1_3(vertical_tile_7_15_to_tile_6_15_3),
		.out_wire_2_0(horizontal_tile_6_15_to_tile_6_14_0),
		.out_wire_2_1(horizontal_tile_6_15_to_tile_6_14_1),
		.out_wire_2_2(horizontal_tile_6_15_to_tile_6_14_2),
		.out_wire_2_3(horizontal_tile_6_15_to_tile_6_14_3),
		.in_wire_2_0(horizontal_tile_6_14_to_tile_6_15_0),
		.in_wire_2_1(horizontal_tile_6_14_to_tile_6_15_1),
		.in_wire_2_2(horizontal_tile_6_14_to_tile_6_15_2),
		.in_wire_2_3(horizontal_tile_6_14_to_tile_6_15_3),
		.out_wire_0_0(horizontal_tile_6_15_to_tile_6_16_0),
		.out_wire_0_1(horizontal_tile_6_15_to_tile_6_16_1),
		.out_wire_0_2(horizontal_tile_6_15_to_tile_6_16_2),
		.out_wire_0_3(horizontal_tile_6_15_to_tile_6_16_3),
		.in_wire_0_0(horizontal_tile_6_16_to_tile_6_15_0),
		.in_wire_0_1(horizontal_tile_6_16_to_tile_6_15_1),
		.in_wire_0_2(horizontal_tile_6_16_to_tile_6_15_2),
		.in_wire_0_3(horizontal_tile_6_16_to_tile_6_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(208)
	);

	pe_tile pe_tile_6_16(
		.out_wire_3_0(vertical_tile_6_16_to_tile_5_16_0),
		.out_wire_3_1(vertical_tile_6_16_to_tile_5_16_1),
		.out_wire_3_2(vertical_tile_6_16_to_tile_5_16_2),
		.out_wire_3_3(vertical_tile_6_16_to_tile_5_16_3),
		.in_wire_3_0(vertical_tile_5_16_to_tile_6_16_0),
		.in_wire_3_1(vertical_tile_5_16_to_tile_6_16_1),
		.in_wire_3_2(vertical_tile_5_16_to_tile_6_16_2),
		.in_wire_3_3(vertical_tile_5_16_to_tile_6_16_3),
		.out_wire_1_0(vertical_tile_6_16_to_tile_7_16_0),
		.out_wire_1_1(vertical_tile_6_16_to_tile_7_16_1),
		.out_wire_1_2(vertical_tile_6_16_to_tile_7_16_2),
		.out_wire_1_3(vertical_tile_6_16_to_tile_7_16_3),
		.in_wire_1_0(vertical_tile_7_16_to_tile_6_16_0),
		.in_wire_1_1(vertical_tile_7_16_to_tile_6_16_1),
		.in_wire_1_2(vertical_tile_7_16_to_tile_6_16_2),
		.in_wire_1_3(vertical_tile_7_16_to_tile_6_16_3),
		.out_wire_2_0(horizontal_tile_6_16_to_tile_6_15_0),
		.out_wire_2_1(horizontal_tile_6_16_to_tile_6_15_1),
		.out_wire_2_2(horizontal_tile_6_16_to_tile_6_15_2),
		.out_wire_2_3(horizontal_tile_6_16_to_tile_6_15_3),
		.in_wire_2_0(horizontal_tile_6_15_to_tile_6_16_0),
		.in_wire_2_1(horizontal_tile_6_15_to_tile_6_16_1),
		.in_wire_2_2(horizontal_tile_6_15_to_tile_6_16_2),
		.in_wire_2_3(horizontal_tile_6_15_to_tile_6_16_3),
		.out_wire_0_0(horizontal_tile_6_16_to_tile_6_17_0),
		.out_wire_0_1(horizontal_tile_6_16_to_tile_6_17_1),
		.out_wire_0_2(horizontal_tile_6_16_to_tile_6_17_2),
		.out_wire_0_3(horizontal_tile_6_16_to_tile_6_17_3),
		.in_wire_0_0(horizontal_tile_6_17_to_tile_6_16_0),
		.in_wire_0_1(horizontal_tile_6_17_to_tile_6_16_1),
		.in_wire_0_2(horizontal_tile_6_17_to_tile_6_16_2),
		.in_wire_0_3(horizontal_tile_6_17_to_tile_6_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(209)
	);

	pe_tile pe_tile_6_17(
		.out_wire_3_0(vertical_tile_6_17_to_tile_5_17_0),
		.out_wire_3_1(vertical_tile_6_17_to_tile_5_17_1),
		.out_wire_3_2(vertical_tile_6_17_to_tile_5_17_2),
		.out_wire_3_3(vertical_tile_6_17_to_tile_5_17_3),
		.in_wire_3_0(vertical_tile_5_17_to_tile_6_17_0),
		.in_wire_3_1(vertical_tile_5_17_to_tile_6_17_1),
		.in_wire_3_2(vertical_tile_5_17_to_tile_6_17_2),
		.in_wire_3_3(vertical_tile_5_17_to_tile_6_17_3),
		.out_wire_1_0(vertical_tile_6_17_to_tile_7_17_0),
		.out_wire_1_1(vertical_tile_6_17_to_tile_7_17_1),
		.out_wire_1_2(vertical_tile_6_17_to_tile_7_17_2),
		.out_wire_1_3(vertical_tile_6_17_to_tile_7_17_3),
		.in_wire_1_0(vertical_tile_7_17_to_tile_6_17_0),
		.in_wire_1_1(vertical_tile_7_17_to_tile_6_17_1),
		.in_wire_1_2(vertical_tile_7_17_to_tile_6_17_2),
		.in_wire_1_3(vertical_tile_7_17_to_tile_6_17_3),
		.out_wire_2_0(horizontal_tile_6_17_to_tile_6_16_0),
		.out_wire_2_1(horizontal_tile_6_17_to_tile_6_16_1),
		.out_wire_2_2(horizontal_tile_6_17_to_tile_6_16_2),
		.out_wire_2_3(horizontal_tile_6_17_to_tile_6_16_3),
		.in_wire_2_0(horizontal_tile_6_16_to_tile_6_17_0),
		.in_wire_2_1(horizontal_tile_6_16_to_tile_6_17_1),
		.in_wire_2_2(horizontal_tile_6_16_to_tile_6_17_2),
		.in_wire_2_3(horizontal_tile_6_16_to_tile_6_17_3),
		.out_wire_0_0(horizontal_tile_6_17_to_tile_6_18_0),
		.out_wire_0_1(horizontal_tile_6_17_to_tile_6_18_1),
		.out_wire_0_2(horizontal_tile_6_17_to_tile_6_18_2),
		.out_wire_0_3(horizontal_tile_6_17_to_tile_6_18_3),
		.in_wire_0_0(horizontal_tile_6_18_to_tile_6_17_0),
		.in_wire_0_1(horizontal_tile_6_18_to_tile_6_17_1),
		.in_wire_0_2(horizontal_tile_6_18_to_tile_6_17_2),
		.in_wire_0_3(horizontal_tile_6_18_to_tile_6_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(210)
	);

	pe_tile pe_tile_6_18(
		.out_wire_3_0(vertical_tile_6_18_to_tile_5_18_0),
		.out_wire_3_1(vertical_tile_6_18_to_tile_5_18_1),
		.out_wire_3_2(vertical_tile_6_18_to_tile_5_18_2),
		.out_wire_3_3(vertical_tile_6_18_to_tile_5_18_3),
		.in_wire_3_0(vertical_tile_5_18_to_tile_6_18_0),
		.in_wire_3_1(vertical_tile_5_18_to_tile_6_18_1),
		.in_wire_3_2(vertical_tile_5_18_to_tile_6_18_2),
		.in_wire_3_3(vertical_tile_5_18_to_tile_6_18_3),
		.out_wire_1_0(vertical_tile_6_18_to_tile_7_18_0),
		.out_wire_1_1(vertical_tile_6_18_to_tile_7_18_1),
		.out_wire_1_2(vertical_tile_6_18_to_tile_7_18_2),
		.out_wire_1_3(vertical_tile_6_18_to_tile_7_18_3),
		.in_wire_1_0(vertical_tile_7_18_to_tile_6_18_0),
		.in_wire_1_1(vertical_tile_7_18_to_tile_6_18_1),
		.in_wire_1_2(vertical_tile_7_18_to_tile_6_18_2),
		.in_wire_1_3(vertical_tile_7_18_to_tile_6_18_3),
		.out_wire_2_0(horizontal_tile_6_18_to_tile_6_17_0),
		.out_wire_2_1(horizontal_tile_6_18_to_tile_6_17_1),
		.out_wire_2_2(horizontal_tile_6_18_to_tile_6_17_2),
		.out_wire_2_3(horizontal_tile_6_18_to_tile_6_17_3),
		.in_wire_2_0(horizontal_tile_6_17_to_tile_6_18_0),
		.in_wire_2_1(horizontal_tile_6_17_to_tile_6_18_1),
		.in_wire_2_2(horizontal_tile_6_17_to_tile_6_18_2),
		.in_wire_2_3(horizontal_tile_6_17_to_tile_6_18_3),
		.out_wire_0_0(horizontal_tile_6_18_to_tile_6_19_0),
		.out_wire_0_1(horizontal_tile_6_18_to_tile_6_19_1),
		.out_wire_0_2(horizontal_tile_6_18_to_tile_6_19_2),
		.out_wire_0_3(horizontal_tile_6_18_to_tile_6_19_3),
		.in_wire_0_0(horizontal_tile_6_19_to_tile_6_18_0),
		.in_wire_0_1(horizontal_tile_6_19_to_tile_6_18_1),
		.in_wire_0_2(horizontal_tile_6_19_to_tile_6_18_2),
		.in_wire_0_3(horizontal_tile_6_19_to_tile_6_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(211)
	);

	pe_tile pe_tile_6_19(
		.out_wire_3_0(vertical_tile_6_19_to_tile_5_19_0),
		.out_wire_3_1(vertical_tile_6_19_to_tile_5_19_1),
		.out_wire_3_2(vertical_tile_6_19_to_tile_5_19_2),
		.out_wire_3_3(vertical_tile_6_19_to_tile_5_19_3),
		.in_wire_3_0(vertical_tile_5_19_to_tile_6_19_0),
		.in_wire_3_1(vertical_tile_5_19_to_tile_6_19_1),
		.in_wire_3_2(vertical_tile_5_19_to_tile_6_19_2),
		.in_wire_3_3(vertical_tile_5_19_to_tile_6_19_3),
		.out_wire_1_0(vertical_tile_6_19_to_tile_7_19_0),
		.out_wire_1_1(vertical_tile_6_19_to_tile_7_19_1),
		.out_wire_1_2(vertical_tile_6_19_to_tile_7_19_2),
		.out_wire_1_3(vertical_tile_6_19_to_tile_7_19_3),
		.in_wire_1_0(vertical_tile_7_19_to_tile_6_19_0),
		.in_wire_1_1(vertical_tile_7_19_to_tile_6_19_1),
		.in_wire_1_2(vertical_tile_7_19_to_tile_6_19_2),
		.in_wire_1_3(vertical_tile_7_19_to_tile_6_19_3),
		.out_wire_2_0(horizontal_tile_6_19_to_tile_6_18_0),
		.out_wire_2_1(horizontal_tile_6_19_to_tile_6_18_1),
		.out_wire_2_2(horizontal_tile_6_19_to_tile_6_18_2),
		.out_wire_2_3(horizontal_tile_6_19_to_tile_6_18_3),
		.in_wire_2_0(horizontal_tile_6_18_to_tile_6_19_0),
		.in_wire_2_1(horizontal_tile_6_18_to_tile_6_19_1),
		.in_wire_2_2(horizontal_tile_6_18_to_tile_6_19_2),
		.in_wire_2_3(horizontal_tile_6_18_to_tile_6_19_3),
		.out_wire_0_0(horizontal_tile_6_19_to_tile_6_20_0),
		.out_wire_0_1(horizontal_tile_6_19_to_tile_6_20_1),
		.out_wire_0_2(horizontal_tile_6_19_to_tile_6_20_2),
		.out_wire_0_3(horizontal_tile_6_19_to_tile_6_20_3),
		.in_wire_0_0(horizontal_tile_6_20_to_tile_6_19_0),
		.in_wire_0_1(horizontal_tile_6_20_to_tile_6_19_1),
		.in_wire_0_2(horizontal_tile_6_20_to_tile_6_19_2),
		.in_wire_0_3(horizontal_tile_6_20_to_tile_6_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(212)
	);

	pe_tile pe_tile_6_20(
		.out_wire_3_0(vertical_tile_6_20_to_tile_5_20_0),
		.out_wire_3_1(vertical_tile_6_20_to_tile_5_20_1),
		.out_wire_3_2(vertical_tile_6_20_to_tile_5_20_2),
		.out_wire_3_3(vertical_tile_6_20_to_tile_5_20_3),
		.in_wire_3_0(vertical_tile_5_20_to_tile_6_20_0),
		.in_wire_3_1(vertical_tile_5_20_to_tile_6_20_1),
		.in_wire_3_2(vertical_tile_5_20_to_tile_6_20_2),
		.in_wire_3_3(vertical_tile_5_20_to_tile_6_20_3),
		.out_wire_1_0(vertical_tile_6_20_to_tile_7_20_0),
		.out_wire_1_1(vertical_tile_6_20_to_tile_7_20_1),
		.out_wire_1_2(vertical_tile_6_20_to_tile_7_20_2),
		.out_wire_1_3(vertical_tile_6_20_to_tile_7_20_3),
		.in_wire_1_0(vertical_tile_7_20_to_tile_6_20_0),
		.in_wire_1_1(vertical_tile_7_20_to_tile_6_20_1),
		.in_wire_1_2(vertical_tile_7_20_to_tile_6_20_2),
		.in_wire_1_3(vertical_tile_7_20_to_tile_6_20_3),
		.out_wire_2_0(horizontal_tile_6_20_to_tile_6_19_0),
		.out_wire_2_1(horizontal_tile_6_20_to_tile_6_19_1),
		.out_wire_2_2(horizontal_tile_6_20_to_tile_6_19_2),
		.out_wire_2_3(horizontal_tile_6_20_to_tile_6_19_3),
		.in_wire_2_0(horizontal_tile_6_19_to_tile_6_20_0),
		.in_wire_2_1(horizontal_tile_6_19_to_tile_6_20_1),
		.in_wire_2_2(horizontal_tile_6_19_to_tile_6_20_2),
		.in_wire_2_3(horizontal_tile_6_19_to_tile_6_20_3),
		.out_wire_0_0(horizontal_tile_6_20_to_tile_6_21_0),
		.out_wire_0_1(horizontal_tile_6_20_to_tile_6_21_1),
		.out_wire_0_2(horizontal_tile_6_20_to_tile_6_21_2),
		.out_wire_0_3(horizontal_tile_6_20_to_tile_6_21_3),
		.in_wire_0_0(horizontal_tile_6_21_to_tile_6_20_0),
		.in_wire_0_1(horizontal_tile_6_21_to_tile_6_20_1),
		.in_wire_0_2(horizontal_tile_6_21_to_tile_6_20_2),
		.in_wire_0_3(horizontal_tile_6_21_to_tile_6_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(213)
	);

	pe_tile pe_tile_6_21(
		.out_wire_3_0(vertical_tile_6_21_to_tile_5_21_0),
		.out_wire_3_1(vertical_tile_6_21_to_tile_5_21_1),
		.out_wire_3_2(vertical_tile_6_21_to_tile_5_21_2),
		.out_wire_3_3(vertical_tile_6_21_to_tile_5_21_3),
		.in_wire_3_0(vertical_tile_5_21_to_tile_6_21_0),
		.in_wire_3_1(vertical_tile_5_21_to_tile_6_21_1),
		.in_wire_3_2(vertical_tile_5_21_to_tile_6_21_2),
		.in_wire_3_3(vertical_tile_5_21_to_tile_6_21_3),
		.out_wire_1_0(vertical_tile_6_21_to_tile_7_21_0),
		.out_wire_1_1(vertical_tile_6_21_to_tile_7_21_1),
		.out_wire_1_2(vertical_tile_6_21_to_tile_7_21_2),
		.out_wire_1_3(vertical_tile_6_21_to_tile_7_21_3),
		.in_wire_1_0(vertical_tile_7_21_to_tile_6_21_0),
		.in_wire_1_1(vertical_tile_7_21_to_tile_6_21_1),
		.in_wire_1_2(vertical_tile_7_21_to_tile_6_21_2),
		.in_wire_1_3(vertical_tile_7_21_to_tile_6_21_3),
		.out_wire_2_0(horizontal_tile_6_21_to_tile_6_20_0),
		.out_wire_2_1(horizontal_tile_6_21_to_tile_6_20_1),
		.out_wire_2_2(horizontal_tile_6_21_to_tile_6_20_2),
		.out_wire_2_3(horizontal_tile_6_21_to_tile_6_20_3),
		.in_wire_2_0(horizontal_tile_6_20_to_tile_6_21_0),
		.in_wire_2_1(horizontal_tile_6_20_to_tile_6_21_1),
		.in_wire_2_2(horizontal_tile_6_20_to_tile_6_21_2),
		.in_wire_2_3(horizontal_tile_6_20_to_tile_6_21_3),
		.out_wire_0_0(horizontal_tile_6_21_to_tile_6_22_0),
		.out_wire_0_1(horizontal_tile_6_21_to_tile_6_22_1),
		.out_wire_0_2(horizontal_tile_6_21_to_tile_6_22_2),
		.out_wire_0_3(horizontal_tile_6_21_to_tile_6_22_3),
		.in_wire_0_0(horizontal_tile_6_22_to_tile_6_21_0),
		.in_wire_0_1(horizontal_tile_6_22_to_tile_6_21_1),
		.in_wire_0_2(horizontal_tile_6_22_to_tile_6_21_2),
		.in_wire_0_3(horizontal_tile_6_22_to_tile_6_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(214)
	);

	pe_tile pe_tile_6_22(
		.out_wire_3_0(vertical_tile_6_22_to_tile_5_22_0),
		.out_wire_3_1(vertical_tile_6_22_to_tile_5_22_1),
		.out_wire_3_2(vertical_tile_6_22_to_tile_5_22_2),
		.out_wire_3_3(vertical_tile_6_22_to_tile_5_22_3),
		.in_wire_3_0(vertical_tile_5_22_to_tile_6_22_0),
		.in_wire_3_1(vertical_tile_5_22_to_tile_6_22_1),
		.in_wire_3_2(vertical_tile_5_22_to_tile_6_22_2),
		.in_wire_3_3(vertical_tile_5_22_to_tile_6_22_3),
		.out_wire_1_0(vertical_tile_6_22_to_tile_7_22_0),
		.out_wire_1_1(vertical_tile_6_22_to_tile_7_22_1),
		.out_wire_1_2(vertical_tile_6_22_to_tile_7_22_2),
		.out_wire_1_3(vertical_tile_6_22_to_tile_7_22_3),
		.in_wire_1_0(vertical_tile_7_22_to_tile_6_22_0),
		.in_wire_1_1(vertical_tile_7_22_to_tile_6_22_1),
		.in_wire_1_2(vertical_tile_7_22_to_tile_6_22_2),
		.in_wire_1_3(vertical_tile_7_22_to_tile_6_22_3),
		.out_wire_2_0(horizontal_tile_6_22_to_tile_6_21_0),
		.out_wire_2_1(horizontal_tile_6_22_to_tile_6_21_1),
		.out_wire_2_2(horizontal_tile_6_22_to_tile_6_21_2),
		.out_wire_2_3(horizontal_tile_6_22_to_tile_6_21_3),
		.in_wire_2_0(horizontal_tile_6_21_to_tile_6_22_0),
		.in_wire_2_1(horizontal_tile_6_21_to_tile_6_22_1),
		.in_wire_2_2(horizontal_tile_6_21_to_tile_6_22_2),
		.in_wire_2_3(horizontal_tile_6_21_to_tile_6_22_3),
		.out_wire_0_0(horizontal_tile_6_22_to_tile_6_23_0),
		.out_wire_0_1(horizontal_tile_6_22_to_tile_6_23_1),
		.out_wire_0_2(horizontal_tile_6_22_to_tile_6_23_2),
		.out_wire_0_3(horizontal_tile_6_22_to_tile_6_23_3),
		.in_wire_0_0(horizontal_tile_6_23_to_tile_6_22_0),
		.in_wire_0_1(horizontal_tile_6_23_to_tile_6_22_1),
		.in_wire_0_2(horizontal_tile_6_23_to_tile_6_22_2),
		.in_wire_0_3(horizontal_tile_6_23_to_tile_6_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(215)
	);

	pe_tile pe_tile_6_23(
		.out_wire_3_0(vertical_tile_6_23_to_tile_5_23_0),
		.out_wire_3_1(vertical_tile_6_23_to_tile_5_23_1),
		.out_wire_3_2(vertical_tile_6_23_to_tile_5_23_2),
		.out_wire_3_3(vertical_tile_6_23_to_tile_5_23_3),
		.in_wire_3_0(vertical_tile_5_23_to_tile_6_23_0),
		.in_wire_3_1(vertical_tile_5_23_to_tile_6_23_1),
		.in_wire_3_2(vertical_tile_5_23_to_tile_6_23_2),
		.in_wire_3_3(vertical_tile_5_23_to_tile_6_23_3),
		.out_wire_1_0(vertical_tile_6_23_to_tile_7_23_0),
		.out_wire_1_1(vertical_tile_6_23_to_tile_7_23_1),
		.out_wire_1_2(vertical_tile_6_23_to_tile_7_23_2),
		.out_wire_1_3(vertical_tile_6_23_to_tile_7_23_3),
		.in_wire_1_0(vertical_tile_7_23_to_tile_6_23_0),
		.in_wire_1_1(vertical_tile_7_23_to_tile_6_23_1),
		.in_wire_1_2(vertical_tile_7_23_to_tile_6_23_2),
		.in_wire_1_3(vertical_tile_7_23_to_tile_6_23_3),
		.out_wire_2_0(horizontal_tile_6_23_to_tile_6_22_0),
		.out_wire_2_1(horizontal_tile_6_23_to_tile_6_22_1),
		.out_wire_2_2(horizontal_tile_6_23_to_tile_6_22_2),
		.out_wire_2_3(horizontal_tile_6_23_to_tile_6_22_3),
		.in_wire_2_0(horizontal_tile_6_22_to_tile_6_23_0),
		.in_wire_2_1(horizontal_tile_6_22_to_tile_6_23_1),
		.in_wire_2_2(horizontal_tile_6_22_to_tile_6_23_2),
		.in_wire_2_3(horizontal_tile_6_22_to_tile_6_23_3),
		.out_wire_0_0(horizontal_tile_6_23_to_tile_6_24_0),
		.out_wire_0_1(horizontal_tile_6_23_to_tile_6_24_1),
		.out_wire_0_2(horizontal_tile_6_23_to_tile_6_24_2),
		.out_wire_0_3(horizontal_tile_6_23_to_tile_6_24_3),
		.in_wire_0_0(horizontal_tile_6_24_to_tile_6_23_0),
		.in_wire_0_1(horizontal_tile_6_24_to_tile_6_23_1),
		.in_wire_0_2(horizontal_tile_6_24_to_tile_6_23_2),
		.in_wire_0_3(horizontal_tile_6_24_to_tile_6_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(216)
	);

	pe_tile pe_tile_6_24(
		.out_wire_3_0(vertical_tile_6_24_to_tile_5_24_0),
		.out_wire_3_1(vertical_tile_6_24_to_tile_5_24_1),
		.out_wire_3_2(vertical_tile_6_24_to_tile_5_24_2),
		.out_wire_3_3(vertical_tile_6_24_to_tile_5_24_3),
		.in_wire_3_0(vertical_tile_5_24_to_tile_6_24_0),
		.in_wire_3_1(vertical_tile_5_24_to_tile_6_24_1),
		.in_wire_3_2(vertical_tile_5_24_to_tile_6_24_2),
		.in_wire_3_3(vertical_tile_5_24_to_tile_6_24_3),
		.out_wire_1_0(vertical_tile_6_24_to_tile_7_24_0),
		.out_wire_1_1(vertical_tile_6_24_to_tile_7_24_1),
		.out_wire_1_2(vertical_tile_6_24_to_tile_7_24_2),
		.out_wire_1_3(vertical_tile_6_24_to_tile_7_24_3),
		.in_wire_1_0(vertical_tile_7_24_to_tile_6_24_0),
		.in_wire_1_1(vertical_tile_7_24_to_tile_6_24_1),
		.in_wire_1_2(vertical_tile_7_24_to_tile_6_24_2),
		.in_wire_1_3(vertical_tile_7_24_to_tile_6_24_3),
		.out_wire_2_0(horizontal_tile_6_24_to_tile_6_23_0),
		.out_wire_2_1(horizontal_tile_6_24_to_tile_6_23_1),
		.out_wire_2_2(horizontal_tile_6_24_to_tile_6_23_2),
		.out_wire_2_3(horizontal_tile_6_24_to_tile_6_23_3),
		.in_wire_2_0(horizontal_tile_6_23_to_tile_6_24_0),
		.in_wire_2_1(horizontal_tile_6_23_to_tile_6_24_1),
		.in_wire_2_2(horizontal_tile_6_23_to_tile_6_24_2),
		.in_wire_2_3(horizontal_tile_6_23_to_tile_6_24_3),
		.out_wire_0_0(horizontal_tile_6_24_to_tile_6_25_0),
		.out_wire_0_1(horizontal_tile_6_24_to_tile_6_25_1),
		.out_wire_0_2(horizontal_tile_6_24_to_tile_6_25_2),
		.out_wire_0_3(horizontal_tile_6_24_to_tile_6_25_3),
		.in_wire_0_0(horizontal_tile_6_25_to_tile_6_24_0),
		.in_wire_0_1(horizontal_tile_6_25_to_tile_6_24_1),
		.in_wire_0_2(horizontal_tile_6_25_to_tile_6_24_2),
		.in_wire_0_3(horizontal_tile_6_25_to_tile_6_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(217)
	);

	pe_tile pe_tile_6_25(
		.out_wire_3_0(vertical_tile_6_25_to_tile_5_25_0),
		.out_wire_3_1(vertical_tile_6_25_to_tile_5_25_1),
		.out_wire_3_2(vertical_tile_6_25_to_tile_5_25_2),
		.out_wire_3_3(vertical_tile_6_25_to_tile_5_25_3),
		.in_wire_3_0(vertical_tile_5_25_to_tile_6_25_0),
		.in_wire_3_1(vertical_tile_5_25_to_tile_6_25_1),
		.in_wire_3_2(vertical_tile_5_25_to_tile_6_25_2),
		.in_wire_3_3(vertical_tile_5_25_to_tile_6_25_3),
		.out_wire_1_0(vertical_tile_6_25_to_tile_7_25_0),
		.out_wire_1_1(vertical_tile_6_25_to_tile_7_25_1),
		.out_wire_1_2(vertical_tile_6_25_to_tile_7_25_2),
		.out_wire_1_3(vertical_tile_6_25_to_tile_7_25_3),
		.in_wire_1_0(vertical_tile_7_25_to_tile_6_25_0),
		.in_wire_1_1(vertical_tile_7_25_to_tile_6_25_1),
		.in_wire_1_2(vertical_tile_7_25_to_tile_6_25_2),
		.in_wire_1_3(vertical_tile_7_25_to_tile_6_25_3),
		.out_wire_2_0(horizontal_tile_6_25_to_tile_6_24_0),
		.out_wire_2_1(horizontal_tile_6_25_to_tile_6_24_1),
		.out_wire_2_2(horizontal_tile_6_25_to_tile_6_24_2),
		.out_wire_2_3(horizontal_tile_6_25_to_tile_6_24_3),
		.in_wire_2_0(horizontal_tile_6_24_to_tile_6_25_0),
		.in_wire_2_1(horizontal_tile_6_24_to_tile_6_25_1),
		.in_wire_2_2(horizontal_tile_6_24_to_tile_6_25_2),
		.in_wire_2_3(horizontal_tile_6_24_to_tile_6_25_3),
		.out_wire_0_0(horizontal_tile_6_25_to_tile_6_26_0),
		.out_wire_0_1(horizontal_tile_6_25_to_tile_6_26_1),
		.out_wire_0_2(horizontal_tile_6_25_to_tile_6_26_2),
		.out_wire_0_3(horizontal_tile_6_25_to_tile_6_26_3),
		.in_wire_0_0(horizontal_tile_6_26_to_tile_6_25_0),
		.in_wire_0_1(horizontal_tile_6_26_to_tile_6_25_1),
		.in_wire_0_2(horizontal_tile_6_26_to_tile_6_25_2),
		.in_wire_0_3(horizontal_tile_6_26_to_tile_6_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(218)
	);

	pe_tile pe_tile_6_26(
		.out_wire_3_0(vertical_tile_6_26_to_tile_5_26_0),
		.out_wire_3_1(vertical_tile_6_26_to_tile_5_26_1),
		.out_wire_3_2(vertical_tile_6_26_to_tile_5_26_2),
		.out_wire_3_3(vertical_tile_6_26_to_tile_5_26_3),
		.in_wire_3_0(vertical_tile_5_26_to_tile_6_26_0),
		.in_wire_3_1(vertical_tile_5_26_to_tile_6_26_1),
		.in_wire_3_2(vertical_tile_5_26_to_tile_6_26_2),
		.in_wire_3_3(vertical_tile_5_26_to_tile_6_26_3),
		.out_wire_1_0(vertical_tile_6_26_to_tile_7_26_0),
		.out_wire_1_1(vertical_tile_6_26_to_tile_7_26_1),
		.out_wire_1_2(vertical_tile_6_26_to_tile_7_26_2),
		.out_wire_1_3(vertical_tile_6_26_to_tile_7_26_3),
		.in_wire_1_0(vertical_tile_7_26_to_tile_6_26_0),
		.in_wire_1_1(vertical_tile_7_26_to_tile_6_26_1),
		.in_wire_1_2(vertical_tile_7_26_to_tile_6_26_2),
		.in_wire_1_3(vertical_tile_7_26_to_tile_6_26_3),
		.out_wire_2_0(horizontal_tile_6_26_to_tile_6_25_0),
		.out_wire_2_1(horizontal_tile_6_26_to_tile_6_25_1),
		.out_wire_2_2(horizontal_tile_6_26_to_tile_6_25_2),
		.out_wire_2_3(horizontal_tile_6_26_to_tile_6_25_3),
		.in_wire_2_0(horizontal_tile_6_25_to_tile_6_26_0),
		.in_wire_2_1(horizontal_tile_6_25_to_tile_6_26_1),
		.in_wire_2_2(horizontal_tile_6_25_to_tile_6_26_2),
		.in_wire_2_3(horizontal_tile_6_25_to_tile_6_26_3),
		.out_wire_0_0(horizontal_tile_6_26_to_tile_6_27_0),
		.out_wire_0_1(horizontal_tile_6_26_to_tile_6_27_1),
		.out_wire_0_2(horizontal_tile_6_26_to_tile_6_27_2),
		.out_wire_0_3(horizontal_tile_6_26_to_tile_6_27_3),
		.in_wire_0_0(horizontal_tile_6_27_to_tile_6_26_0),
		.in_wire_0_1(horizontal_tile_6_27_to_tile_6_26_1),
		.in_wire_0_2(horizontal_tile_6_27_to_tile_6_26_2),
		.in_wire_0_3(horizontal_tile_6_27_to_tile_6_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(219)
	);

	pe_tile pe_tile_6_27(
		.out_wire_3_0(vertical_tile_6_27_to_tile_5_27_0),
		.out_wire_3_1(vertical_tile_6_27_to_tile_5_27_1),
		.out_wire_3_2(vertical_tile_6_27_to_tile_5_27_2),
		.out_wire_3_3(vertical_tile_6_27_to_tile_5_27_3),
		.in_wire_3_0(vertical_tile_5_27_to_tile_6_27_0),
		.in_wire_3_1(vertical_tile_5_27_to_tile_6_27_1),
		.in_wire_3_2(vertical_tile_5_27_to_tile_6_27_2),
		.in_wire_3_3(vertical_tile_5_27_to_tile_6_27_3),
		.out_wire_1_0(vertical_tile_6_27_to_tile_7_27_0),
		.out_wire_1_1(vertical_tile_6_27_to_tile_7_27_1),
		.out_wire_1_2(vertical_tile_6_27_to_tile_7_27_2),
		.out_wire_1_3(vertical_tile_6_27_to_tile_7_27_3),
		.in_wire_1_0(vertical_tile_7_27_to_tile_6_27_0),
		.in_wire_1_1(vertical_tile_7_27_to_tile_6_27_1),
		.in_wire_1_2(vertical_tile_7_27_to_tile_6_27_2),
		.in_wire_1_3(vertical_tile_7_27_to_tile_6_27_3),
		.out_wire_2_0(horizontal_tile_6_27_to_tile_6_26_0),
		.out_wire_2_1(horizontal_tile_6_27_to_tile_6_26_1),
		.out_wire_2_2(horizontal_tile_6_27_to_tile_6_26_2),
		.out_wire_2_3(horizontal_tile_6_27_to_tile_6_26_3),
		.in_wire_2_0(horizontal_tile_6_26_to_tile_6_27_0),
		.in_wire_2_1(horizontal_tile_6_26_to_tile_6_27_1),
		.in_wire_2_2(horizontal_tile_6_26_to_tile_6_27_2),
		.in_wire_2_3(horizontal_tile_6_26_to_tile_6_27_3),
		.out_wire_0_0(horizontal_tile_6_27_to_tile_6_28_0),
		.out_wire_0_1(horizontal_tile_6_27_to_tile_6_28_1),
		.out_wire_0_2(horizontal_tile_6_27_to_tile_6_28_2),
		.out_wire_0_3(horizontal_tile_6_27_to_tile_6_28_3),
		.in_wire_0_0(horizontal_tile_6_28_to_tile_6_27_0),
		.in_wire_0_1(horizontal_tile_6_28_to_tile_6_27_1),
		.in_wire_0_2(horizontal_tile_6_28_to_tile_6_27_2),
		.in_wire_0_3(horizontal_tile_6_28_to_tile_6_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(220)
	);

	pe_tile pe_tile_6_28(
		.out_wire_3_0(vertical_tile_6_28_to_tile_5_28_0),
		.out_wire_3_1(vertical_tile_6_28_to_tile_5_28_1),
		.out_wire_3_2(vertical_tile_6_28_to_tile_5_28_2),
		.out_wire_3_3(vertical_tile_6_28_to_tile_5_28_3),
		.in_wire_3_0(vertical_tile_5_28_to_tile_6_28_0),
		.in_wire_3_1(vertical_tile_5_28_to_tile_6_28_1),
		.in_wire_3_2(vertical_tile_5_28_to_tile_6_28_2),
		.in_wire_3_3(vertical_tile_5_28_to_tile_6_28_3),
		.out_wire_1_0(vertical_tile_6_28_to_tile_7_28_0),
		.out_wire_1_1(vertical_tile_6_28_to_tile_7_28_1),
		.out_wire_1_2(vertical_tile_6_28_to_tile_7_28_2),
		.out_wire_1_3(vertical_tile_6_28_to_tile_7_28_3),
		.in_wire_1_0(vertical_tile_7_28_to_tile_6_28_0),
		.in_wire_1_1(vertical_tile_7_28_to_tile_6_28_1),
		.in_wire_1_2(vertical_tile_7_28_to_tile_6_28_2),
		.in_wire_1_3(vertical_tile_7_28_to_tile_6_28_3),
		.out_wire_2_0(horizontal_tile_6_28_to_tile_6_27_0),
		.out_wire_2_1(horizontal_tile_6_28_to_tile_6_27_1),
		.out_wire_2_2(horizontal_tile_6_28_to_tile_6_27_2),
		.out_wire_2_3(horizontal_tile_6_28_to_tile_6_27_3),
		.in_wire_2_0(horizontal_tile_6_27_to_tile_6_28_0),
		.in_wire_2_1(horizontal_tile_6_27_to_tile_6_28_1),
		.in_wire_2_2(horizontal_tile_6_27_to_tile_6_28_2),
		.in_wire_2_3(horizontal_tile_6_27_to_tile_6_28_3),
		.out_wire_0_0(horizontal_tile_6_28_to_tile_6_29_0),
		.out_wire_0_1(horizontal_tile_6_28_to_tile_6_29_1),
		.out_wire_0_2(horizontal_tile_6_28_to_tile_6_29_2),
		.out_wire_0_3(horizontal_tile_6_28_to_tile_6_29_3),
		.in_wire_0_0(horizontal_tile_6_29_to_tile_6_28_0),
		.in_wire_0_1(horizontal_tile_6_29_to_tile_6_28_1),
		.in_wire_0_2(horizontal_tile_6_29_to_tile_6_28_2),
		.in_wire_0_3(horizontal_tile_6_29_to_tile_6_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(221)
	);

	pe_tile pe_tile_6_29(
		.out_wire_3_0(vertical_tile_6_29_to_tile_5_29_0),
		.out_wire_3_1(vertical_tile_6_29_to_tile_5_29_1),
		.out_wire_3_2(vertical_tile_6_29_to_tile_5_29_2),
		.out_wire_3_3(vertical_tile_6_29_to_tile_5_29_3),
		.in_wire_3_0(vertical_tile_5_29_to_tile_6_29_0),
		.in_wire_3_1(vertical_tile_5_29_to_tile_6_29_1),
		.in_wire_3_2(vertical_tile_5_29_to_tile_6_29_2),
		.in_wire_3_3(vertical_tile_5_29_to_tile_6_29_3),
		.out_wire_1_0(vertical_tile_6_29_to_tile_7_29_0),
		.out_wire_1_1(vertical_tile_6_29_to_tile_7_29_1),
		.out_wire_1_2(vertical_tile_6_29_to_tile_7_29_2),
		.out_wire_1_3(vertical_tile_6_29_to_tile_7_29_3),
		.in_wire_1_0(vertical_tile_7_29_to_tile_6_29_0),
		.in_wire_1_1(vertical_tile_7_29_to_tile_6_29_1),
		.in_wire_1_2(vertical_tile_7_29_to_tile_6_29_2),
		.in_wire_1_3(vertical_tile_7_29_to_tile_6_29_3),
		.out_wire_2_0(horizontal_tile_6_29_to_tile_6_28_0),
		.out_wire_2_1(horizontal_tile_6_29_to_tile_6_28_1),
		.out_wire_2_2(horizontal_tile_6_29_to_tile_6_28_2),
		.out_wire_2_3(horizontal_tile_6_29_to_tile_6_28_3),
		.in_wire_2_0(horizontal_tile_6_28_to_tile_6_29_0),
		.in_wire_2_1(horizontal_tile_6_28_to_tile_6_29_1),
		.in_wire_2_2(horizontal_tile_6_28_to_tile_6_29_2),
		.in_wire_2_3(horizontal_tile_6_28_to_tile_6_29_3),
		.out_wire_0_0(horizontal_tile_6_29_to_tile_6_30_0),
		.out_wire_0_1(horizontal_tile_6_29_to_tile_6_30_1),
		.out_wire_0_2(horizontal_tile_6_29_to_tile_6_30_2),
		.out_wire_0_3(horizontal_tile_6_29_to_tile_6_30_3),
		.in_wire_0_0(horizontal_tile_6_30_to_tile_6_29_0),
		.in_wire_0_1(horizontal_tile_6_30_to_tile_6_29_1),
		.in_wire_0_2(horizontal_tile_6_30_to_tile_6_29_2),
		.in_wire_0_3(horizontal_tile_6_30_to_tile_6_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(222)
	);

	pe_tile pe_tile_6_30(
		.out_wire_3_0(vertical_tile_6_30_to_tile_5_30_0),
		.out_wire_3_1(vertical_tile_6_30_to_tile_5_30_1),
		.out_wire_3_2(vertical_tile_6_30_to_tile_5_30_2),
		.out_wire_3_3(vertical_tile_6_30_to_tile_5_30_3),
		.in_wire_3_0(vertical_tile_5_30_to_tile_6_30_0),
		.in_wire_3_1(vertical_tile_5_30_to_tile_6_30_1),
		.in_wire_3_2(vertical_tile_5_30_to_tile_6_30_2),
		.in_wire_3_3(vertical_tile_5_30_to_tile_6_30_3),
		.out_wire_1_0(vertical_tile_6_30_to_tile_7_30_0),
		.out_wire_1_1(vertical_tile_6_30_to_tile_7_30_1),
		.out_wire_1_2(vertical_tile_6_30_to_tile_7_30_2),
		.out_wire_1_3(vertical_tile_6_30_to_tile_7_30_3),
		.in_wire_1_0(vertical_tile_7_30_to_tile_6_30_0),
		.in_wire_1_1(vertical_tile_7_30_to_tile_6_30_1),
		.in_wire_1_2(vertical_tile_7_30_to_tile_6_30_2),
		.in_wire_1_3(vertical_tile_7_30_to_tile_6_30_3),
		.out_wire_2_0(horizontal_tile_6_30_to_tile_6_29_0),
		.out_wire_2_1(horizontal_tile_6_30_to_tile_6_29_1),
		.out_wire_2_2(horizontal_tile_6_30_to_tile_6_29_2),
		.out_wire_2_3(horizontal_tile_6_30_to_tile_6_29_3),
		.in_wire_2_0(horizontal_tile_6_29_to_tile_6_30_0),
		.in_wire_2_1(horizontal_tile_6_29_to_tile_6_30_1),
		.in_wire_2_2(horizontal_tile_6_29_to_tile_6_30_2),
		.in_wire_2_3(horizontal_tile_6_29_to_tile_6_30_3),
		.out_wire_0_0(horizontal_tile_6_30_to_tile_6_31_0),
		.out_wire_0_1(horizontal_tile_6_30_to_tile_6_31_1),
		.out_wire_0_2(horizontal_tile_6_30_to_tile_6_31_2),
		.out_wire_0_3(horizontal_tile_6_30_to_tile_6_31_3),
		.in_wire_0_0(horizontal_tile_6_31_to_tile_6_30_0),
		.in_wire_0_1(horizontal_tile_6_31_to_tile_6_30_1),
		.in_wire_0_2(horizontal_tile_6_31_to_tile_6_30_2),
		.in_wire_0_3(horizontal_tile_6_31_to_tile_6_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(223)
	);

	pe_tile_right pe_tile_6_31(
		.out_wire_3_0(vertical_tile_6_31_to_tile_5_31_0),
		.out_wire_3_1(vertical_tile_6_31_to_tile_5_31_1),
		.out_wire_3_2(vertical_tile_6_31_to_tile_5_31_2),
		.out_wire_3_3(vertical_tile_6_31_to_tile_5_31_3),
		.in_wire_3_0(vertical_tile_5_31_to_tile_6_31_0),
		.in_wire_3_1(vertical_tile_5_31_to_tile_6_31_1),
		.in_wire_3_2(vertical_tile_5_31_to_tile_6_31_2),
		.in_wire_3_3(vertical_tile_5_31_to_tile_6_31_3),
		.out_wire_1_0(vertical_tile_6_31_to_tile_7_31_0),
		.out_wire_1_1(vertical_tile_6_31_to_tile_7_31_1),
		.out_wire_1_2(vertical_tile_6_31_to_tile_7_31_2),
		.out_wire_1_3(vertical_tile_6_31_to_tile_7_31_3),
		.in_wire_1_0(vertical_tile_7_31_to_tile_6_31_0),
		.in_wire_1_1(vertical_tile_7_31_to_tile_6_31_1),
		.in_wire_1_2(vertical_tile_7_31_to_tile_6_31_2),
		.in_wire_1_3(vertical_tile_7_31_to_tile_6_31_3),
		.out_wire_2_0(horizontal_tile_6_31_to_tile_6_30_0),
		.out_wire_2_1(horizontal_tile_6_31_to_tile_6_30_1),
		.out_wire_2_2(horizontal_tile_6_31_to_tile_6_30_2),
		.out_wire_2_3(horizontal_tile_6_31_to_tile_6_30_3),
		.in_wire_2_0(horizontal_tile_6_30_to_tile_6_31_0),
		.in_wire_2_1(horizontal_tile_6_30_to_tile_6_31_1),
		.in_wire_2_2(horizontal_tile_6_30_to_tile_6_31_2),
		.in_wire_2_3(horizontal_tile_6_30_to_tile_6_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(224)
	);

	pe_tile_left pe_tile_7_0(
		.out_wire_3_0(vertical_tile_7_0_to_tile_6_0_0),
		.out_wire_3_1(vertical_tile_7_0_to_tile_6_0_1),
		.out_wire_3_2(vertical_tile_7_0_to_tile_6_0_2),
		.out_wire_3_3(vertical_tile_7_0_to_tile_6_0_3),
		.in_wire_3_0(vertical_tile_6_0_to_tile_7_0_0),
		.in_wire_3_1(vertical_tile_6_0_to_tile_7_0_1),
		.in_wire_3_2(vertical_tile_6_0_to_tile_7_0_2),
		.in_wire_3_3(vertical_tile_6_0_to_tile_7_0_3),
		.out_wire_1_0(vertical_tile_7_0_to_tile_8_0_0),
		.out_wire_1_1(vertical_tile_7_0_to_tile_8_0_1),
		.out_wire_1_2(vertical_tile_7_0_to_tile_8_0_2),
		.out_wire_1_3(vertical_tile_7_0_to_tile_8_0_3),
		.in_wire_1_0(vertical_tile_8_0_to_tile_7_0_0),
		.in_wire_1_1(vertical_tile_8_0_to_tile_7_0_1),
		.in_wire_1_2(vertical_tile_8_0_to_tile_7_0_2),
		.in_wire_1_3(vertical_tile_8_0_to_tile_7_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_7_0_to_tile_7_1_0),
		.out_wire_0_1(horizontal_tile_7_0_to_tile_7_1_1),
		.out_wire_0_2(horizontal_tile_7_0_to_tile_7_1_2),
		.out_wire_0_3(horizontal_tile_7_0_to_tile_7_1_3),
		.in_wire_0_0(horizontal_tile_7_1_to_tile_7_0_0),
		.in_wire_0_1(horizontal_tile_7_1_to_tile_7_0_1),
		.in_wire_0_2(horizontal_tile_7_1_to_tile_7_0_2),
		.in_wire_0_3(horizontal_tile_7_1_to_tile_7_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(225)
	);

	pe_tile pe_tile_7_1(
		.out_wire_3_0(vertical_tile_7_1_to_tile_6_1_0),
		.out_wire_3_1(vertical_tile_7_1_to_tile_6_1_1),
		.out_wire_3_2(vertical_tile_7_1_to_tile_6_1_2),
		.out_wire_3_3(vertical_tile_7_1_to_tile_6_1_3),
		.in_wire_3_0(vertical_tile_6_1_to_tile_7_1_0),
		.in_wire_3_1(vertical_tile_6_1_to_tile_7_1_1),
		.in_wire_3_2(vertical_tile_6_1_to_tile_7_1_2),
		.in_wire_3_3(vertical_tile_6_1_to_tile_7_1_3),
		.out_wire_1_0(vertical_tile_7_1_to_tile_8_1_0),
		.out_wire_1_1(vertical_tile_7_1_to_tile_8_1_1),
		.out_wire_1_2(vertical_tile_7_1_to_tile_8_1_2),
		.out_wire_1_3(vertical_tile_7_1_to_tile_8_1_3),
		.in_wire_1_0(vertical_tile_8_1_to_tile_7_1_0),
		.in_wire_1_1(vertical_tile_8_1_to_tile_7_1_1),
		.in_wire_1_2(vertical_tile_8_1_to_tile_7_1_2),
		.in_wire_1_3(vertical_tile_8_1_to_tile_7_1_3),
		.out_wire_2_0(horizontal_tile_7_1_to_tile_7_0_0),
		.out_wire_2_1(horizontal_tile_7_1_to_tile_7_0_1),
		.out_wire_2_2(horizontal_tile_7_1_to_tile_7_0_2),
		.out_wire_2_3(horizontal_tile_7_1_to_tile_7_0_3),
		.in_wire_2_0(horizontal_tile_7_0_to_tile_7_1_0),
		.in_wire_2_1(horizontal_tile_7_0_to_tile_7_1_1),
		.in_wire_2_2(horizontal_tile_7_0_to_tile_7_1_2),
		.in_wire_2_3(horizontal_tile_7_0_to_tile_7_1_3),
		.out_wire_0_0(horizontal_tile_7_1_to_tile_7_2_0),
		.out_wire_0_1(horizontal_tile_7_1_to_tile_7_2_1),
		.out_wire_0_2(horizontal_tile_7_1_to_tile_7_2_2),
		.out_wire_0_3(horizontal_tile_7_1_to_tile_7_2_3),
		.in_wire_0_0(horizontal_tile_7_2_to_tile_7_1_0),
		.in_wire_0_1(horizontal_tile_7_2_to_tile_7_1_1),
		.in_wire_0_2(horizontal_tile_7_2_to_tile_7_1_2),
		.in_wire_0_3(horizontal_tile_7_2_to_tile_7_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(226)
	);

	pe_tile pe_tile_7_2(
		.out_wire_3_0(vertical_tile_7_2_to_tile_6_2_0),
		.out_wire_3_1(vertical_tile_7_2_to_tile_6_2_1),
		.out_wire_3_2(vertical_tile_7_2_to_tile_6_2_2),
		.out_wire_3_3(vertical_tile_7_2_to_tile_6_2_3),
		.in_wire_3_0(vertical_tile_6_2_to_tile_7_2_0),
		.in_wire_3_1(vertical_tile_6_2_to_tile_7_2_1),
		.in_wire_3_2(vertical_tile_6_2_to_tile_7_2_2),
		.in_wire_3_3(vertical_tile_6_2_to_tile_7_2_3),
		.out_wire_1_0(vertical_tile_7_2_to_tile_8_2_0),
		.out_wire_1_1(vertical_tile_7_2_to_tile_8_2_1),
		.out_wire_1_2(vertical_tile_7_2_to_tile_8_2_2),
		.out_wire_1_3(vertical_tile_7_2_to_tile_8_2_3),
		.in_wire_1_0(vertical_tile_8_2_to_tile_7_2_0),
		.in_wire_1_1(vertical_tile_8_2_to_tile_7_2_1),
		.in_wire_1_2(vertical_tile_8_2_to_tile_7_2_2),
		.in_wire_1_3(vertical_tile_8_2_to_tile_7_2_3),
		.out_wire_2_0(horizontal_tile_7_2_to_tile_7_1_0),
		.out_wire_2_1(horizontal_tile_7_2_to_tile_7_1_1),
		.out_wire_2_2(horizontal_tile_7_2_to_tile_7_1_2),
		.out_wire_2_3(horizontal_tile_7_2_to_tile_7_1_3),
		.in_wire_2_0(horizontal_tile_7_1_to_tile_7_2_0),
		.in_wire_2_1(horizontal_tile_7_1_to_tile_7_2_1),
		.in_wire_2_2(horizontal_tile_7_1_to_tile_7_2_2),
		.in_wire_2_3(horizontal_tile_7_1_to_tile_7_2_3),
		.out_wire_0_0(horizontal_tile_7_2_to_tile_7_3_0),
		.out_wire_0_1(horizontal_tile_7_2_to_tile_7_3_1),
		.out_wire_0_2(horizontal_tile_7_2_to_tile_7_3_2),
		.out_wire_0_3(horizontal_tile_7_2_to_tile_7_3_3),
		.in_wire_0_0(horizontal_tile_7_3_to_tile_7_2_0),
		.in_wire_0_1(horizontal_tile_7_3_to_tile_7_2_1),
		.in_wire_0_2(horizontal_tile_7_3_to_tile_7_2_2),
		.in_wire_0_3(horizontal_tile_7_3_to_tile_7_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(227)
	);

	pe_tile pe_tile_7_3(
		.out_wire_3_0(vertical_tile_7_3_to_tile_6_3_0),
		.out_wire_3_1(vertical_tile_7_3_to_tile_6_3_1),
		.out_wire_3_2(vertical_tile_7_3_to_tile_6_3_2),
		.out_wire_3_3(vertical_tile_7_3_to_tile_6_3_3),
		.in_wire_3_0(vertical_tile_6_3_to_tile_7_3_0),
		.in_wire_3_1(vertical_tile_6_3_to_tile_7_3_1),
		.in_wire_3_2(vertical_tile_6_3_to_tile_7_3_2),
		.in_wire_3_3(vertical_tile_6_3_to_tile_7_3_3),
		.out_wire_1_0(vertical_tile_7_3_to_tile_8_3_0),
		.out_wire_1_1(vertical_tile_7_3_to_tile_8_3_1),
		.out_wire_1_2(vertical_tile_7_3_to_tile_8_3_2),
		.out_wire_1_3(vertical_tile_7_3_to_tile_8_3_3),
		.in_wire_1_0(vertical_tile_8_3_to_tile_7_3_0),
		.in_wire_1_1(vertical_tile_8_3_to_tile_7_3_1),
		.in_wire_1_2(vertical_tile_8_3_to_tile_7_3_2),
		.in_wire_1_3(vertical_tile_8_3_to_tile_7_3_3),
		.out_wire_2_0(horizontal_tile_7_3_to_tile_7_2_0),
		.out_wire_2_1(horizontal_tile_7_3_to_tile_7_2_1),
		.out_wire_2_2(horizontal_tile_7_3_to_tile_7_2_2),
		.out_wire_2_3(horizontal_tile_7_3_to_tile_7_2_3),
		.in_wire_2_0(horizontal_tile_7_2_to_tile_7_3_0),
		.in_wire_2_1(horizontal_tile_7_2_to_tile_7_3_1),
		.in_wire_2_2(horizontal_tile_7_2_to_tile_7_3_2),
		.in_wire_2_3(horizontal_tile_7_2_to_tile_7_3_3),
		.out_wire_0_0(horizontal_tile_7_3_to_tile_7_4_0),
		.out_wire_0_1(horizontal_tile_7_3_to_tile_7_4_1),
		.out_wire_0_2(horizontal_tile_7_3_to_tile_7_4_2),
		.out_wire_0_3(horizontal_tile_7_3_to_tile_7_4_3),
		.in_wire_0_0(horizontal_tile_7_4_to_tile_7_3_0),
		.in_wire_0_1(horizontal_tile_7_4_to_tile_7_3_1),
		.in_wire_0_2(horizontal_tile_7_4_to_tile_7_3_2),
		.in_wire_0_3(horizontal_tile_7_4_to_tile_7_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(228)
	);

	pe_tile pe_tile_7_4(
		.out_wire_3_0(vertical_tile_7_4_to_tile_6_4_0),
		.out_wire_3_1(vertical_tile_7_4_to_tile_6_4_1),
		.out_wire_3_2(vertical_tile_7_4_to_tile_6_4_2),
		.out_wire_3_3(vertical_tile_7_4_to_tile_6_4_3),
		.in_wire_3_0(vertical_tile_6_4_to_tile_7_4_0),
		.in_wire_3_1(vertical_tile_6_4_to_tile_7_4_1),
		.in_wire_3_2(vertical_tile_6_4_to_tile_7_4_2),
		.in_wire_3_3(vertical_tile_6_4_to_tile_7_4_3),
		.out_wire_1_0(vertical_tile_7_4_to_tile_8_4_0),
		.out_wire_1_1(vertical_tile_7_4_to_tile_8_4_1),
		.out_wire_1_2(vertical_tile_7_4_to_tile_8_4_2),
		.out_wire_1_3(vertical_tile_7_4_to_tile_8_4_3),
		.in_wire_1_0(vertical_tile_8_4_to_tile_7_4_0),
		.in_wire_1_1(vertical_tile_8_4_to_tile_7_4_1),
		.in_wire_1_2(vertical_tile_8_4_to_tile_7_4_2),
		.in_wire_1_3(vertical_tile_8_4_to_tile_7_4_3),
		.out_wire_2_0(horizontal_tile_7_4_to_tile_7_3_0),
		.out_wire_2_1(horizontal_tile_7_4_to_tile_7_3_1),
		.out_wire_2_2(horizontal_tile_7_4_to_tile_7_3_2),
		.out_wire_2_3(horizontal_tile_7_4_to_tile_7_3_3),
		.in_wire_2_0(horizontal_tile_7_3_to_tile_7_4_0),
		.in_wire_2_1(horizontal_tile_7_3_to_tile_7_4_1),
		.in_wire_2_2(horizontal_tile_7_3_to_tile_7_4_2),
		.in_wire_2_3(horizontal_tile_7_3_to_tile_7_4_3),
		.out_wire_0_0(horizontal_tile_7_4_to_tile_7_5_0),
		.out_wire_0_1(horizontal_tile_7_4_to_tile_7_5_1),
		.out_wire_0_2(horizontal_tile_7_4_to_tile_7_5_2),
		.out_wire_0_3(horizontal_tile_7_4_to_tile_7_5_3),
		.in_wire_0_0(horizontal_tile_7_5_to_tile_7_4_0),
		.in_wire_0_1(horizontal_tile_7_5_to_tile_7_4_1),
		.in_wire_0_2(horizontal_tile_7_5_to_tile_7_4_2),
		.in_wire_0_3(horizontal_tile_7_5_to_tile_7_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(229)
	);

	pe_tile pe_tile_7_5(
		.out_wire_3_0(vertical_tile_7_5_to_tile_6_5_0),
		.out_wire_3_1(vertical_tile_7_5_to_tile_6_5_1),
		.out_wire_3_2(vertical_tile_7_5_to_tile_6_5_2),
		.out_wire_3_3(vertical_tile_7_5_to_tile_6_5_3),
		.in_wire_3_0(vertical_tile_6_5_to_tile_7_5_0),
		.in_wire_3_1(vertical_tile_6_5_to_tile_7_5_1),
		.in_wire_3_2(vertical_tile_6_5_to_tile_7_5_2),
		.in_wire_3_3(vertical_tile_6_5_to_tile_7_5_3),
		.out_wire_1_0(vertical_tile_7_5_to_tile_8_5_0),
		.out_wire_1_1(vertical_tile_7_5_to_tile_8_5_1),
		.out_wire_1_2(vertical_tile_7_5_to_tile_8_5_2),
		.out_wire_1_3(vertical_tile_7_5_to_tile_8_5_3),
		.in_wire_1_0(vertical_tile_8_5_to_tile_7_5_0),
		.in_wire_1_1(vertical_tile_8_5_to_tile_7_5_1),
		.in_wire_1_2(vertical_tile_8_5_to_tile_7_5_2),
		.in_wire_1_3(vertical_tile_8_5_to_tile_7_5_3),
		.out_wire_2_0(horizontal_tile_7_5_to_tile_7_4_0),
		.out_wire_2_1(horizontal_tile_7_5_to_tile_7_4_1),
		.out_wire_2_2(horizontal_tile_7_5_to_tile_7_4_2),
		.out_wire_2_3(horizontal_tile_7_5_to_tile_7_4_3),
		.in_wire_2_0(horizontal_tile_7_4_to_tile_7_5_0),
		.in_wire_2_1(horizontal_tile_7_4_to_tile_7_5_1),
		.in_wire_2_2(horizontal_tile_7_4_to_tile_7_5_2),
		.in_wire_2_3(horizontal_tile_7_4_to_tile_7_5_3),
		.out_wire_0_0(horizontal_tile_7_5_to_tile_7_6_0),
		.out_wire_0_1(horizontal_tile_7_5_to_tile_7_6_1),
		.out_wire_0_2(horizontal_tile_7_5_to_tile_7_6_2),
		.out_wire_0_3(horizontal_tile_7_5_to_tile_7_6_3),
		.in_wire_0_0(horizontal_tile_7_6_to_tile_7_5_0),
		.in_wire_0_1(horizontal_tile_7_6_to_tile_7_5_1),
		.in_wire_0_2(horizontal_tile_7_6_to_tile_7_5_2),
		.in_wire_0_3(horizontal_tile_7_6_to_tile_7_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(230)
	);

	pe_tile pe_tile_7_6(
		.out_wire_3_0(vertical_tile_7_6_to_tile_6_6_0),
		.out_wire_3_1(vertical_tile_7_6_to_tile_6_6_1),
		.out_wire_3_2(vertical_tile_7_6_to_tile_6_6_2),
		.out_wire_3_3(vertical_tile_7_6_to_tile_6_6_3),
		.in_wire_3_0(vertical_tile_6_6_to_tile_7_6_0),
		.in_wire_3_1(vertical_tile_6_6_to_tile_7_6_1),
		.in_wire_3_2(vertical_tile_6_6_to_tile_7_6_2),
		.in_wire_3_3(vertical_tile_6_6_to_tile_7_6_3),
		.out_wire_1_0(vertical_tile_7_6_to_tile_8_6_0),
		.out_wire_1_1(vertical_tile_7_6_to_tile_8_6_1),
		.out_wire_1_2(vertical_tile_7_6_to_tile_8_6_2),
		.out_wire_1_3(vertical_tile_7_6_to_tile_8_6_3),
		.in_wire_1_0(vertical_tile_8_6_to_tile_7_6_0),
		.in_wire_1_1(vertical_tile_8_6_to_tile_7_6_1),
		.in_wire_1_2(vertical_tile_8_6_to_tile_7_6_2),
		.in_wire_1_3(vertical_tile_8_6_to_tile_7_6_3),
		.out_wire_2_0(horizontal_tile_7_6_to_tile_7_5_0),
		.out_wire_2_1(horizontal_tile_7_6_to_tile_7_5_1),
		.out_wire_2_2(horizontal_tile_7_6_to_tile_7_5_2),
		.out_wire_2_3(horizontal_tile_7_6_to_tile_7_5_3),
		.in_wire_2_0(horizontal_tile_7_5_to_tile_7_6_0),
		.in_wire_2_1(horizontal_tile_7_5_to_tile_7_6_1),
		.in_wire_2_2(horizontal_tile_7_5_to_tile_7_6_2),
		.in_wire_2_3(horizontal_tile_7_5_to_tile_7_6_3),
		.out_wire_0_0(horizontal_tile_7_6_to_tile_7_7_0),
		.out_wire_0_1(horizontal_tile_7_6_to_tile_7_7_1),
		.out_wire_0_2(horizontal_tile_7_6_to_tile_7_7_2),
		.out_wire_0_3(horizontal_tile_7_6_to_tile_7_7_3),
		.in_wire_0_0(horizontal_tile_7_7_to_tile_7_6_0),
		.in_wire_0_1(horizontal_tile_7_7_to_tile_7_6_1),
		.in_wire_0_2(horizontal_tile_7_7_to_tile_7_6_2),
		.in_wire_0_3(horizontal_tile_7_7_to_tile_7_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(231)
	);

	pe_tile pe_tile_7_7(
		.out_wire_3_0(vertical_tile_7_7_to_tile_6_7_0),
		.out_wire_3_1(vertical_tile_7_7_to_tile_6_7_1),
		.out_wire_3_2(vertical_tile_7_7_to_tile_6_7_2),
		.out_wire_3_3(vertical_tile_7_7_to_tile_6_7_3),
		.in_wire_3_0(vertical_tile_6_7_to_tile_7_7_0),
		.in_wire_3_1(vertical_tile_6_7_to_tile_7_7_1),
		.in_wire_3_2(vertical_tile_6_7_to_tile_7_7_2),
		.in_wire_3_3(vertical_tile_6_7_to_tile_7_7_3),
		.out_wire_1_0(vertical_tile_7_7_to_tile_8_7_0),
		.out_wire_1_1(vertical_tile_7_7_to_tile_8_7_1),
		.out_wire_1_2(vertical_tile_7_7_to_tile_8_7_2),
		.out_wire_1_3(vertical_tile_7_7_to_tile_8_7_3),
		.in_wire_1_0(vertical_tile_8_7_to_tile_7_7_0),
		.in_wire_1_1(vertical_tile_8_7_to_tile_7_7_1),
		.in_wire_1_2(vertical_tile_8_7_to_tile_7_7_2),
		.in_wire_1_3(vertical_tile_8_7_to_tile_7_7_3),
		.out_wire_2_0(horizontal_tile_7_7_to_tile_7_6_0),
		.out_wire_2_1(horizontal_tile_7_7_to_tile_7_6_1),
		.out_wire_2_2(horizontal_tile_7_7_to_tile_7_6_2),
		.out_wire_2_3(horizontal_tile_7_7_to_tile_7_6_3),
		.in_wire_2_0(horizontal_tile_7_6_to_tile_7_7_0),
		.in_wire_2_1(horizontal_tile_7_6_to_tile_7_7_1),
		.in_wire_2_2(horizontal_tile_7_6_to_tile_7_7_2),
		.in_wire_2_3(horizontal_tile_7_6_to_tile_7_7_3),
		.out_wire_0_0(horizontal_tile_7_7_to_tile_7_8_0),
		.out_wire_0_1(horizontal_tile_7_7_to_tile_7_8_1),
		.out_wire_0_2(horizontal_tile_7_7_to_tile_7_8_2),
		.out_wire_0_3(horizontal_tile_7_7_to_tile_7_8_3),
		.in_wire_0_0(horizontal_tile_7_8_to_tile_7_7_0),
		.in_wire_0_1(horizontal_tile_7_8_to_tile_7_7_1),
		.in_wire_0_2(horizontal_tile_7_8_to_tile_7_7_2),
		.in_wire_0_3(horizontal_tile_7_8_to_tile_7_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(232)
	);

	pe_tile pe_tile_7_8(
		.out_wire_3_0(vertical_tile_7_8_to_tile_6_8_0),
		.out_wire_3_1(vertical_tile_7_8_to_tile_6_8_1),
		.out_wire_3_2(vertical_tile_7_8_to_tile_6_8_2),
		.out_wire_3_3(vertical_tile_7_8_to_tile_6_8_3),
		.in_wire_3_0(vertical_tile_6_8_to_tile_7_8_0),
		.in_wire_3_1(vertical_tile_6_8_to_tile_7_8_1),
		.in_wire_3_2(vertical_tile_6_8_to_tile_7_8_2),
		.in_wire_3_3(vertical_tile_6_8_to_tile_7_8_3),
		.out_wire_1_0(vertical_tile_7_8_to_tile_8_8_0),
		.out_wire_1_1(vertical_tile_7_8_to_tile_8_8_1),
		.out_wire_1_2(vertical_tile_7_8_to_tile_8_8_2),
		.out_wire_1_3(vertical_tile_7_8_to_tile_8_8_3),
		.in_wire_1_0(vertical_tile_8_8_to_tile_7_8_0),
		.in_wire_1_1(vertical_tile_8_8_to_tile_7_8_1),
		.in_wire_1_2(vertical_tile_8_8_to_tile_7_8_2),
		.in_wire_1_3(vertical_tile_8_8_to_tile_7_8_3),
		.out_wire_2_0(horizontal_tile_7_8_to_tile_7_7_0),
		.out_wire_2_1(horizontal_tile_7_8_to_tile_7_7_1),
		.out_wire_2_2(horizontal_tile_7_8_to_tile_7_7_2),
		.out_wire_2_3(horizontal_tile_7_8_to_tile_7_7_3),
		.in_wire_2_0(horizontal_tile_7_7_to_tile_7_8_0),
		.in_wire_2_1(horizontal_tile_7_7_to_tile_7_8_1),
		.in_wire_2_2(horizontal_tile_7_7_to_tile_7_8_2),
		.in_wire_2_3(horizontal_tile_7_7_to_tile_7_8_3),
		.out_wire_0_0(horizontal_tile_7_8_to_tile_7_9_0),
		.out_wire_0_1(horizontal_tile_7_8_to_tile_7_9_1),
		.out_wire_0_2(horizontal_tile_7_8_to_tile_7_9_2),
		.out_wire_0_3(horizontal_tile_7_8_to_tile_7_9_3),
		.in_wire_0_0(horizontal_tile_7_9_to_tile_7_8_0),
		.in_wire_0_1(horizontal_tile_7_9_to_tile_7_8_1),
		.in_wire_0_2(horizontal_tile_7_9_to_tile_7_8_2),
		.in_wire_0_3(horizontal_tile_7_9_to_tile_7_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(233)
	);

	pe_tile pe_tile_7_9(
		.out_wire_3_0(vertical_tile_7_9_to_tile_6_9_0),
		.out_wire_3_1(vertical_tile_7_9_to_tile_6_9_1),
		.out_wire_3_2(vertical_tile_7_9_to_tile_6_9_2),
		.out_wire_3_3(vertical_tile_7_9_to_tile_6_9_3),
		.in_wire_3_0(vertical_tile_6_9_to_tile_7_9_0),
		.in_wire_3_1(vertical_tile_6_9_to_tile_7_9_1),
		.in_wire_3_2(vertical_tile_6_9_to_tile_7_9_2),
		.in_wire_3_3(vertical_tile_6_9_to_tile_7_9_3),
		.out_wire_1_0(vertical_tile_7_9_to_tile_8_9_0),
		.out_wire_1_1(vertical_tile_7_9_to_tile_8_9_1),
		.out_wire_1_2(vertical_tile_7_9_to_tile_8_9_2),
		.out_wire_1_3(vertical_tile_7_9_to_tile_8_9_3),
		.in_wire_1_0(vertical_tile_8_9_to_tile_7_9_0),
		.in_wire_1_1(vertical_tile_8_9_to_tile_7_9_1),
		.in_wire_1_2(vertical_tile_8_9_to_tile_7_9_2),
		.in_wire_1_3(vertical_tile_8_9_to_tile_7_9_3),
		.out_wire_2_0(horizontal_tile_7_9_to_tile_7_8_0),
		.out_wire_2_1(horizontal_tile_7_9_to_tile_7_8_1),
		.out_wire_2_2(horizontal_tile_7_9_to_tile_7_8_2),
		.out_wire_2_3(horizontal_tile_7_9_to_tile_7_8_3),
		.in_wire_2_0(horizontal_tile_7_8_to_tile_7_9_0),
		.in_wire_2_1(horizontal_tile_7_8_to_tile_7_9_1),
		.in_wire_2_2(horizontal_tile_7_8_to_tile_7_9_2),
		.in_wire_2_3(horizontal_tile_7_8_to_tile_7_9_3),
		.out_wire_0_0(horizontal_tile_7_9_to_tile_7_10_0),
		.out_wire_0_1(horizontal_tile_7_9_to_tile_7_10_1),
		.out_wire_0_2(horizontal_tile_7_9_to_tile_7_10_2),
		.out_wire_0_3(horizontal_tile_7_9_to_tile_7_10_3),
		.in_wire_0_0(horizontal_tile_7_10_to_tile_7_9_0),
		.in_wire_0_1(horizontal_tile_7_10_to_tile_7_9_1),
		.in_wire_0_2(horizontal_tile_7_10_to_tile_7_9_2),
		.in_wire_0_3(horizontal_tile_7_10_to_tile_7_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(234)
	);

	pe_tile pe_tile_7_10(
		.out_wire_3_0(vertical_tile_7_10_to_tile_6_10_0),
		.out_wire_3_1(vertical_tile_7_10_to_tile_6_10_1),
		.out_wire_3_2(vertical_tile_7_10_to_tile_6_10_2),
		.out_wire_3_3(vertical_tile_7_10_to_tile_6_10_3),
		.in_wire_3_0(vertical_tile_6_10_to_tile_7_10_0),
		.in_wire_3_1(vertical_tile_6_10_to_tile_7_10_1),
		.in_wire_3_2(vertical_tile_6_10_to_tile_7_10_2),
		.in_wire_3_3(vertical_tile_6_10_to_tile_7_10_3),
		.out_wire_1_0(vertical_tile_7_10_to_tile_8_10_0),
		.out_wire_1_1(vertical_tile_7_10_to_tile_8_10_1),
		.out_wire_1_2(vertical_tile_7_10_to_tile_8_10_2),
		.out_wire_1_3(vertical_tile_7_10_to_tile_8_10_3),
		.in_wire_1_0(vertical_tile_8_10_to_tile_7_10_0),
		.in_wire_1_1(vertical_tile_8_10_to_tile_7_10_1),
		.in_wire_1_2(vertical_tile_8_10_to_tile_7_10_2),
		.in_wire_1_3(vertical_tile_8_10_to_tile_7_10_3),
		.out_wire_2_0(horizontal_tile_7_10_to_tile_7_9_0),
		.out_wire_2_1(horizontal_tile_7_10_to_tile_7_9_1),
		.out_wire_2_2(horizontal_tile_7_10_to_tile_7_9_2),
		.out_wire_2_3(horizontal_tile_7_10_to_tile_7_9_3),
		.in_wire_2_0(horizontal_tile_7_9_to_tile_7_10_0),
		.in_wire_2_1(horizontal_tile_7_9_to_tile_7_10_1),
		.in_wire_2_2(horizontal_tile_7_9_to_tile_7_10_2),
		.in_wire_2_3(horizontal_tile_7_9_to_tile_7_10_3),
		.out_wire_0_0(horizontal_tile_7_10_to_tile_7_11_0),
		.out_wire_0_1(horizontal_tile_7_10_to_tile_7_11_1),
		.out_wire_0_2(horizontal_tile_7_10_to_tile_7_11_2),
		.out_wire_0_3(horizontal_tile_7_10_to_tile_7_11_3),
		.in_wire_0_0(horizontal_tile_7_11_to_tile_7_10_0),
		.in_wire_0_1(horizontal_tile_7_11_to_tile_7_10_1),
		.in_wire_0_2(horizontal_tile_7_11_to_tile_7_10_2),
		.in_wire_0_3(horizontal_tile_7_11_to_tile_7_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(235)
	);

	pe_tile pe_tile_7_11(
		.out_wire_3_0(vertical_tile_7_11_to_tile_6_11_0),
		.out_wire_3_1(vertical_tile_7_11_to_tile_6_11_1),
		.out_wire_3_2(vertical_tile_7_11_to_tile_6_11_2),
		.out_wire_3_3(vertical_tile_7_11_to_tile_6_11_3),
		.in_wire_3_0(vertical_tile_6_11_to_tile_7_11_0),
		.in_wire_3_1(vertical_tile_6_11_to_tile_7_11_1),
		.in_wire_3_2(vertical_tile_6_11_to_tile_7_11_2),
		.in_wire_3_3(vertical_tile_6_11_to_tile_7_11_3),
		.out_wire_1_0(vertical_tile_7_11_to_tile_8_11_0),
		.out_wire_1_1(vertical_tile_7_11_to_tile_8_11_1),
		.out_wire_1_2(vertical_tile_7_11_to_tile_8_11_2),
		.out_wire_1_3(vertical_tile_7_11_to_tile_8_11_3),
		.in_wire_1_0(vertical_tile_8_11_to_tile_7_11_0),
		.in_wire_1_1(vertical_tile_8_11_to_tile_7_11_1),
		.in_wire_1_2(vertical_tile_8_11_to_tile_7_11_2),
		.in_wire_1_3(vertical_tile_8_11_to_tile_7_11_3),
		.out_wire_2_0(horizontal_tile_7_11_to_tile_7_10_0),
		.out_wire_2_1(horizontal_tile_7_11_to_tile_7_10_1),
		.out_wire_2_2(horizontal_tile_7_11_to_tile_7_10_2),
		.out_wire_2_3(horizontal_tile_7_11_to_tile_7_10_3),
		.in_wire_2_0(horizontal_tile_7_10_to_tile_7_11_0),
		.in_wire_2_1(horizontal_tile_7_10_to_tile_7_11_1),
		.in_wire_2_2(horizontal_tile_7_10_to_tile_7_11_2),
		.in_wire_2_3(horizontal_tile_7_10_to_tile_7_11_3),
		.out_wire_0_0(horizontal_tile_7_11_to_tile_7_12_0),
		.out_wire_0_1(horizontal_tile_7_11_to_tile_7_12_1),
		.out_wire_0_2(horizontal_tile_7_11_to_tile_7_12_2),
		.out_wire_0_3(horizontal_tile_7_11_to_tile_7_12_3),
		.in_wire_0_0(horizontal_tile_7_12_to_tile_7_11_0),
		.in_wire_0_1(horizontal_tile_7_12_to_tile_7_11_1),
		.in_wire_0_2(horizontal_tile_7_12_to_tile_7_11_2),
		.in_wire_0_3(horizontal_tile_7_12_to_tile_7_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(236)
	);

	pe_tile pe_tile_7_12(
		.out_wire_3_0(vertical_tile_7_12_to_tile_6_12_0),
		.out_wire_3_1(vertical_tile_7_12_to_tile_6_12_1),
		.out_wire_3_2(vertical_tile_7_12_to_tile_6_12_2),
		.out_wire_3_3(vertical_tile_7_12_to_tile_6_12_3),
		.in_wire_3_0(vertical_tile_6_12_to_tile_7_12_0),
		.in_wire_3_1(vertical_tile_6_12_to_tile_7_12_1),
		.in_wire_3_2(vertical_tile_6_12_to_tile_7_12_2),
		.in_wire_3_3(vertical_tile_6_12_to_tile_7_12_3),
		.out_wire_1_0(vertical_tile_7_12_to_tile_8_12_0),
		.out_wire_1_1(vertical_tile_7_12_to_tile_8_12_1),
		.out_wire_1_2(vertical_tile_7_12_to_tile_8_12_2),
		.out_wire_1_3(vertical_tile_7_12_to_tile_8_12_3),
		.in_wire_1_0(vertical_tile_8_12_to_tile_7_12_0),
		.in_wire_1_1(vertical_tile_8_12_to_tile_7_12_1),
		.in_wire_1_2(vertical_tile_8_12_to_tile_7_12_2),
		.in_wire_1_3(vertical_tile_8_12_to_tile_7_12_3),
		.out_wire_2_0(horizontal_tile_7_12_to_tile_7_11_0),
		.out_wire_2_1(horizontal_tile_7_12_to_tile_7_11_1),
		.out_wire_2_2(horizontal_tile_7_12_to_tile_7_11_2),
		.out_wire_2_3(horizontal_tile_7_12_to_tile_7_11_3),
		.in_wire_2_0(horizontal_tile_7_11_to_tile_7_12_0),
		.in_wire_2_1(horizontal_tile_7_11_to_tile_7_12_1),
		.in_wire_2_2(horizontal_tile_7_11_to_tile_7_12_2),
		.in_wire_2_3(horizontal_tile_7_11_to_tile_7_12_3),
		.out_wire_0_0(horizontal_tile_7_12_to_tile_7_13_0),
		.out_wire_0_1(horizontal_tile_7_12_to_tile_7_13_1),
		.out_wire_0_2(horizontal_tile_7_12_to_tile_7_13_2),
		.out_wire_0_3(horizontal_tile_7_12_to_tile_7_13_3),
		.in_wire_0_0(horizontal_tile_7_13_to_tile_7_12_0),
		.in_wire_0_1(horizontal_tile_7_13_to_tile_7_12_1),
		.in_wire_0_2(horizontal_tile_7_13_to_tile_7_12_2),
		.in_wire_0_3(horizontal_tile_7_13_to_tile_7_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(237)
	);

	pe_tile pe_tile_7_13(
		.out_wire_3_0(vertical_tile_7_13_to_tile_6_13_0),
		.out_wire_3_1(vertical_tile_7_13_to_tile_6_13_1),
		.out_wire_3_2(vertical_tile_7_13_to_tile_6_13_2),
		.out_wire_3_3(vertical_tile_7_13_to_tile_6_13_3),
		.in_wire_3_0(vertical_tile_6_13_to_tile_7_13_0),
		.in_wire_3_1(vertical_tile_6_13_to_tile_7_13_1),
		.in_wire_3_2(vertical_tile_6_13_to_tile_7_13_2),
		.in_wire_3_3(vertical_tile_6_13_to_tile_7_13_3),
		.out_wire_1_0(vertical_tile_7_13_to_tile_8_13_0),
		.out_wire_1_1(vertical_tile_7_13_to_tile_8_13_1),
		.out_wire_1_2(vertical_tile_7_13_to_tile_8_13_2),
		.out_wire_1_3(vertical_tile_7_13_to_tile_8_13_3),
		.in_wire_1_0(vertical_tile_8_13_to_tile_7_13_0),
		.in_wire_1_1(vertical_tile_8_13_to_tile_7_13_1),
		.in_wire_1_2(vertical_tile_8_13_to_tile_7_13_2),
		.in_wire_1_3(vertical_tile_8_13_to_tile_7_13_3),
		.out_wire_2_0(horizontal_tile_7_13_to_tile_7_12_0),
		.out_wire_2_1(horizontal_tile_7_13_to_tile_7_12_1),
		.out_wire_2_2(horizontal_tile_7_13_to_tile_7_12_2),
		.out_wire_2_3(horizontal_tile_7_13_to_tile_7_12_3),
		.in_wire_2_0(horizontal_tile_7_12_to_tile_7_13_0),
		.in_wire_2_1(horizontal_tile_7_12_to_tile_7_13_1),
		.in_wire_2_2(horizontal_tile_7_12_to_tile_7_13_2),
		.in_wire_2_3(horizontal_tile_7_12_to_tile_7_13_3),
		.out_wire_0_0(horizontal_tile_7_13_to_tile_7_14_0),
		.out_wire_0_1(horizontal_tile_7_13_to_tile_7_14_1),
		.out_wire_0_2(horizontal_tile_7_13_to_tile_7_14_2),
		.out_wire_0_3(horizontal_tile_7_13_to_tile_7_14_3),
		.in_wire_0_0(horizontal_tile_7_14_to_tile_7_13_0),
		.in_wire_0_1(horizontal_tile_7_14_to_tile_7_13_1),
		.in_wire_0_2(horizontal_tile_7_14_to_tile_7_13_2),
		.in_wire_0_3(horizontal_tile_7_14_to_tile_7_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(238)
	);

	pe_tile pe_tile_7_14(
		.out_wire_3_0(vertical_tile_7_14_to_tile_6_14_0),
		.out_wire_3_1(vertical_tile_7_14_to_tile_6_14_1),
		.out_wire_3_2(vertical_tile_7_14_to_tile_6_14_2),
		.out_wire_3_3(vertical_tile_7_14_to_tile_6_14_3),
		.in_wire_3_0(vertical_tile_6_14_to_tile_7_14_0),
		.in_wire_3_1(vertical_tile_6_14_to_tile_7_14_1),
		.in_wire_3_2(vertical_tile_6_14_to_tile_7_14_2),
		.in_wire_3_3(vertical_tile_6_14_to_tile_7_14_3),
		.out_wire_1_0(vertical_tile_7_14_to_tile_8_14_0),
		.out_wire_1_1(vertical_tile_7_14_to_tile_8_14_1),
		.out_wire_1_2(vertical_tile_7_14_to_tile_8_14_2),
		.out_wire_1_3(vertical_tile_7_14_to_tile_8_14_3),
		.in_wire_1_0(vertical_tile_8_14_to_tile_7_14_0),
		.in_wire_1_1(vertical_tile_8_14_to_tile_7_14_1),
		.in_wire_1_2(vertical_tile_8_14_to_tile_7_14_2),
		.in_wire_1_3(vertical_tile_8_14_to_tile_7_14_3),
		.out_wire_2_0(horizontal_tile_7_14_to_tile_7_13_0),
		.out_wire_2_1(horizontal_tile_7_14_to_tile_7_13_1),
		.out_wire_2_2(horizontal_tile_7_14_to_tile_7_13_2),
		.out_wire_2_3(horizontal_tile_7_14_to_tile_7_13_3),
		.in_wire_2_0(horizontal_tile_7_13_to_tile_7_14_0),
		.in_wire_2_1(horizontal_tile_7_13_to_tile_7_14_1),
		.in_wire_2_2(horizontal_tile_7_13_to_tile_7_14_2),
		.in_wire_2_3(horizontal_tile_7_13_to_tile_7_14_3),
		.out_wire_0_0(horizontal_tile_7_14_to_tile_7_15_0),
		.out_wire_0_1(horizontal_tile_7_14_to_tile_7_15_1),
		.out_wire_0_2(horizontal_tile_7_14_to_tile_7_15_2),
		.out_wire_0_3(horizontal_tile_7_14_to_tile_7_15_3),
		.in_wire_0_0(horizontal_tile_7_15_to_tile_7_14_0),
		.in_wire_0_1(horizontal_tile_7_15_to_tile_7_14_1),
		.in_wire_0_2(horizontal_tile_7_15_to_tile_7_14_2),
		.in_wire_0_3(horizontal_tile_7_15_to_tile_7_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(239)
	);

	pe_tile pe_tile_7_15(
		.out_wire_3_0(vertical_tile_7_15_to_tile_6_15_0),
		.out_wire_3_1(vertical_tile_7_15_to_tile_6_15_1),
		.out_wire_3_2(vertical_tile_7_15_to_tile_6_15_2),
		.out_wire_3_3(vertical_tile_7_15_to_tile_6_15_3),
		.in_wire_3_0(vertical_tile_6_15_to_tile_7_15_0),
		.in_wire_3_1(vertical_tile_6_15_to_tile_7_15_1),
		.in_wire_3_2(vertical_tile_6_15_to_tile_7_15_2),
		.in_wire_3_3(vertical_tile_6_15_to_tile_7_15_3),
		.out_wire_1_0(vertical_tile_7_15_to_tile_8_15_0),
		.out_wire_1_1(vertical_tile_7_15_to_tile_8_15_1),
		.out_wire_1_2(vertical_tile_7_15_to_tile_8_15_2),
		.out_wire_1_3(vertical_tile_7_15_to_tile_8_15_3),
		.in_wire_1_0(vertical_tile_8_15_to_tile_7_15_0),
		.in_wire_1_1(vertical_tile_8_15_to_tile_7_15_1),
		.in_wire_1_2(vertical_tile_8_15_to_tile_7_15_2),
		.in_wire_1_3(vertical_tile_8_15_to_tile_7_15_3),
		.out_wire_2_0(horizontal_tile_7_15_to_tile_7_14_0),
		.out_wire_2_1(horizontal_tile_7_15_to_tile_7_14_1),
		.out_wire_2_2(horizontal_tile_7_15_to_tile_7_14_2),
		.out_wire_2_3(horizontal_tile_7_15_to_tile_7_14_3),
		.in_wire_2_0(horizontal_tile_7_14_to_tile_7_15_0),
		.in_wire_2_1(horizontal_tile_7_14_to_tile_7_15_1),
		.in_wire_2_2(horizontal_tile_7_14_to_tile_7_15_2),
		.in_wire_2_3(horizontal_tile_7_14_to_tile_7_15_3),
		.out_wire_0_0(horizontal_tile_7_15_to_tile_7_16_0),
		.out_wire_0_1(horizontal_tile_7_15_to_tile_7_16_1),
		.out_wire_0_2(horizontal_tile_7_15_to_tile_7_16_2),
		.out_wire_0_3(horizontal_tile_7_15_to_tile_7_16_3),
		.in_wire_0_0(horizontal_tile_7_16_to_tile_7_15_0),
		.in_wire_0_1(horizontal_tile_7_16_to_tile_7_15_1),
		.in_wire_0_2(horizontal_tile_7_16_to_tile_7_15_2),
		.in_wire_0_3(horizontal_tile_7_16_to_tile_7_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(240)
	);

	pe_tile pe_tile_7_16(
		.out_wire_3_0(vertical_tile_7_16_to_tile_6_16_0),
		.out_wire_3_1(vertical_tile_7_16_to_tile_6_16_1),
		.out_wire_3_2(vertical_tile_7_16_to_tile_6_16_2),
		.out_wire_3_3(vertical_tile_7_16_to_tile_6_16_3),
		.in_wire_3_0(vertical_tile_6_16_to_tile_7_16_0),
		.in_wire_3_1(vertical_tile_6_16_to_tile_7_16_1),
		.in_wire_3_2(vertical_tile_6_16_to_tile_7_16_2),
		.in_wire_3_3(vertical_tile_6_16_to_tile_7_16_3),
		.out_wire_1_0(vertical_tile_7_16_to_tile_8_16_0),
		.out_wire_1_1(vertical_tile_7_16_to_tile_8_16_1),
		.out_wire_1_2(vertical_tile_7_16_to_tile_8_16_2),
		.out_wire_1_3(vertical_tile_7_16_to_tile_8_16_3),
		.in_wire_1_0(vertical_tile_8_16_to_tile_7_16_0),
		.in_wire_1_1(vertical_tile_8_16_to_tile_7_16_1),
		.in_wire_1_2(vertical_tile_8_16_to_tile_7_16_2),
		.in_wire_1_3(vertical_tile_8_16_to_tile_7_16_3),
		.out_wire_2_0(horizontal_tile_7_16_to_tile_7_15_0),
		.out_wire_2_1(horizontal_tile_7_16_to_tile_7_15_1),
		.out_wire_2_2(horizontal_tile_7_16_to_tile_7_15_2),
		.out_wire_2_3(horizontal_tile_7_16_to_tile_7_15_3),
		.in_wire_2_0(horizontal_tile_7_15_to_tile_7_16_0),
		.in_wire_2_1(horizontal_tile_7_15_to_tile_7_16_1),
		.in_wire_2_2(horizontal_tile_7_15_to_tile_7_16_2),
		.in_wire_2_3(horizontal_tile_7_15_to_tile_7_16_3),
		.out_wire_0_0(horizontal_tile_7_16_to_tile_7_17_0),
		.out_wire_0_1(horizontal_tile_7_16_to_tile_7_17_1),
		.out_wire_0_2(horizontal_tile_7_16_to_tile_7_17_2),
		.out_wire_0_3(horizontal_tile_7_16_to_tile_7_17_3),
		.in_wire_0_0(horizontal_tile_7_17_to_tile_7_16_0),
		.in_wire_0_1(horizontal_tile_7_17_to_tile_7_16_1),
		.in_wire_0_2(horizontal_tile_7_17_to_tile_7_16_2),
		.in_wire_0_3(horizontal_tile_7_17_to_tile_7_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(241)
	);

	pe_tile pe_tile_7_17(
		.out_wire_3_0(vertical_tile_7_17_to_tile_6_17_0),
		.out_wire_3_1(vertical_tile_7_17_to_tile_6_17_1),
		.out_wire_3_2(vertical_tile_7_17_to_tile_6_17_2),
		.out_wire_3_3(vertical_tile_7_17_to_tile_6_17_3),
		.in_wire_3_0(vertical_tile_6_17_to_tile_7_17_0),
		.in_wire_3_1(vertical_tile_6_17_to_tile_7_17_1),
		.in_wire_3_2(vertical_tile_6_17_to_tile_7_17_2),
		.in_wire_3_3(vertical_tile_6_17_to_tile_7_17_3),
		.out_wire_1_0(vertical_tile_7_17_to_tile_8_17_0),
		.out_wire_1_1(vertical_tile_7_17_to_tile_8_17_1),
		.out_wire_1_2(vertical_tile_7_17_to_tile_8_17_2),
		.out_wire_1_3(vertical_tile_7_17_to_tile_8_17_3),
		.in_wire_1_0(vertical_tile_8_17_to_tile_7_17_0),
		.in_wire_1_1(vertical_tile_8_17_to_tile_7_17_1),
		.in_wire_1_2(vertical_tile_8_17_to_tile_7_17_2),
		.in_wire_1_3(vertical_tile_8_17_to_tile_7_17_3),
		.out_wire_2_0(horizontal_tile_7_17_to_tile_7_16_0),
		.out_wire_2_1(horizontal_tile_7_17_to_tile_7_16_1),
		.out_wire_2_2(horizontal_tile_7_17_to_tile_7_16_2),
		.out_wire_2_3(horizontal_tile_7_17_to_tile_7_16_3),
		.in_wire_2_0(horizontal_tile_7_16_to_tile_7_17_0),
		.in_wire_2_1(horizontal_tile_7_16_to_tile_7_17_1),
		.in_wire_2_2(horizontal_tile_7_16_to_tile_7_17_2),
		.in_wire_2_3(horizontal_tile_7_16_to_tile_7_17_3),
		.out_wire_0_0(horizontal_tile_7_17_to_tile_7_18_0),
		.out_wire_0_1(horizontal_tile_7_17_to_tile_7_18_1),
		.out_wire_0_2(horizontal_tile_7_17_to_tile_7_18_2),
		.out_wire_0_3(horizontal_tile_7_17_to_tile_7_18_3),
		.in_wire_0_0(horizontal_tile_7_18_to_tile_7_17_0),
		.in_wire_0_1(horizontal_tile_7_18_to_tile_7_17_1),
		.in_wire_0_2(horizontal_tile_7_18_to_tile_7_17_2),
		.in_wire_0_3(horizontal_tile_7_18_to_tile_7_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(242)
	);

	pe_tile pe_tile_7_18(
		.out_wire_3_0(vertical_tile_7_18_to_tile_6_18_0),
		.out_wire_3_1(vertical_tile_7_18_to_tile_6_18_1),
		.out_wire_3_2(vertical_tile_7_18_to_tile_6_18_2),
		.out_wire_3_3(vertical_tile_7_18_to_tile_6_18_3),
		.in_wire_3_0(vertical_tile_6_18_to_tile_7_18_0),
		.in_wire_3_1(vertical_tile_6_18_to_tile_7_18_1),
		.in_wire_3_2(vertical_tile_6_18_to_tile_7_18_2),
		.in_wire_3_3(vertical_tile_6_18_to_tile_7_18_3),
		.out_wire_1_0(vertical_tile_7_18_to_tile_8_18_0),
		.out_wire_1_1(vertical_tile_7_18_to_tile_8_18_1),
		.out_wire_1_2(vertical_tile_7_18_to_tile_8_18_2),
		.out_wire_1_3(vertical_tile_7_18_to_tile_8_18_3),
		.in_wire_1_0(vertical_tile_8_18_to_tile_7_18_0),
		.in_wire_1_1(vertical_tile_8_18_to_tile_7_18_1),
		.in_wire_1_2(vertical_tile_8_18_to_tile_7_18_2),
		.in_wire_1_3(vertical_tile_8_18_to_tile_7_18_3),
		.out_wire_2_0(horizontal_tile_7_18_to_tile_7_17_0),
		.out_wire_2_1(horizontal_tile_7_18_to_tile_7_17_1),
		.out_wire_2_2(horizontal_tile_7_18_to_tile_7_17_2),
		.out_wire_2_3(horizontal_tile_7_18_to_tile_7_17_3),
		.in_wire_2_0(horizontal_tile_7_17_to_tile_7_18_0),
		.in_wire_2_1(horizontal_tile_7_17_to_tile_7_18_1),
		.in_wire_2_2(horizontal_tile_7_17_to_tile_7_18_2),
		.in_wire_2_3(horizontal_tile_7_17_to_tile_7_18_3),
		.out_wire_0_0(horizontal_tile_7_18_to_tile_7_19_0),
		.out_wire_0_1(horizontal_tile_7_18_to_tile_7_19_1),
		.out_wire_0_2(horizontal_tile_7_18_to_tile_7_19_2),
		.out_wire_0_3(horizontal_tile_7_18_to_tile_7_19_3),
		.in_wire_0_0(horizontal_tile_7_19_to_tile_7_18_0),
		.in_wire_0_1(horizontal_tile_7_19_to_tile_7_18_1),
		.in_wire_0_2(horizontal_tile_7_19_to_tile_7_18_2),
		.in_wire_0_3(horizontal_tile_7_19_to_tile_7_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(243)
	);

	pe_tile pe_tile_7_19(
		.out_wire_3_0(vertical_tile_7_19_to_tile_6_19_0),
		.out_wire_3_1(vertical_tile_7_19_to_tile_6_19_1),
		.out_wire_3_2(vertical_tile_7_19_to_tile_6_19_2),
		.out_wire_3_3(vertical_tile_7_19_to_tile_6_19_3),
		.in_wire_3_0(vertical_tile_6_19_to_tile_7_19_0),
		.in_wire_3_1(vertical_tile_6_19_to_tile_7_19_1),
		.in_wire_3_2(vertical_tile_6_19_to_tile_7_19_2),
		.in_wire_3_3(vertical_tile_6_19_to_tile_7_19_3),
		.out_wire_1_0(vertical_tile_7_19_to_tile_8_19_0),
		.out_wire_1_1(vertical_tile_7_19_to_tile_8_19_1),
		.out_wire_1_2(vertical_tile_7_19_to_tile_8_19_2),
		.out_wire_1_3(vertical_tile_7_19_to_tile_8_19_3),
		.in_wire_1_0(vertical_tile_8_19_to_tile_7_19_0),
		.in_wire_1_1(vertical_tile_8_19_to_tile_7_19_1),
		.in_wire_1_2(vertical_tile_8_19_to_tile_7_19_2),
		.in_wire_1_3(vertical_tile_8_19_to_tile_7_19_3),
		.out_wire_2_0(horizontal_tile_7_19_to_tile_7_18_0),
		.out_wire_2_1(horizontal_tile_7_19_to_tile_7_18_1),
		.out_wire_2_2(horizontal_tile_7_19_to_tile_7_18_2),
		.out_wire_2_3(horizontal_tile_7_19_to_tile_7_18_3),
		.in_wire_2_0(horizontal_tile_7_18_to_tile_7_19_0),
		.in_wire_2_1(horizontal_tile_7_18_to_tile_7_19_1),
		.in_wire_2_2(horizontal_tile_7_18_to_tile_7_19_2),
		.in_wire_2_3(horizontal_tile_7_18_to_tile_7_19_3),
		.out_wire_0_0(horizontal_tile_7_19_to_tile_7_20_0),
		.out_wire_0_1(horizontal_tile_7_19_to_tile_7_20_1),
		.out_wire_0_2(horizontal_tile_7_19_to_tile_7_20_2),
		.out_wire_0_3(horizontal_tile_7_19_to_tile_7_20_3),
		.in_wire_0_0(horizontal_tile_7_20_to_tile_7_19_0),
		.in_wire_0_1(horizontal_tile_7_20_to_tile_7_19_1),
		.in_wire_0_2(horizontal_tile_7_20_to_tile_7_19_2),
		.in_wire_0_3(horizontal_tile_7_20_to_tile_7_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(244)
	);

	pe_tile pe_tile_7_20(
		.out_wire_3_0(vertical_tile_7_20_to_tile_6_20_0),
		.out_wire_3_1(vertical_tile_7_20_to_tile_6_20_1),
		.out_wire_3_2(vertical_tile_7_20_to_tile_6_20_2),
		.out_wire_3_3(vertical_tile_7_20_to_tile_6_20_3),
		.in_wire_3_0(vertical_tile_6_20_to_tile_7_20_0),
		.in_wire_3_1(vertical_tile_6_20_to_tile_7_20_1),
		.in_wire_3_2(vertical_tile_6_20_to_tile_7_20_2),
		.in_wire_3_3(vertical_tile_6_20_to_tile_7_20_3),
		.out_wire_1_0(vertical_tile_7_20_to_tile_8_20_0),
		.out_wire_1_1(vertical_tile_7_20_to_tile_8_20_1),
		.out_wire_1_2(vertical_tile_7_20_to_tile_8_20_2),
		.out_wire_1_3(vertical_tile_7_20_to_tile_8_20_3),
		.in_wire_1_0(vertical_tile_8_20_to_tile_7_20_0),
		.in_wire_1_1(vertical_tile_8_20_to_tile_7_20_1),
		.in_wire_1_2(vertical_tile_8_20_to_tile_7_20_2),
		.in_wire_1_3(vertical_tile_8_20_to_tile_7_20_3),
		.out_wire_2_0(horizontal_tile_7_20_to_tile_7_19_0),
		.out_wire_2_1(horizontal_tile_7_20_to_tile_7_19_1),
		.out_wire_2_2(horizontal_tile_7_20_to_tile_7_19_2),
		.out_wire_2_3(horizontal_tile_7_20_to_tile_7_19_3),
		.in_wire_2_0(horizontal_tile_7_19_to_tile_7_20_0),
		.in_wire_2_1(horizontal_tile_7_19_to_tile_7_20_1),
		.in_wire_2_2(horizontal_tile_7_19_to_tile_7_20_2),
		.in_wire_2_3(horizontal_tile_7_19_to_tile_7_20_3),
		.out_wire_0_0(horizontal_tile_7_20_to_tile_7_21_0),
		.out_wire_0_1(horizontal_tile_7_20_to_tile_7_21_1),
		.out_wire_0_2(horizontal_tile_7_20_to_tile_7_21_2),
		.out_wire_0_3(horizontal_tile_7_20_to_tile_7_21_3),
		.in_wire_0_0(horizontal_tile_7_21_to_tile_7_20_0),
		.in_wire_0_1(horizontal_tile_7_21_to_tile_7_20_1),
		.in_wire_0_2(horizontal_tile_7_21_to_tile_7_20_2),
		.in_wire_0_3(horizontal_tile_7_21_to_tile_7_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(245)
	);

	pe_tile pe_tile_7_21(
		.out_wire_3_0(vertical_tile_7_21_to_tile_6_21_0),
		.out_wire_3_1(vertical_tile_7_21_to_tile_6_21_1),
		.out_wire_3_2(vertical_tile_7_21_to_tile_6_21_2),
		.out_wire_3_3(vertical_tile_7_21_to_tile_6_21_3),
		.in_wire_3_0(vertical_tile_6_21_to_tile_7_21_0),
		.in_wire_3_1(vertical_tile_6_21_to_tile_7_21_1),
		.in_wire_3_2(vertical_tile_6_21_to_tile_7_21_2),
		.in_wire_3_3(vertical_tile_6_21_to_tile_7_21_3),
		.out_wire_1_0(vertical_tile_7_21_to_tile_8_21_0),
		.out_wire_1_1(vertical_tile_7_21_to_tile_8_21_1),
		.out_wire_1_2(vertical_tile_7_21_to_tile_8_21_2),
		.out_wire_1_3(vertical_tile_7_21_to_tile_8_21_3),
		.in_wire_1_0(vertical_tile_8_21_to_tile_7_21_0),
		.in_wire_1_1(vertical_tile_8_21_to_tile_7_21_1),
		.in_wire_1_2(vertical_tile_8_21_to_tile_7_21_2),
		.in_wire_1_3(vertical_tile_8_21_to_tile_7_21_3),
		.out_wire_2_0(horizontal_tile_7_21_to_tile_7_20_0),
		.out_wire_2_1(horizontal_tile_7_21_to_tile_7_20_1),
		.out_wire_2_2(horizontal_tile_7_21_to_tile_7_20_2),
		.out_wire_2_3(horizontal_tile_7_21_to_tile_7_20_3),
		.in_wire_2_0(horizontal_tile_7_20_to_tile_7_21_0),
		.in_wire_2_1(horizontal_tile_7_20_to_tile_7_21_1),
		.in_wire_2_2(horizontal_tile_7_20_to_tile_7_21_2),
		.in_wire_2_3(horizontal_tile_7_20_to_tile_7_21_3),
		.out_wire_0_0(horizontal_tile_7_21_to_tile_7_22_0),
		.out_wire_0_1(horizontal_tile_7_21_to_tile_7_22_1),
		.out_wire_0_2(horizontal_tile_7_21_to_tile_7_22_2),
		.out_wire_0_3(horizontal_tile_7_21_to_tile_7_22_3),
		.in_wire_0_0(horizontal_tile_7_22_to_tile_7_21_0),
		.in_wire_0_1(horizontal_tile_7_22_to_tile_7_21_1),
		.in_wire_0_2(horizontal_tile_7_22_to_tile_7_21_2),
		.in_wire_0_3(horizontal_tile_7_22_to_tile_7_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(246)
	);

	pe_tile pe_tile_7_22(
		.out_wire_3_0(vertical_tile_7_22_to_tile_6_22_0),
		.out_wire_3_1(vertical_tile_7_22_to_tile_6_22_1),
		.out_wire_3_2(vertical_tile_7_22_to_tile_6_22_2),
		.out_wire_3_3(vertical_tile_7_22_to_tile_6_22_3),
		.in_wire_3_0(vertical_tile_6_22_to_tile_7_22_0),
		.in_wire_3_1(vertical_tile_6_22_to_tile_7_22_1),
		.in_wire_3_2(vertical_tile_6_22_to_tile_7_22_2),
		.in_wire_3_3(vertical_tile_6_22_to_tile_7_22_3),
		.out_wire_1_0(vertical_tile_7_22_to_tile_8_22_0),
		.out_wire_1_1(vertical_tile_7_22_to_tile_8_22_1),
		.out_wire_1_2(vertical_tile_7_22_to_tile_8_22_2),
		.out_wire_1_3(vertical_tile_7_22_to_tile_8_22_3),
		.in_wire_1_0(vertical_tile_8_22_to_tile_7_22_0),
		.in_wire_1_1(vertical_tile_8_22_to_tile_7_22_1),
		.in_wire_1_2(vertical_tile_8_22_to_tile_7_22_2),
		.in_wire_1_3(vertical_tile_8_22_to_tile_7_22_3),
		.out_wire_2_0(horizontal_tile_7_22_to_tile_7_21_0),
		.out_wire_2_1(horizontal_tile_7_22_to_tile_7_21_1),
		.out_wire_2_2(horizontal_tile_7_22_to_tile_7_21_2),
		.out_wire_2_3(horizontal_tile_7_22_to_tile_7_21_3),
		.in_wire_2_0(horizontal_tile_7_21_to_tile_7_22_0),
		.in_wire_2_1(horizontal_tile_7_21_to_tile_7_22_1),
		.in_wire_2_2(horizontal_tile_7_21_to_tile_7_22_2),
		.in_wire_2_3(horizontal_tile_7_21_to_tile_7_22_3),
		.out_wire_0_0(horizontal_tile_7_22_to_tile_7_23_0),
		.out_wire_0_1(horizontal_tile_7_22_to_tile_7_23_1),
		.out_wire_0_2(horizontal_tile_7_22_to_tile_7_23_2),
		.out_wire_0_3(horizontal_tile_7_22_to_tile_7_23_3),
		.in_wire_0_0(horizontal_tile_7_23_to_tile_7_22_0),
		.in_wire_0_1(horizontal_tile_7_23_to_tile_7_22_1),
		.in_wire_0_2(horizontal_tile_7_23_to_tile_7_22_2),
		.in_wire_0_3(horizontal_tile_7_23_to_tile_7_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(247)
	);

	pe_tile pe_tile_7_23(
		.out_wire_3_0(vertical_tile_7_23_to_tile_6_23_0),
		.out_wire_3_1(vertical_tile_7_23_to_tile_6_23_1),
		.out_wire_3_2(vertical_tile_7_23_to_tile_6_23_2),
		.out_wire_3_3(vertical_tile_7_23_to_tile_6_23_3),
		.in_wire_3_0(vertical_tile_6_23_to_tile_7_23_0),
		.in_wire_3_1(vertical_tile_6_23_to_tile_7_23_1),
		.in_wire_3_2(vertical_tile_6_23_to_tile_7_23_2),
		.in_wire_3_3(vertical_tile_6_23_to_tile_7_23_3),
		.out_wire_1_0(vertical_tile_7_23_to_tile_8_23_0),
		.out_wire_1_1(vertical_tile_7_23_to_tile_8_23_1),
		.out_wire_1_2(vertical_tile_7_23_to_tile_8_23_2),
		.out_wire_1_3(vertical_tile_7_23_to_tile_8_23_3),
		.in_wire_1_0(vertical_tile_8_23_to_tile_7_23_0),
		.in_wire_1_1(vertical_tile_8_23_to_tile_7_23_1),
		.in_wire_1_2(vertical_tile_8_23_to_tile_7_23_2),
		.in_wire_1_3(vertical_tile_8_23_to_tile_7_23_3),
		.out_wire_2_0(horizontal_tile_7_23_to_tile_7_22_0),
		.out_wire_2_1(horizontal_tile_7_23_to_tile_7_22_1),
		.out_wire_2_2(horizontal_tile_7_23_to_tile_7_22_2),
		.out_wire_2_3(horizontal_tile_7_23_to_tile_7_22_3),
		.in_wire_2_0(horizontal_tile_7_22_to_tile_7_23_0),
		.in_wire_2_1(horizontal_tile_7_22_to_tile_7_23_1),
		.in_wire_2_2(horizontal_tile_7_22_to_tile_7_23_2),
		.in_wire_2_3(horizontal_tile_7_22_to_tile_7_23_3),
		.out_wire_0_0(horizontal_tile_7_23_to_tile_7_24_0),
		.out_wire_0_1(horizontal_tile_7_23_to_tile_7_24_1),
		.out_wire_0_2(horizontal_tile_7_23_to_tile_7_24_2),
		.out_wire_0_3(horizontal_tile_7_23_to_tile_7_24_3),
		.in_wire_0_0(horizontal_tile_7_24_to_tile_7_23_0),
		.in_wire_0_1(horizontal_tile_7_24_to_tile_7_23_1),
		.in_wire_0_2(horizontal_tile_7_24_to_tile_7_23_2),
		.in_wire_0_3(horizontal_tile_7_24_to_tile_7_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(248)
	);

	pe_tile pe_tile_7_24(
		.out_wire_3_0(vertical_tile_7_24_to_tile_6_24_0),
		.out_wire_3_1(vertical_tile_7_24_to_tile_6_24_1),
		.out_wire_3_2(vertical_tile_7_24_to_tile_6_24_2),
		.out_wire_3_3(vertical_tile_7_24_to_tile_6_24_3),
		.in_wire_3_0(vertical_tile_6_24_to_tile_7_24_0),
		.in_wire_3_1(vertical_tile_6_24_to_tile_7_24_1),
		.in_wire_3_2(vertical_tile_6_24_to_tile_7_24_2),
		.in_wire_3_3(vertical_tile_6_24_to_tile_7_24_3),
		.out_wire_1_0(vertical_tile_7_24_to_tile_8_24_0),
		.out_wire_1_1(vertical_tile_7_24_to_tile_8_24_1),
		.out_wire_1_2(vertical_tile_7_24_to_tile_8_24_2),
		.out_wire_1_3(vertical_tile_7_24_to_tile_8_24_3),
		.in_wire_1_0(vertical_tile_8_24_to_tile_7_24_0),
		.in_wire_1_1(vertical_tile_8_24_to_tile_7_24_1),
		.in_wire_1_2(vertical_tile_8_24_to_tile_7_24_2),
		.in_wire_1_3(vertical_tile_8_24_to_tile_7_24_3),
		.out_wire_2_0(horizontal_tile_7_24_to_tile_7_23_0),
		.out_wire_2_1(horizontal_tile_7_24_to_tile_7_23_1),
		.out_wire_2_2(horizontal_tile_7_24_to_tile_7_23_2),
		.out_wire_2_3(horizontal_tile_7_24_to_tile_7_23_3),
		.in_wire_2_0(horizontal_tile_7_23_to_tile_7_24_0),
		.in_wire_2_1(horizontal_tile_7_23_to_tile_7_24_1),
		.in_wire_2_2(horizontal_tile_7_23_to_tile_7_24_2),
		.in_wire_2_3(horizontal_tile_7_23_to_tile_7_24_3),
		.out_wire_0_0(horizontal_tile_7_24_to_tile_7_25_0),
		.out_wire_0_1(horizontal_tile_7_24_to_tile_7_25_1),
		.out_wire_0_2(horizontal_tile_7_24_to_tile_7_25_2),
		.out_wire_0_3(horizontal_tile_7_24_to_tile_7_25_3),
		.in_wire_0_0(horizontal_tile_7_25_to_tile_7_24_0),
		.in_wire_0_1(horizontal_tile_7_25_to_tile_7_24_1),
		.in_wire_0_2(horizontal_tile_7_25_to_tile_7_24_2),
		.in_wire_0_3(horizontal_tile_7_25_to_tile_7_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(249)
	);

	pe_tile pe_tile_7_25(
		.out_wire_3_0(vertical_tile_7_25_to_tile_6_25_0),
		.out_wire_3_1(vertical_tile_7_25_to_tile_6_25_1),
		.out_wire_3_2(vertical_tile_7_25_to_tile_6_25_2),
		.out_wire_3_3(vertical_tile_7_25_to_tile_6_25_3),
		.in_wire_3_0(vertical_tile_6_25_to_tile_7_25_0),
		.in_wire_3_1(vertical_tile_6_25_to_tile_7_25_1),
		.in_wire_3_2(vertical_tile_6_25_to_tile_7_25_2),
		.in_wire_3_3(vertical_tile_6_25_to_tile_7_25_3),
		.out_wire_1_0(vertical_tile_7_25_to_tile_8_25_0),
		.out_wire_1_1(vertical_tile_7_25_to_tile_8_25_1),
		.out_wire_1_2(vertical_tile_7_25_to_tile_8_25_2),
		.out_wire_1_3(vertical_tile_7_25_to_tile_8_25_3),
		.in_wire_1_0(vertical_tile_8_25_to_tile_7_25_0),
		.in_wire_1_1(vertical_tile_8_25_to_tile_7_25_1),
		.in_wire_1_2(vertical_tile_8_25_to_tile_7_25_2),
		.in_wire_1_3(vertical_tile_8_25_to_tile_7_25_3),
		.out_wire_2_0(horizontal_tile_7_25_to_tile_7_24_0),
		.out_wire_2_1(horizontal_tile_7_25_to_tile_7_24_1),
		.out_wire_2_2(horizontal_tile_7_25_to_tile_7_24_2),
		.out_wire_2_3(horizontal_tile_7_25_to_tile_7_24_3),
		.in_wire_2_0(horizontal_tile_7_24_to_tile_7_25_0),
		.in_wire_2_1(horizontal_tile_7_24_to_tile_7_25_1),
		.in_wire_2_2(horizontal_tile_7_24_to_tile_7_25_2),
		.in_wire_2_3(horizontal_tile_7_24_to_tile_7_25_3),
		.out_wire_0_0(horizontal_tile_7_25_to_tile_7_26_0),
		.out_wire_0_1(horizontal_tile_7_25_to_tile_7_26_1),
		.out_wire_0_2(horizontal_tile_7_25_to_tile_7_26_2),
		.out_wire_0_3(horizontal_tile_7_25_to_tile_7_26_3),
		.in_wire_0_0(horizontal_tile_7_26_to_tile_7_25_0),
		.in_wire_0_1(horizontal_tile_7_26_to_tile_7_25_1),
		.in_wire_0_2(horizontal_tile_7_26_to_tile_7_25_2),
		.in_wire_0_3(horizontal_tile_7_26_to_tile_7_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(250)
	);

	pe_tile pe_tile_7_26(
		.out_wire_3_0(vertical_tile_7_26_to_tile_6_26_0),
		.out_wire_3_1(vertical_tile_7_26_to_tile_6_26_1),
		.out_wire_3_2(vertical_tile_7_26_to_tile_6_26_2),
		.out_wire_3_3(vertical_tile_7_26_to_tile_6_26_3),
		.in_wire_3_0(vertical_tile_6_26_to_tile_7_26_0),
		.in_wire_3_1(vertical_tile_6_26_to_tile_7_26_1),
		.in_wire_3_2(vertical_tile_6_26_to_tile_7_26_2),
		.in_wire_3_3(vertical_tile_6_26_to_tile_7_26_3),
		.out_wire_1_0(vertical_tile_7_26_to_tile_8_26_0),
		.out_wire_1_1(vertical_tile_7_26_to_tile_8_26_1),
		.out_wire_1_2(vertical_tile_7_26_to_tile_8_26_2),
		.out_wire_1_3(vertical_tile_7_26_to_tile_8_26_3),
		.in_wire_1_0(vertical_tile_8_26_to_tile_7_26_0),
		.in_wire_1_1(vertical_tile_8_26_to_tile_7_26_1),
		.in_wire_1_2(vertical_tile_8_26_to_tile_7_26_2),
		.in_wire_1_3(vertical_tile_8_26_to_tile_7_26_3),
		.out_wire_2_0(horizontal_tile_7_26_to_tile_7_25_0),
		.out_wire_2_1(horizontal_tile_7_26_to_tile_7_25_1),
		.out_wire_2_2(horizontal_tile_7_26_to_tile_7_25_2),
		.out_wire_2_3(horizontal_tile_7_26_to_tile_7_25_3),
		.in_wire_2_0(horizontal_tile_7_25_to_tile_7_26_0),
		.in_wire_2_1(horizontal_tile_7_25_to_tile_7_26_1),
		.in_wire_2_2(horizontal_tile_7_25_to_tile_7_26_2),
		.in_wire_2_3(horizontal_tile_7_25_to_tile_7_26_3),
		.out_wire_0_0(horizontal_tile_7_26_to_tile_7_27_0),
		.out_wire_0_1(horizontal_tile_7_26_to_tile_7_27_1),
		.out_wire_0_2(horizontal_tile_7_26_to_tile_7_27_2),
		.out_wire_0_3(horizontal_tile_7_26_to_tile_7_27_3),
		.in_wire_0_0(horizontal_tile_7_27_to_tile_7_26_0),
		.in_wire_0_1(horizontal_tile_7_27_to_tile_7_26_1),
		.in_wire_0_2(horizontal_tile_7_27_to_tile_7_26_2),
		.in_wire_0_3(horizontal_tile_7_27_to_tile_7_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(251)
	);

	pe_tile pe_tile_7_27(
		.out_wire_3_0(vertical_tile_7_27_to_tile_6_27_0),
		.out_wire_3_1(vertical_tile_7_27_to_tile_6_27_1),
		.out_wire_3_2(vertical_tile_7_27_to_tile_6_27_2),
		.out_wire_3_3(vertical_tile_7_27_to_tile_6_27_3),
		.in_wire_3_0(vertical_tile_6_27_to_tile_7_27_0),
		.in_wire_3_1(vertical_tile_6_27_to_tile_7_27_1),
		.in_wire_3_2(vertical_tile_6_27_to_tile_7_27_2),
		.in_wire_3_3(vertical_tile_6_27_to_tile_7_27_3),
		.out_wire_1_0(vertical_tile_7_27_to_tile_8_27_0),
		.out_wire_1_1(vertical_tile_7_27_to_tile_8_27_1),
		.out_wire_1_2(vertical_tile_7_27_to_tile_8_27_2),
		.out_wire_1_3(vertical_tile_7_27_to_tile_8_27_3),
		.in_wire_1_0(vertical_tile_8_27_to_tile_7_27_0),
		.in_wire_1_1(vertical_tile_8_27_to_tile_7_27_1),
		.in_wire_1_2(vertical_tile_8_27_to_tile_7_27_2),
		.in_wire_1_3(vertical_tile_8_27_to_tile_7_27_3),
		.out_wire_2_0(horizontal_tile_7_27_to_tile_7_26_0),
		.out_wire_2_1(horizontal_tile_7_27_to_tile_7_26_1),
		.out_wire_2_2(horizontal_tile_7_27_to_tile_7_26_2),
		.out_wire_2_3(horizontal_tile_7_27_to_tile_7_26_3),
		.in_wire_2_0(horizontal_tile_7_26_to_tile_7_27_0),
		.in_wire_2_1(horizontal_tile_7_26_to_tile_7_27_1),
		.in_wire_2_2(horizontal_tile_7_26_to_tile_7_27_2),
		.in_wire_2_3(horizontal_tile_7_26_to_tile_7_27_3),
		.out_wire_0_0(horizontal_tile_7_27_to_tile_7_28_0),
		.out_wire_0_1(horizontal_tile_7_27_to_tile_7_28_1),
		.out_wire_0_2(horizontal_tile_7_27_to_tile_7_28_2),
		.out_wire_0_3(horizontal_tile_7_27_to_tile_7_28_3),
		.in_wire_0_0(horizontal_tile_7_28_to_tile_7_27_0),
		.in_wire_0_1(horizontal_tile_7_28_to_tile_7_27_1),
		.in_wire_0_2(horizontal_tile_7_28_to_tile_7_27_2),
		.in_wire_0_3(horizontal_tile_7_28_to_tile_7_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(252)
	);

	pe_tile pe_tile_7_28(
		.out_wire_3_0(vertical_tile_7_28_to_tile_6_28_0),
		.out_wire_3_1(vertical_tile_7_28_to_tile_6_28_1),
		.out_wire_3_2(vertical_tile_7_28_to_tile_6_28_2),
		.out_wire_3_3(vertical_tile_7_28_to_tile_6_28_3),
		.in_wire_3_0(vertical_tile_6_28_to_tile_7_28_0),
		.in_wire_3_1(vertical_tile_6_28_to_tile_7_28_1),
		.in_wire_3_2(vertical_tile_6_28_to_tile_7_28_2),
		.in_wire_3_3(vertical_tile_6_28_to_tile_7_28_3),
		.out_wire_1_0(vertical_tile_7_28_to_tile_8_28_0),
		.out_wire_1_1(vertical_tile_7_28_to_tile_8_28_1),
		.out_wire_1_2(vertical_tile_7_28_to_tile_8_28_2),
		.out_wire_1_3(vertical_tile_7_28_to_tile_8_28_3),
		.in_wire_1_0(vertical_tile_8_28_to_tile_7_28_0),
		.in_wire_1_1(vertical_tile_8_28_to_tile_7_28_1),
		.in_wire_1_2(vertical_tile_8_28_to_tile_7_28_2),
		.in_wire_1_3(vertical_tile_8_28_to_tile_7_28_3),
		.out_wire_2_0(horizontal_tile_7_28_to_tile_7_27_0),
		.out_wire_2_1(horizontal_tile_7_28_to_tile_7_27_1),
		.out_wire_2_2(horizontal_tile_7_28_to_tile_7_27_2),
		.out_wire_2_3(horizontal_tile_7_28_to_tile_7_27_3),
		.in_wire_2_0(horizontal_tile_7_27_to_tile_7_28_0),
		.in_wire_2_1(horizontal_tile_7_27_to_tile_7_28_1),
		.in_wire_2_2(horizontal_tile_7_27_to_tile_7_28_2),
		.in_wire_2_3(horizontal_tile_7_27_to_tile_7_28_3),
		.out_wire_0_0(horizontal_tile_7_28_to_tile_7_29_0),
		.out_wire_0_1(horizontal_tile_7_28_to_tile_7_29_1),
		.out_wire_0_2(horizontal_tile_7_28_to_tile_7_29_2),
		.out_wire_0_3(horizontal_tile_7_28_to_tile_7_29_3),
		.in_wire_0_0(horizontal_tile_7_29_to_tile_7_28_0),
		.in_wire_0_1(horizontal_tile_7_29_to_tile_7_28_1),
		.in_wire_0_2(horizontal_tile_7_29_to_tile_7_28_2),
		.in_wire_0_3(horizontal_tile_7_29_to_tile_7_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(253)
	);

	pe_tile pe_tile_7_29(
		.out_wire_3_0(vertical_tile_7_29_to_tile_6_29_0),
		.out_wire_3_1(vertical_tile_7_29_to_tile_6_29_1),
		.out_wire_3_2(vertical_tile_7_29_to_tile_6_29_2),
		.out_wire_3_3(vertical_tile_7_29_to_tile_6_29_3),
		.in_wire_3_0(vertical_tile_6_29_to_tile_7_29_0),
		.in_wire_3_1(vertical_tile_6_29_to_tile_7_29_1),
		.in_wire_3_2(vertical_tile_6_29_to_tile_7_29_2),
		.in_wire_3_3(vertical_tile_6_29_to_tile_7_29_3),
		.out_wire_1_0(vertical_tile_7_29_to_tile_8_29_0),
		.out_wire_1_1(vertical_tile_7_29_to_tile_8_29_1),
		.out_wire_1_2(vertical_tile_7_29_to_tile_8_29_2),
		.out_wire_1_3(vertical_tile_7_29_to_tile_8_29_3),
		.in_wire_1_0(vertical_tile_8_29_to_tile_7_29_0),
		.in_wire_1_1(vertical_tile_8_29_to_tile_7_29_1),
		.in_wire_1_2(vertical_tile_8_29_to_tile_7_29_2),
		.in_wire_1_3(vertical_tile_8_29_to_tile_7_29_3),
		.out_wire_2_0(horizontal_tile_7_29_to_tile_7_28_0),
		.out_wire_2_1(horizontal_tile_7_29_to_tile_7_28_1),
		.out_wire_2_2(horizontal_tile_7_29_to_tile_7_28_2),
		.out_wire_2_3(horizontal_tile_7_29_to_tile_7_28_3),
		.in_wire_2_0(horizontal_tile_7_28_to_tile_7_29_0),
		.in_wire_2_1(horizontal_tile_7_28_to_tile_7_29_1),
		.in_wire_2_2(horizontal_tile_7_28_to_tile_7_29_2),
		.in_wire_2_3(horizontal_tile_7_28_to_tile_7_29_3),
		.out_wire_0_0(horizontal_tile_7_29_to_tile_7_30_0),
		.out_wire_0_1(horizontal_tile_7_29_to_tile_7_30_1),
		.out_wire_0_2(horizontal_tile_7_29_to_tile_7_30_2),
		.out_wire_0_3(horizontal_tile_7_29_to_tile_7_30_3),
		.in_wire_0_0(horizontal_tile_7_30_to_tile_7_29_0),
		.in_wire_0_1(horizontal_tile_7_30_to_tile_7_29_1),
		.in_wire_0_2(horizontal_tile_7_30_to_tile_7_29_2),
		.in_wire_0_3(horizontal_tile_7_30_to_tile_7_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(254)
	);

	pe_tile pe_tile_7_30(
		.out_wire_3_0(vertical_tile_7_30_to_tile_6_30_0),
		.out_wire_3_1(vertical_tile_7_30_to_tile_6_30_1),
		.out_wire_3_2(vertical_tile_7_30_to_tile_6_30_2),
		.out_wire_3_3(vertical_tile_7_30_to_tile_6_30_3),
		.in_wire_3_0(vertical_tile_6_30_to_tile_7_30_0),
		.in_wire_3_1(vertical_tile_6_30_to_tile_7_30_1),
		.in_wire_3_2(vertical_tile_6_30_to_tile_7_30_2),
		.in_wire_3_3(vertical_tile_6_30_to_tile_7_30_3),
		.out_wire_1_0(vertical_tile_7_30_to_tile_8_30_0),
		.out_wire_1_1(vertical_tile_7_30_to_tile_8_30_1),
		.out_wire_1_2(vertical_tile_7_30_to_tile_8_30_2),
		.out_wire_1_3(vertical_tile_7_30_to_tile_8_30_3),
		.in_wire_1_0(vertical_tile_8_30_to_tile_7_30_0),
		.in_wire_1_1(vertical_tile_8_30_to_tile_7_30_1),
		.in_wire_1_2(vertical_tile_8_30_to_tile_7_30_2),
		.in_wire_1_3(vertical_tile_8_30_to_tile_7_30_3),
		.out_wire_2_0(horizontal_tile_7_30_to_tile_7_29_0),
		.out_wire_2_1(horizontal_tile_7_30_to_tile_7_29_1),
		.out_wire_2_2(horizontal_tile_7_30_to_tile_7_29_2),
		.out_wire_2_3(horizontal_tile_7_30_to_tile_7_29_3),
		.in_wire_2_0(horizontal_tile_7_29_to_tile_7_30_0),
		.in_wire_2_1(horizontal_tile_7_29_to_tile_7_30_1),
		.in_wire_2_2(horizontal_tile_7_29_to_tile_7_30_2),
		.in_wire_2_3(horizontal_tile_7_29_to_tile_7_30_3),
		.out_wire_0_0(horizontal_tile_7_30_to_tile_7_31_0),
		.out_wire_0_1(horizontal_tile_7_30_to_tile_7_31_1),
		.out_wire_0_2(horizontal_tile_7_30_to_tile_7_31_2),
		.out_wire_0_3(horizontal_tile_7_30_to_tile_7_31_3),
		.in_wire_0_0(horizontal_tile_7_31_to_tile_7_30_0),
		.in_wire_0_1(horizontal_tile_7_31_to_tile_7_30_1),
		.in_wire_0_2(horizontal_tile_7_31_to_tile_7_30_2),
		.in_wire_0_3(horizontal_tile_7_31_to_tile_7_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(255)
	);

	pe_tile_right pe_tile_7_31(
		.out_wire_3_0(vertical_tile_7_31_to_tile_6_31_0),
		.out_wire_3_1(vertical_tile_7_31_to_tile_6_31_1),
		.out_wire_3_2(vertical_tile_7_31_to_tile_6_31_2),
		.out_wire_3_3(vertical_tile_7_31_to_tile_6_31_3),
		.in_wire_3_0(vertical_tile_6_31_to_tile_7_31_0),
		.in_wire_3_1(vertical_tile_6_31_to_tile_7_31_1),
		.in_wire_3_2(vertical_tile_6_31_to_tile_7_31_2),
		.in_wire_3_3(vertical_tile_6_31_to_tile_7_31_3),
		.out_wire_1_0(vertical_tile_7_31_to_tile_8_31_0),
		.out_wire_1_1(vertical_tile_7_31_to_tile_8_31_1),
		.out_wire_1_2(vertical_tile_7_31_to_tile_8_31_2),
		.out_wire_1_3(vertical_tile_7_31_to_tile_8_31_3),
		.in_wire_1_0(vertical_tile_8_31_to_tile_7_31_0),
		.in_wire_1_1(vertical_tile_8_31_to_tile_7_31_1),
		.in_wire_1_2(vertical_tile_8_31_to_tile_7_31_2),
		.in_wire_1_3(vertical_tile_8_31_to_tile_7_31_3),
		.out_wire_2_0(horizontal_tile_7_31_to_tile_7_30_0),
		.out_wire_2_1(horizontal_tile_7_31_to_tile_7_30_1),
		.out_wire_2_2(horizontal_tile_7_31_to_tile_7_30_2),
		.out_wire_2_3(horizontal_tile_7_31_to_tile_7_30_3),
		.in_wire_2_0(horizontal_tile_7_30_to_tile_7_31_0),
		.in_wire_2_1(horizontal_tile_7_30_to_tile_7_31_1),
		.in_wire_2_2(horizontal_tile_7_30_to_tile_7_31_2),
		.in_wire_2_3(horizontal_tile_7_30_to_tile_7_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(256)
	);

	pe_tile_left pe_tile_8_0(
		.out_wire_3_0(vertical_tile_8_0_to_tile_7_0_0),
		.out_wire_3_1(vertical_tile_8_0_to_tile_7_0_1),
		.out_wire_3_2(vertical_tile_8_0_to_tile_7_0_2),
		.out_wire_3_3(vertical_tile_8_0_to_tile_7_0_3),
		.in_wire_3_0(vertical_tile_7_0_to_tile_8_0_0),
		.in_wire_3_1(vertical_tile_7_0_to_tile_8_0_1),
		.in_wire_3_2(vertical_tile_7_0_to_tile_8_0_2),
		.in_wire_3_3(vertical_tile_7_0_to_tile_8_0_3),
		.out_wire_1_0(vertical_tile_8_0_to_tile_9_0_0),
		.out_wire_1_1(vertical_tile_8_0_to_tile_9_0_1),
		.out_wire_1_2(vertical_tile_8_0_to_tile_9_0_2),
		.out_wire_1_3(vertical_tile_8_0_to_tile_9_0_3),
		.in_wire_1_0(vertical_tile_9_0_to_tile_8_0_0),
		.in_wire_1_1(vertical_tile_9_0_to_tile_8_0_1),
		.in_wire_1_2(vertical_tile_9_0_to_tile_8_0_2),
		.in_wire_1_3(vertical_tile_9_0_to_tile_8_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_8_0_to_tile_8_1_0),
		.out_wire_0_1(horizontal_tile_8_0_to_tile_8_1_1),
		.out_wire_0_2(horizontal_tile_8_0_to_tile_8_1_2),
		.out_wire_0_3(horizontal_tile_8_0_to_tile_8_1_3),
		.in_wire_0_0(horizontal_tile_8_1_to_tile_8_0_0),
		.in_wire_0_1(horizontal_tile_8_1_to_tile_8_0_1),
		.in_wire_0_2(horizontal_tile_8_1_to_tile_8_0_2),
		.in_wire_0_3(horizontal_tile_8_1_to_tile_8_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(257)
	);

	pe_tile pe_tile_8_1(
		.out_wire_3_0(vertical_tile_8_1_to_tile_7_1_0),
		.out_wire_3_1(vertical_tile_8_1_to_tile_7_1_1),
		.out_wire_3_2(vertical_tile_8_1_to_tile_7_1_2),
		.out_wire_3_3(vertical_tile_8_1_to_tile_7_1_3),
		.in_wire_3_0(vertical_tile_7_1_to_tile_8_1_0),
		.in_wire_3_1(vertical_tile_7_1_to_tile_8_1_1),
		.in_wire_3_2(vertical_tile_7_1_to_tile_8_1_2),
		.in_wire_3_3(vertical_tile_7_1_to_tile_8_1_3),
		.out_wire_1_0(vertical_tile_8_1_to_tile_9_1_0),
		.out_wire_1_1(vertical_tile_8_1_to_tile_9_1_1),
		.out_wire_1_2(vertical_tile_8_1_to_tile_9_1_2),
		.out_wire_1_3(vertical_tile_8_1_to_tile_9_1_3),
		.in_wire_1_0(vertical_tile_9_1_to_tile_8_1_0),
		.in_wire_1_1(vertical_tile_9_1_to_tile_8_1_1),
		.in_wire_1_2(vertical_tile_9_1_to_tile_8_1_2),
		.in_wire_1_3(vertical_tile_9_1_to_tile_8_1_3),
		.out_wire_2_0(horizontal_tile_8_1_to_tile_8_0_0),
		.out_wire_2_1(horizontal_tile_8_1_to_tile_8_0_1),
		.out_wire_2_2(horizontal_tile_8_1_to_tile_8_0_2),
		.out_wire_2_3(horizontal_tile_8_1_to_tile_8_0_3),
		.in_wire_2_0(horizontal_tile_8_0_to_tile_8_1_0),
		.in_wire_2_1(horizontal_tile_8_0_to_tile_8_1_1),
		.in_wire_2_2(horizontal_tile_8_0_to_tile_8_1_2),
		.in_wire_2_3(horizontal_tile_8_0_to_tile_8_1_3),
		.out_wire_0_0(horizontal_tile_8_1_to_tile_8_2_0),
		.out_wire_0_1(horizontal_tile_8_1_to_tile_8_2_1),
		.out_wire_0_2(horizontal_tile_8_1_to_tile_8_2_2),
		.out_wire_0_3(horizontal_tile_8_1_to_tile_8_2_3),
		.in_wire_0_0(horizontal_tile_8_2_to_tile_8_1_0),
		.in_wire_0_1(horizontal_tile_8_2_to_tile_8_1_1),
		.in_wire_0_2(horizontal_tile_8_2_to_tile_8_1_2),
		.in_wire_0_3(horizontal_tile_8_2_to_tile_8_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(258)
	);

	pe_tile pe_tile_8_2(
		.out_wire_3_0(vertical_tile_8_2_to_tile_7_2_0),
		.out_wire_3_1(vertical_tile_8_2_to_tile_7_2_1),
		.out_wire_3_2(vertical_tile_8_2_to_tile_7_2_2),
		.out_wire_3_3(vertical_tile_8_2_to_tile_7_2_3),
		.in_wire_3_0(vertical_tile_7_2_to_tile_8_2_0),
		.in_wire_3_1(vertical_tile_7_2_to_tile_8_2_1),
		.in_wire_3_2(vertical_tile_7_2_to_tile_8_2_2),
		.in_wire_3_3(vertical_tile_7_2_to_tile_8_2_3),
		.out_wire_1_0(vertical_tile_8_2_to_tile_9_2_0),
		.out_wire_1_1(vertical_tile_8_2_to_tile_9_2_1),
		.out_wire_1_2(vertical_tile_8_2_to_tile_9_2_2),
		.out_wire_1_3(vertical_tile_8_2_to_tile_9_2_3),
		.in_wire_1_0(vertical_tile_9_2_to_tile_8_2_0),
		.in_wire_1_1(vertical_tile_9_2_to_tile_8_2_1),
		.in_wire_1_2(vertical_tile_9_2_to_tile_8_2_2),
		.in_wire_1_3(vertical_tile_9_2_to_tile_8_2_3),
		.out_wire_2_0(horizontal_tile_8_2_to_tile_8_1_0),
		.out_wire_2_1(horizontal_tile_8_2_to_tile_8_1_1),
		.out_wire_2_2(horizontal_tile_8_2_to_tile_8_1_2),
		.out_wire_2_3(horizontal_tile_8_2_to_tile_8_1_3),
		.in_wire_2_0(horizontal_tile_8_1_to_tile_8_2_0),
		.in_wire_2_1(horizontal_tile_8_1_to_tile_8_2_1),
		.in_wire_2_2(horizontal_tile_8_1_to_tile_8_2_2),
		.in_wire_2_3(horizontal_tile_8_1_to_tile_8_2_3),
		.out_wire_0_0(horizontal_tile_8_2_to_tile_8_3_0),
		.out_wire_0_1(horizontal_tile_8_2_to_tile_8_3_1),
		.out_wire_0_2(horizontal_tile_8_2_to_tile_8_3_2),
		.out_wire_0_3(horizontal_tile_8_2_to_tile_8_3_3),
		.in_wire_0_0(horizontal_tile_8_3_to_tile_8_2_0),
		.in_wire_0_1(horizontal_tile_8_3_to_tile_8_2_1),
		.in_wire_0_2(horizontal_tile_8_3_to_tile_8_2_2),
		.in_wire_0_3(horizontal_tile_8_3_to_tile_8_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(259)
	);

	pe_tile pe_tile_8_3(
		.out_wire_3_0(vertical_tile_8_3_to_tile_7_3_0),
		.out_wire_3_1(vertical_tile_8_3_to_tile_7_3_1),
		.out_wire_3_2(vertical_tile_8_3_to_tile_7_3_2),
		.out_wire_3_3(vertical_tile_8_3_to_tile_7_3_3),
		.in_wire_3_0(vertical_tile_7_3_to_tile_8_3_0),
		.in_wire_3_1(vertical_tile_7_3_to_tile_8_3_1),
		.in_wire_3_2(vertical_tile_7_3_to_tile_8_3_2),
		.in_wire_3_3(vertical_tile_7_3_to_tile_8_3_3),
		.out_wire_1_0(vertical_tile_8_3_to_tile_9_3_0),
		.out_wire_1_1(vertical_tile_8_3_to_tile_9_3_1),
		.out_wire_1_2(vertical_tile_8_3_to_tile_9_3_2),
		.out_wire_1_3(vertical_tile_8_3_to_tile_9_3_3),
		.in_wire_1_0(vertical_tile_9_3_to_tile_8_3_0),
		.in_wire_1_1(vertical_tile_9_3_to_tile_8_3_1),
		.in_wire_1_2(vertical_tile_9_3_to_tile_8_3_2),
		.in_wire_1_3(vertical_tile_9_3_to_tile_8_3_3),
		.out_wire_2_0(horizontal_tile_8_3_to_tile_8_2_0),
		.out_wire_2_1(horizontal_tile_8_3_to_tile_8_2_1),
		.out_wire_2_2(horizontal_tile_8_3_to_tile_8_2_2),
		.out_wire_2_3(horizontal_tile_8_3_to_tile_8_2_3),
		.in_wire_2_0(horizontal_tile_8_2_to_tile_8_3_0),
		.in_wire_2_1(horizontal_tile_8_2_to_tile_8_3_1),
		.in_wire_2_2(horizontal_tile_8_2_to_tile_8_3_2),
		.in_wire_2_3(horizontal_tile_8_2_to_tile_8_3_3),
		.out_wire_0_0(horizontal_tile_8_3_to_tile_8_4_0),
		.out_wire_0_1(horizontal_tile_8_3_to_tile_8_4_1),
		.out_wire_0_2(horizontal_tile_8_3_to_tile_8_4_2),
		.out_wire_0_3(horizontal_tile_8_3_to_tile_8_4_3),
		.in_wire_0_0(horizontal_tile_8_4_to_tile_8_3_0),
		.in_wire_0_1(horizontal_tile_8_4_to_tile_8_3_1),
		.in_wire_0_2(horizontal_tile_8_4_to_tile_8_3_2),
		.in_wire_0_3(horizontal_tile_8_4_to_tile_8_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(260)
	);

	pe_tile pe_tile_8_4(
		.out_wire_3_0(vertical_tile_8_4_to_tile_7_4_0),
		.out_wire_3_1(vertical_tile_8_4_to_tile_7_4_1),
		.out_wire_3_2(vertical_tile_8_4_to_tile_7_4_2),
		.out_wire_3_3(vertical_tile_8_4_to_tile_7_4_3),
		.in_wire_3_0(vertical_tile_7_4_to_tile_8_4_0),
		.in_wire_3_1(vertical_tile_7_4_to_tile_8_4_1),
		.in_wire_3_2(vertical_tile_7_4_to_tile_8_4_2),
		.in_wire_3_3(vertical_tile_7_4_to_tile_8_4_3),
		.out_wire_1_0(vertical_tile_8_4_to_tile_9_4_0),
		.out_wire_1_1(vertical_tile_8_4_to_tile_9_4_1),
		.out_wire_1_2(vertical_tile_8_4_to_tile_9_4_2),
		.out_wire_1_3(vertical_tile_8_4_to_tile_9_4_3),
		.in_wire_1_0(vertical_tile_9_4_to_tile_8_4_0),
		.in_wire_1_1(vertical_tile_9_4_to_tile_8_4_1),
		.in_wire_1_2(vertical_tile_9_4_to_tile_8_4_2),
		.in_wire_1_3(vertical_tile_9_4_to_tile_8_4_3),
		.out_wire_2_0(horizontal_tile_8_4_to_tile_8_3_0),
		.out_wire_2_1(horizontal_tile_8_4_to_tile_8_3_1),
		.out_wire_2_2(horizontal_tile_8_4_to_tile_8_3_2),
		.out_wire_2_3(horizontal_tile_8_4_to_tile_8_3_3),
		.in_wire_2_0(horizontal_tile_8_3_to_tile_8_4_0),
		.in_wire_2_1(horizontal_tile_8_3_to_tile_8_4_1),
		.in_wire_2_2(horizontal_tile_8_3_to_tile_8_4_2),
		.in_wire_2_3(horizontal_tile_8_3_to_tile_8_4_3),
		.out_wire_0_0(horizontal_tile_8_4_to_tile_8_5_0),
		.out_wire_0_1(horizontal_tile_8_4_to_tile_8_5_1),
		.out_wire_0_2(horizontal_tile_8_4_to_tile_8_5_2),
		.out_wire_0_3(horizontal_tile_8_4_to_tile_8_5_3),
		.in_wire_0_0(horizontal_tile_8_5_to_tile_8_4_0),
		.in_wire_0_1(horizontal_tile_8_5_to_tile_8_4_1),
		.in_wire_0_2(horizontal_tile_8_5_to_tile_8_4_2),
		.in_wire_0_3(horizontal_tile_8_5_to_tile_8_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(261)
	);

	pe_tile pe_tile_8_5(
		.out_wire_3_0(vertical_tile_8_5_to_tile_7_5_0),
		.out_wire_3_1(vertical_tile_8_5_to_tile_7_5_1),
		.out_wire_3_2(vertical_tile_8_5_to_tile_7_5_2),
		.out_wire_3_3(vertical_tile_8_5_to_tile_7_5_3),
		.in_wire_3_0(vertical_tile_7_5_to_tile_8_5_0),
		.in_wire_3_1(vertical_tile_7_5_to_tile_8_5_1),
		.in_wire_3_2(vertical_tile_7_5_to_tile_8_5_2),
		.in_wire_3_3(vertical_tile_7_5_to_tile_8_5_3),
		.out_wire_1_0(vertical_tile_8_5_to_tile_9_5_0),
		.out_wire_1_1(vertical_tile_8_5_to_tile_9_5_1),
		.out_wire_1_2(vertical_tile_8_5_to_tile_9_5_2),
		.out_wire_1_3(vertical_tile_8_5_to_tile_9_5_3),
		.in_wire_1_0(vertical_tile_9_5_to_tile_8_5_0),
		.in_wire_1_1(vertical_tile_9_5_to_tile_8_5_1),
		.in_wire_1_2(vertical_tile_9_5_to_tile_8_5_2),
		.in_wire_1_3(vertical_tile_9_5_to_tile_8_5_3),
		.out_wire_2_0(horizontal_tile_8_5_to_tile_8_4_0),
		.out_wire_2_1(horizontal_tile_8_5_to_tile_8_4_1),
		.out_wire_2_2(horizontal_tile_8_5_to_tile_8_4_2),
		.out_wire_2_3(horizontal_tile_8_5_to_tile_8_4_3),
		.in_wire_2_0(horizontal_tile_8_4_to_tile_8_5_0),
		.in_wire_2_1(horizontal_tile_8_4_to_tile_8_5_1),
		.in_wire_2_2(horizontal_tile_8_4_to_tile_8_5_2),
		.in_wire_2_3(horizontal_tile_8_4_to_tile_8_5_3),
		.out_wire_0_0(horizontal_tile_8_5_to_tile_8_6_0),
		.out_wire_0_1(horizontal_tile_8_5_to_tile_8_6_1),
		.out_wire_0_2(horizontal_tile_8_5_to_tile_8_6_2),
		.out_wire_0_3(horizontal_tile_8_5_to_tile_8_6_3),
		.in_wire_0_0(horizontal_tile_8_6_to_tile_8_5_0),
		.in_wire_0_1(horizontal_tile_8_6_to_tile_8_5_1),
		.in_wire_0_2(horizontal_tile_8_6_to_tile_8_5_2),
		.in_wire_0_3(horizontal_tile_8_6_to_tile_8_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(262)
	);

	pe_tile pe_tile_8_6(
		.out_wire_3_0(vertical_tile_8_6_to_tile_7_6_0),
		.out_wire_3_1(vertical_tile_8_6_to_tile_7_6_1),
		.out_wire_3_2(vertical_tile_8_6_to_tile_7_6_2),
		.out_wire_3_3(vertical_tile_8_6_to_tile_7_6_3),
		.in_wire_3_0(vertical_tile_7_6_to_tile_8_6_0),
		.in_wire_3_1(vertical_tile_7_6_to_tile_8_6_1),
		.in_wire_3_2(vertical_tile_7_6_to_tile_8_6_2),
		.in_wire_3_3(vertical_tile_7_6_to_tile_8_6_3),
		.out_wire_1_0(vertical_tile_8_6_to_tile_9_6_0),
		.out_wire_1_1(vertical_tile_8_6_to_tile_9_6_1),
		.out_wire_1_2(vertical_tile_8_6_to_tile_9_6_2),
		.out_wire_1_3(vertical_tile_8_6_to_tile_9_6_3),
		.in_wire_1_0(vertical_tile_9_6_to_tile_8_6_0),
		.in_wire_1_1(vertical_tile_9_6_to_tile_8_6_1),
		.in_wire_1_2(vertical_tile_9_6_to_tile_8_6_2),
		.in_wire_1_3(vertical_tile_9_6_to_tile_8_6_3),
		.out_wire_2_0(horizontal_tile_8_6_to_tile_8_5_0),
		.out_wire_2_1(horizontal_tile_8_6_to_tile_8_5_1),
		.out_wire_2_2(horizontal_tile_8_6_to_tile_8_5_2),
		.out_wire_2_3(horizontal_tile_8_6_to_tile_8_5_3),
		.in_wire_2_0(horizontal_tile_8_5_to_tile_8_6_0),
		.in_wire_2_1(horizontal_tile_8_5_to_tile_8_6_1),
		.in_wire_2_2(horizontal_tile_8_5_to_tile_8_6_2),
		.in_wire_2_3(horizontal_tile_8_5_to_tile_8_6_3),
		.out_wire_0_0(horizontal_tile_8_6_to_tile_8_7_0),
		.out_wire_0_1(horizontal_tile_8_6_to_tile_8_7_1),
		.out_wire_0_2(horizontal_tile_8_6_to_tile_8_7_2),
		.out_wire_0_3(horizontal_tile_8_6_to_tile_8_7_3),
		.in_wire_0_0(horizontal_tile_8_7_to_tile_8_6_0),
		.in_wire_0_1(horizontal_tile_8_7_to_tile_8_6_1),
		.in_wire_0_2(horizontal_tile_8_7_to_tile_8_6_2),
		.in_wire_0_3(horizontal_tile_8_7_to_tile_8_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(263)
	);

	pe_tile pe_tile_8_7(
		.out_wire_3_0(vertical_tile_8_7_to_tile_7_7_0),
		.out_wire_3_1(vertical_tile_8_7_to_tile_7_7_1),
		.out_wire_3_2(vertical_tile_8_7_to_tile_7_7_2),
		.out_wire_3_3(vertical_tile_8_7_to_tile_7_7_3),
		.in_wire_3_0(vertical_tile_7_7_to_tile_8_7_0),
		.in_wire_3_1(vertical_tile_7_7_to_tile_8_7_1),
		.in_wire_3_2(vertical_tile_7_7_to_tile_8_7_2),
		.in_wire_3_3(vertical_tile_7_7_to_tile_8_7_3),
		.out_wire_1_0(vertical_tile_8_7_to_tile_9_7_0),
		.out_wire_1_1(vertical_tile_8_7_to_tile_9_7_1),
		.out_wire_1_2(vertical_tile_8_7_to_tile_9_7_2),
		.out_wire_1_3(vertical_tile_8_7_to_tile_9_7_3),
		.in_wire_1_0(vertical_tile_9_7_to_tile_8_7_0),
		.in_wire_1_1(vertical_tile_9_7_to_tile_8_7_1),
		.in_wire_1_2(vertical_tile_9_7_to_tile_8_7_2),
		.in_wire_1_3(vertical_tile_9_7_to_tile_8_7_3),
		.out_wire_2_0(horizontal_tile_8_7_to_tile_8_6_0),
		.out_wire_2_1(horizontal_tile_8_7_to_tile_8_6_1),
		.out_wire_2_2(horizontal_tile_8_7_to_tile_8_6_2),
		.out_wire_2_3(horizontal_tile_8_7_to_tile_8_6_3),
		.in_wire_2_0(horizontal_tile_8_6_to_tile_8_7_0),
		.in_wire_2_1(horizontal_tile_8_6_to_tile_8_7_1),
		.in_wire_2_2(horizontal_tile_8_6_to_tile_8_7_2),
		.in_wire_2_3(horizontal_tile_8_6_to_tile_8_7_3),
		.out_wire_0_0(horizontal_tile_8_7_to_tile_8_8_0),
		.out_wire_0_1(horizontal_tile_8_7_to_tile_8_8_1),
		.out_wire_0_2(horizontal_tile_8_7_to_tile_8_8_2),
		.out_wire_0_3(horizontal_tile_8_7_to_tile_8_8_3),
		.in_wire_0_0(horizontal_tile_8_8_to_tile_8_7_0),
		.in_wire_0_1(horizontal_tile_8_8_to_tile_8_7_1),
		.in_wire_0_2(horizontal_tile_8_8_to_tile_8_7_2),
		.in_wire_0_3(horizontal_tile_8_8_to_tile_8_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(264)
	);

	pe_tile pe_tile_8_8(
		.out_wire_3_0(vertical_tile_8_8_to_tile_7_8_0),
		.out_wire_3_1(vertical_tile_8_8_to_tile_7_8_1),
		.out_wire_3_2(vertical_tile_8_8_to_tile_7_8_2),
		.out_wire_3_3(vertical_tile_8_8_to_tile_7_8_3),
		.in_wire_3_0(vertical_tile_7_8_to_tile_8_8_0),
		.in_wire_3_1(vertical_tile_7_8_to_tile_8_8_1),
		.in_wire_3_2(vertical_tile_7_8_to_tile_8_8_2),
		.in_wire_3_3(vertical_tile_7_8_to_tile_8_8_3),
		.out_wire_1_0(vertical_tile_8_8_to_tile_9_8_0),
		.out_wire_1_1(vertical_tile_8_8_to_tile_9_8_1),
		.out_wire_1_2(vertical_tile_8_8_to_tile_9_8_2),
		.out_wire_1_3(vertical_tile_8_8_to_tile_9_8_3),
		.in_wire_1_0(vertical_tile_9_8_to_tile_8_8_0),
		.in_wire_1_1(vertical_tile_9_8_to_tile_8_8_1),
		.in_wire_1_2(vertical_tile_9_8_to_tile_8_8_2),
		.in_wire_1_3(vertical_tile_9_8_to_tile_8_8_3),
		.out_wire_2_0(horizontal_tile_8_8_to_tile_8_7_0),
		.out_wire_2_1(horizontal_tile_8_8_to_tile_8_7_1),
		.out_wire_2_2(horizontal_tile_8_8_to_tile_8_7_2),
		.out_wire_2_3(horizontal_tile_8_8_to_tile_8_7_3),
		.in_wire_2_0(horizontal_tile_8_7_to_tile_8_8_0),
		.in_wire_2_1(horizontal_tile_8_7_to_tile_8_8_1),
		.in_wire_2_2(horizontal_tile_8_7_to_tile_8_8_2),
		.in_wire_2_3(horizontal_tile_8_7_to_tile_8_8_3),
		.out_wire_0_0(horizontal_tile_8_8_to_tile_8_9_0),
		.out_wire_0_1(horizontal_tile_8_8_to_tile_8_9_1),
		.out_wire_0_2(horizontal_tile_8_8_to_tile_8_9_2),
		.out_wire_0_3(horizontal_tile_8_8_to_tile_8_9_3),
		.in_wire_0_0(horizontal_tile_8_9_to_tile_8_8_0),
		.in_wire_0_1(horizontal_tile_8_9_to_tile_8_8_1),
		.in_wire_0_2(horizontal_tile_8_9_to_tile_8_8_2),
		.in_wire_0_3(horizontal_tile_8_9_to_tile_8_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(265)
	);

	pe_tile pe_tile_8_9(
		.out_wire_3_0(vertical_tile_8_9_to_tile_7_9_0),
		.out_wire_3_1(vertical_tile_8_9_to_tile_7_9_1),
		.out_wire_3_2(vertical_tile_8_9_to_tile_7_9_2),
		.out_wire_3_3(vertical_tile_8_9_to_tile_7_9_3),
		.in_wire_3_0(vertical_tile_7_9_to_tile_8_9_0),
		.in_wire_3_1(vertical_tile_7_9_to_tile_8_9_1),
		.in_wire_3_2(vertical_tile_7_9_to_tile_8_9_2),
		.in_wire_3_3(vertical_tile_7_9_to_tile_8_9_3),
		.out_wire_1_0(vertical_tile_8_9_to_tile_9_9_0),
		.out_wire_1_1(vertical_tile_8_9_to_tile_9_9_1),
		.out_wire_1_2(vertical_tile_8_9_to_tile_9_9_2),
		.out_wire_1_3(vertical_tile_8_9_to_tile_9_9_3),
		.in_wire_1_0(vertical_tile_9_9_to_tile_8_9_0),
		.in_wire_1_1(vertical_tile_9_9_to_tile_8_9_1),
		.in_wire_1_2(vertical_tile_9_9_to_tile_8_9_2),
		.in_wire_1_3(vertical_tile_9_9_to_tile_8_9_3),
		.out_wire_2_0(horizontal_tile_8_9_to_tile_8_8_0),
		.out_wire_2_1(horizontal_tile_8_9_to_tile_8_8_1),
		.out_wire_2_2(horizontal_tile_8_9_to_tile_8_8_2),
		.out_wire_2_3(horizontal_tile_8_9_to_tile_8_8_3),
		.in_wire_2_0(horizontal_tile_8_8_to_tile_8_9_0),
		.in_wire_2_1(horizontal_tile_8_8_to_tile_8_9_1),
		.in_wire_2_2(horizontal_tile_8_8_to_tile_8_9_2),
		.in_wire_2_3(horizontal_tile_8_8_to_tile_8_9_3),
		.out_wire_0_0(horizontal_tile_8_9_to_tile_8_10_0),
		.out_wire_0_1(horizontal_tile_8_9_to_tile_8_10_1),
		.out_wire_0_2(horizontal_tile_8_9_to_tile_8_10_2),
		.out_wire_0_3(horizontal_tile_8_9_to_tile_8_10_3),
		.in_wire_0_0(horizontal_tile_8_10_to_tile_8_9_0),
		.in_wire_0_1(horizontal_tile_8_10_to_tile_8_9_1),
		.in_wire_0_2(horizontal_tile_8_10_to_tile_8_9_2),
		.in_wire_0_3(horizontal_tile_8_10_to_tile_8_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(266)
	);

	pe_tile pe_tile_8_10(
		.out_wire_3_0(vertical_tile_8_10_to_tile_7_10_0),
		.out_wire_3_1(vertical_tile_8_10_to_tile_7_10_1),
		.out_wire_3_2(vertical_tile_8_10_to_tile_7_10_2),
		.out_wire_3_3(vertical_tile_8_10_to_tile_7_10_3),
		.in_wire_3_0(vertical_tile_7_10_to_tile_8_10_0),
		.in_wire_3_1(vertical_tile_7_10_to_tile_8_10_1),
		.in_wire_3_2(vertical_tile_7_10_to_tile_8_10_2),
		.in_wire_3_3(vertical_tile_7_10_to_tile_8_10_3),
		.out_wire_1_0(vertical_tile_8_10_to_tile_9_10_0),
		.out_wire_1_1(vertical_tile_8_10_to_tile_9_10_1),
		.out_wire_1_2(vertical_tile_8_10_to_tile_9_10_2),
		.out_wire_1_3(vertical_tile_8_10_to_tile_9_10_3),
		.in_wire_1_0(vertical_tile_9_10_to_tile_8_10_0),
		.in_wire_1_1(vertical_tile_9_10_to_tile_8_10_1),
		.in_wire_1_2(vertical_tile_9_10_to_tile_8_10_2),
		.in_wire_1_3(vertical_tile_9_10_to_tile_8_10_3),
		.out_wire_2_0(horizontal_tile_8_10_to_tile_8_9_0),
		.out_wire_2_1(horizontal_tile_8_10_to_tile_8_9_1),
		.out_wire_2_2(horizontal_tile_8_10_to_tile_8_9_2),
		.out_wire_2_3(horizontal_tile_8_10_to_tile_8_9_3),
		.in_wire_2_0(horizontal_tile_8_9_to_tile_8_10_0),
		.in_wire_2_1(horizontal_tile_8_9_to_tile_8_10_1),
		.in_wire_2_2(horizontal_tile_8_9_to_tile_8_10_2),
		.in_wire_2_3(horizontal_tile_8_9_to_tile_8_10_3),
		.out_wire_0_0(horizontal_tile_8_10_to_tile_8_11_0),
		.out_wire_0_1(horizontal_tile_8_10_to_tile_8_11_1),
		.out_wire_0_2(horizontal_tile_8_10_to_tile_8_11_2),
		.out_wire_0_3(horizontal_tile_8_10_to_tile_8_11_3),
		.in_wire_0_0(horizontal_tile_8_11_to_tile_8_10_0),
		.in_wire_0_1(horizontal_tile_8_11_to_tile_8_10_1),
		.in_wire_0_2(horizontal_tile_8_11_to_tile_8_10_2),
		.in_wire_0_3(horizontal_tile_8_11_to_tile_8_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(267)
	);

	pe_tile pe_tile_8_11(
		.out_wire_3_0(vertical_tile_8_11_to_tile_7_11_0),
		.out_wire_3_1(vertical_tile_8_11_to_tile_7_11_1),
		.out_wire_3_2(vertical_tile_8_11_to_tile_7_11_2),
		.out_wire_3_3(vertical_tile_8_11_to_tile_7_11_3),
		.in_wire_3_0(vertical_tile_7_11_to_tile_8_11_0),
		.in_wire_3_1(vertical_tile_7_11_to_tile_8_11_1),
		.in_wire_3_2(vertical_tile_7_11_to_tile_8_11_2),
		.in_wire_3_3(vertical_tile_7_11_to_tile_8_11_3),
		.out_wire_1_0(vertical_tile_8_11_to_tile_9_11_0),
		.out_wire_1_1(vertical_tile_8_11_to_tile_9_11_1),
		.out_wire_1_2(vertical_tile_8_11_to_tile_9_11_2),
		.out_wire_1_3(vertical_tile_8_11_to_tile_9_11_3),
		.in_wire_1_0(vertical_tile_9_11_to_tile_8_11_0),
		.in_wire_1_1(vertical_tile_9_11_to_tile_8_11_1),
		.in_wire_1_2(vertical_tile_9_11_to_tile_8_11_2),
		.in_wire_1_3(vertical_tile_9_11_to_tile_8_11_3),
		.out_wire_2_0(horizontal_tile_8_11_to_tile_8_10_0),
		.out_wire_2_1(horizontal_tile_8_11_to_tile_8_10_1),
		.out_wire_2_2(horizontal_tile_8_11_to_tile_8_10_2),
		.out_wire_2_3(horizontal_tile_8_11_to_tile_8_10_3),
		.in_wire_2_0(horizontal_tile_8_10_to_tile_8_11_0),
		.in_wire_2_1(horizontal_tile_8_10_to_tile_8_11_1),
		.in_wire_2_2(horizontal_tile_8_10_to_tile_8_11_2),
		.in_wire_2_3(horizontal_tile_8_10_to_tile_8_11_3),
		.out_wire_0_0(horizontal_tile_8_11_to_tile_8_12_0),
		.out_wire_0_1(horizontal_tile_8_11_to_tile_8_12_1),
		.out_wire_0_2(horizontal_tile_8_11_to_tile_8_12_2),
		.out_wire_0_3(horizontal_tile_8_11_to_tile_8_12_3),
		.in_wire_0_0(horizontal_tile_8_12_to_tile_8_11_0),
		.in_wire_0_1(horizontal_tile_8_12_to_tile_8_11_1),
		.in_wire_0_2(horizontal_tile_8_12_to_tile_8_11_2),
		.in_wire_0_3(horizontal_tile_8_12_to_tile_8_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(268)
	);

	pe_tile pe_tile_8_12(
		.out_wire_3_0(vertical_tile_8_12_to_tile_7_12_0),
		.out_wire_3_1(vertical_tile_8_12_to_tile_7_12_1),
		.out_wire_3_2(vertical_tile_8_12_to_tile_7_12_2),
		.out_wire_3_3(vertical_tile_8_12_to_tile_7_12_3),
		.in_wire_3_0(vertical_tile_7_12_to_tile_8_12_0),
		.in_wire_3_1(vertical_tile_7_12_to_tile_8_12_1),
		.in_wire_3_2(vertical_tile_7_12_to_tile_8_12_2),
		.in_wire_3_3(vertical_tile_7_12_to_tile_8_12_3),
		.out_wire_1_0(vertical_tile_8_12_to_tile_9_12_0),
		.out_wire_1_1(vertical_tile_8_12_to_tile_9_12_1),
		.out_wire_1_2(vertical_tile_8_12_to_tile_9_12_2),
		.out_wire_1_3(vertical_tile_8_12_to_tile_9_12_3),
		.in_wire_1_0(vertical_tile_9_12_to_tile_8_12_0),
		.in_wire_1_1(vertical_tile_9_12_to_tile_8_12_1),
		.in_wire_1_2(vertical_tile_9_12_to_tile_8_12_2),
		.in_wire_1_3(vertical_tile_9_12_to_tile_8_12_3),
		.out_wire_2_0(horizontal_tile_8_12_to_tile_8_11_0),
		.out_wire_2_1(horizontal_tile_8_12_to_tile_8_11_1),
		.out_wire_2_2(horizontal_tile_8_12_to_tile_8_11_2),
		.out_wire_2_3(horizontal_tile_8_12_to_tile_8_11_3),
		.in_wire_2_0(horizontal_tile_8_11_to_tile_8_12_0),
		.in_wire_2_1(horizontal_tile_8_11_to_tile_8_12_1),
		.in_wire_2_2(horizontal_tile_8_11_to_tile_8_12_2),
		.in_wire_2_3(horizontal_tile_8_11_to_tile_8_12_3),
		.out_wire_0_0(horizontal_tile_8_12_to_tile_8_13_0),
		.out_wire_0_1(horizontal_tile_8_12_to_tile_8_13_1),
		.out_wire_0_2(horizontal_tile_8_12_to_tile_8_13_2),
		.out_wire_0_3(horizontal_tile_8_12_to_tile_8_13_3),
		.in_wire_0_0(horizontal_tile_8_13_to_tile_8_12_0),
		.in_wire_0_1(horizontal_tile_8_13_to_tile_8_12_1),
		.in_wire_0_2(horizontal_tile_8_13_to_tile_8_12_2),
		.in_wire_0_3(horizontal_tile_8_13_to_tile_8_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(269)
	);

	pe_tile pe_tile_8_13(
		.out_wire_3_0(vertical_tile_8_13_to_tile_7_13_0),
		.out_wire_3_1(vertical_tile_8_13_to_tile_7_13_1),
		.out_wire_3_2(vertical_tile_8_13_to_tile_7_13_2),
		.out_wire_3_3(vertical_tile_8_13_to_tile_7_13_3),
		.in_wire_3_0(vertical_tile_7_13_to_tile_8_13_0),
		.in_wire_3_1(vertical_tile_7_13_to_tile_8_13_1),
		.in_wire_3_2(vertical_tile_7_13_to_tile_8_13_2),
		.in_wire_3_3(vertical_tile_7_13_to_tile_8_13_3),
		.out_wire_1_0(vertical_tile_8_13_to_tile_9_13_0),
		.out_wire_1_1(vertical_tile_8_13_to_tile_9_13_1),
		.out_wire_1_2(vertical_tile_8_13_to_tile_9_13_2),
		.out_wire_1_3(vertical_tile_8_13_to_tile_9_13_3),
		.in_wire_1_0(vertical_tile_9_13_to_tile_8_13_0),
		.in_wire_1_1(vertical_tile_9_13_to_tile_8_13_1),
		.in_wire_1_2(vertical_tile_9_13_to_tile_8_13_2),
		.in_wire_1_3(vertical_tile_9_13_to_tile_8_13_3),
		.out_wire_2_0(horizontal_tile_8_13_to_tile_8_12_0),
		.out_wire_2_1(horizontal_tile_8_13_to_tile_8_12_1),
		.out_wire_2_2(horizontal_tile_8_13_to_tile_8_12_2),
		.out_wire_2_3(horizontal_tile_8_13_to_tile_8_12_3),
		.in_wire_2_0(horizontal_tile_8_12_to_tile_8_13_0),
		.in_wire_2_1(horizontal_tile_8_12_to_tile_8_13_1),
		.in_wire_2_2(horizontal_tile_8_12_to_tile_8_13_2),
		.in_wire_2_3(horizontal_tile_8_12_to_tile_8_13_3),
		.out_wire_0_0(horizontal_tile_8_13_to_tile_8_14_0),
		.out_wire_0_1(horizontal_tile_8_13_to_tile_8_14_1),
		.out_wire_0_2(horizontal_tile_8_13_to_tile_8_14_2),
		.out_wire_0_3(horizontal_tile_8_13_to_tile_8_14_3),
		.in_wire_0_0(horizontal_tile_8_14_to_tile_8_13_0),
		.in_wire_0_1(horizontal_tile_8_14_to_tile_8_13_1),
		.in_wire_0_2(horizontal_tile_8_14_to_tile_8_13_2),
		.in_wire_0_3(horizontal_tile_8_14_to_tile_8_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(270)
	);

	pe_tile pe_tile_8_14(
		.out_wire_3_0(vertical_tile_8_14_to_tile_7_14_0),
		.out_wire_3_1(vertical_tile_8_14_to_tile_7_14_1),
		.out_wire_3_2(vertical_tile_8_14_to_tile_7_14_2),
		.out_wire_3_3(vertical_tile_8_14_to_tile_7_14_3),
		.in_wire_3_0(vertical_tile_7_14_to_tile_8_14_0),
		.in_wire_3_1(vertical_tile_7_14_to_tile_8_14_1),
		.in_wire_3_2(vertical_tile_7_14_to_tile_8_14_2),
		.in_wire_3_3(vertical_tile_7_14_to_tile_8_14_3),
		.out_wire_1_0(vertical_tile_8_14_to_tile_9_14_0),
		.out_wire_1_1(vertical_tile_8_14_to_tile_9_14_1),
		.out_wire_1_2(vertical_tile_8_14_to_tile_9_14_2),
		.out_wire_1_3(vertical_tile_8_14_to_tile_9_14_3),
		.in_wire_1_0(vertical_tile_9_14_to_tile_8_14_0),
		.in_wire_1_1(vertical_tile_9_14_to_tile_8_14_1),
		.in_wire_1_2(vertical_tile_9_14_to_tile_8_14_2),
		.in_wire_1_3(vertical_tile_9_14_to_tile_8_14_3),
		.out_wire_2_0(horizontal_tile_8_14_to_tile_8_13_0),
		.out_wire_2_1(horizontal_tile_8_14_to_tile_8_13_1),
		.out_wire_2_2(horizontal_tile_8_14_to_tile_8_13_2),
		.out_wire_2_3(horizontal_tile_8_14_to_tile_8_13_3),
		.in_wire_2_0(horizontal_tile_8_13_to_tile_8_14_0),
		.in_wire_2_1(horizontal_tile_8_13_to_tile_8_14_1),
		.in_wire_2_2(horizontal_tile_8_13_to_tile_8_14_2),
		.in_wire_2_3(horizontal_tile_8_13_to_tile_8_14_3),
		.out_wire_0_0(horizontal_tile_8_14_to_tile_8_15_0),
		.out_wire_0_1(horizontal_tile_8_14_to_tile_8_15_1),
		.out_wire_0_2(horizontal_tile_8_14_to_tile_8_15_2),
		.out_wire_0_3(horizontal_tile_8_14_to_tile_8_15_3),
		.in_wire_0_0(horizontal_tile_8_15_to_tile_8_14_0),
		.in_wire_0_1(horizontal_tile_8_15_to_tile_8_14_1),
		.in_wire_0_2(horizontal_tile_8_15_to_tile_8_14_2),
		.in_wire_0_3(horizontal_tile_8_15_to_tile_8_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(271)
	);

	pe_tile pe_tile_8_15(
		.out_wire_3_0(vertical_tile_8_15_to_tile_7_15_0),
		.out_wire_3_1(vertical_tile_8_15_to_tile_7_15_1),
		.out_wire_3_2(vertical_tile_8_15_to_tile_7_15_2),
		.out_wire_3_3(vertical_tile_8_15_to_tile_7_15_3),
		.in_wire_3_0(vertical_tile_7_15_to_tile_8_15_0),
		.in_wire_3_1(vertical_tile_7_15_to_tile_8_15_1),
		.in_wire_3_2(vertical_tile_7_15_to_tile_8_15_2),
		.in_wire_3_3(vertical_tile_7_15_to_tile_8_15_3),
		.out_wire_1_0(vertical_tile_8_15_to_tile_9_15_0),
		.out_wire_1_1(vertical_tile_8_15_to_tile_9_15_1),
		.out_wire_1_2(vertical_tile_8_15_to_tile_9_15_2),
		.out_wire_1_3(vertical_tile_8_15_to_tile_9_15_3),
		.in_wire_1_0(vertical_tile_9_15_to_tile_8_15_0),
		.in_wire_1_1(vertical_tile_9_15_to_tile_8_15_1),
		.in_wire_1_2(vertical_tile_9_15_to_tile_8_15_2),
		.in_wire_1_3(vertical_tile_9_15_to_tile_8_15_3),
		.out_wire_2_0(horizontal_tile_8_15_to_tile_8_14_0),
		.out_wire_2_1(horizontal_tile_8_15_to_tile_8_14_1),
		.out_wire_2_2(horizontal_tile_8_15_to_tile_8_14_2),
		.out_wire_2_3(horizontal_tile_8_15_to_tile_8_14_3),
		.in_wire_2_0(horizontal_tile_8_14_to_tile_8_15_0),
		.in_wire_2_1(horizontal_tile_8_14_to_tile_8_15_1),
		.in_wire_2_2(horizontal_tile_8_14_to_tile_8_15_2),
		.in_wire_2_3(horizontal_tile_8_14_to_tile_8_15_3),
		.out_wire_0_0(horizontal_tile_8_15_to_tile_8_16_0),
		.out_wire_0_1(horizontal_tile_8_15_to_tile_8_16_1),
		.out_wire_0_2(horizontal_tile_8_15_to_tile_8_16_2),
		.out_wire_0_3(horizontal_tile_8_15_to_tile_8_16_3),
		.in_wire_0_0(horizontal_tile_8_16_to_tile_8_15_0),
		.in_wire_0_1(horizontal_tile_8_16_to_tile_8_15_1),
		.in_wire_0_2(horizontal_tile_8_16_to_tile_8_15_2),
		.in_wire_0_3(horizontal_tile_8_16_to_tile_8_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(272)
	);

	pe_tile pe_tile_8_16(
		.out_wire_3_0(vertical_tile_8_16_to_tile_7_16_0),
		.out_wire_3_1(vertical_tile_8_16_to_tile_7_16_1),
		.out_wire_3_2(vertical_tile_8_16_to_tile_7_16_2),
		.out_wire_3_3(vertical_tile_8_16_to_tile_7_16_3),
		.in_wire_3_0(vertical_tile_7_16_to_tile_8_16_0),
		.in_wire_3_1(vertical_tile_7_16_to_tile_8_16_1),
		.in_wire_3_2(vertical_tile_7_16_to_tile_8_16_2),
		.in_wire_3_3(vertical_tile_7_16_to_tile_8_16_3),
		.out_wire_1_0(vertical_tile_8_16_to_tile_9_16_0),
		.out_wire_1_1(vertical_tile_8_16_to_tile_9_16_1),
		.out_wire_1_2(vertical_tile_8_16_to_tile_9_16_2),
		.out_wire_1_3(vertical_tile_8_16_to_tile_9_16_3),
		.in_wire_1_0(vertical_tile_9_16_to_tile_8_16_0),
		.in_wire_1_1(vertical_tile_9_16_to_tile_8_16_1),
		.in_wire_1_2(vertical_tile_9_16_to_tile_8_16_2),
		.in_wire_1_3(vertical_tile_9_16_to_tile_8_16_3),
		.out_wire_2_0(horizontal_tile_8_16_to_tile_8_15_0),
		.out_wire_2_1(horizontal_tile_8_16_to_tile_8_15_1),
		.out_wire_2_2(horizontal_tile_8_16_to_tile_8_15_2),
		.out_wire_2_3(horizontal_tile_8_16_to_tile_8_15_3),
		.in_wire_2_0(horizontal_tile_8_15_to_tile_8_16_0),
		.in_wire_2_1(horizontal_tile_8_15_to_tile_8_16_1),
		.in_wire_2_2(horizontal_tile_8_15_to_tile_8_16_2),
		.in_wire_2_3(horizontal_tile_8_15_to_tile_8_16_3),
		.out_wire_0_0(horizontal_tile_8_16_to_tile_8_17_0),
		.out_wire_0_1(horizontal_tile_8_16_to_tile_8_17_1),
		.out_wire_0_2(horizontal_tile_8_16_to_tile_8_17_2),
		.out_wire_0_3(horizontal_tile_8_16_to_tile_8_17_3),
		.in_wire_0_0(horizontal_tile_8_17_to_tile_8_16_0),
		.in_wire_0_1(horizontal_tile_8_17_to_tile_8_16_1),
		.in_wire_0_2(horizontal_tile_8_17_to_tile_8_16_2),
		.in_wire_0_3(horizontal_tile_8_17_to_tile_8_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(273)
	);

	pe_tile pe_tile_8_17(
		.out_wire_3_0(vertical_tile_8_17_to_tile_7_17_0),
		.out_wire_3_1(vertical_tile_8_17_to_tile_7_17_1),
		.out_wire_3_2(vertical_tile_8_17_to_tile_7_17_2),
		.out_wire_3_3(vertical_tile_8_17_to_tile_7_17_3),
		.in_wire_3_0(vertical_tile_7_17_to_tile_8_17_0),
		.in_wire_3_1(vertical_tile_7_17_to_tile_8_17_1),
		.in_wire_3_2(vertical_tile_7_17_to_tile_8_17_2),
		.in_wire_3_3(vertical_tile_7_17_to_tile_8_17_3),
		.out_wire_1_0(vertical_tile_8_17_to_tile_9_17_0),
		.out_wire_1_1(vertical_tile_8_17_to_tile_9_17_1),
		.out_wire_1_2(vertical_tile_8_17_to_tile_9_17_2),
		.out_wire_1_3(vertical_tile_8_17_to_tile_9_17_3),
		.in_wire_1_0(vertical_tile_9_17_to_tile_8_17_0),
		.in_wire_1_1(vertical_tile_9_17_to_tile_8_17_1),
		.in_wire_1_2(vertical_tile_9_17_to_tile_8_17_2),
		.in_wire_1_3(vertical_tile_9_17_to_tile_8_17_3),
		.out_wire_2_0(horizontal_tile_8_17_to_tile_8_16_0),
		.out_wire_2_1(horizontal_tile_8_17_to_tile_8_16_1),
		.out_wire_2_2(horizontal_tile_8_17_to_tile_8_16_2),
		.out_wire_2_3(horizontal_tile_8_17_to_tile_8_16_3),
		.in_wire_2_0(horizontal_tile_8_16_to_tile_8_17_0),
		.in_wire_2_1(horizontal_tile_8_16_to_tile_8_17_1),
		.in_wire_2_2(horizontal_tile_8_16_to_tile_8_17_2),
		.in_wire_2_3(horizontal_tile_8_16_to_tile_8_17_3),
		.out_wire_0_0(horizontal_tile_8_17_to_tile_8_18_0),
		.out_wire_0_1(horizontal_tile_8_17_to_tile_8_18_1),
		.out_wire_0_2(horizontal_tile_8_17_to_tile_8_18_2),
		.out_wire_0_3(horizontal_tile_8_17_to_tile_8_18_3),
		.in_wire_0_0(horizontal_tile_8_18_to_tile_8_17_0),
		.in_wire_0_1(horizontal_tile_8_18_to_tile_8_17_1),
		.in_wire_0_2(horizontal_tile_8_18_to_tile_8_17_2),
		.in_wire_0_3(horizontal_tile_8_18_to_tile_8_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(274)
	);

	pe_tile pe_tile_8_18(
		.out_wire_3_0(vertical_tile_8_18_to_tile_7_18_0),
		.out_wire_3_1(vertical_tile_8_18_to_tile_7_18_1),
		.out_wire_3_2(vertical_tile_8_18_to_tile_7_18_2),
		.out_wire_3_3(vertical_tile_8_18_to_tile_7_18_3),
		.in_wire_3_0(vertical_tile_7_18_to_tile_8_18_0),
		.in_wire_3_1(vertical_tile_7_18_to_tile_8_18_1),
		.in_wire_3_2(vertical_tile_7_18_to_tile_8_18_2),
		.in_wire_3_3(vertical_tile_7_18_to_tile_8_18_3),
		.out_wire_1_0(vertical_tile_8_18_to_tile_9_18_0),
		.out_wire_1_1(vertical_tile_8_18_to_tile_9_18_1),
		.out_wire_1_2(vertical_tile_8_18_to_tile_9_18_2),
		.out_wire_1_3(vertical_tile_8_18_to_tile_9_18_3),
		.in_wire_1_0(vertical_tile_9_18_to_tile_8_18_0),
		.in_wire_1_1(vertical_tile_9_18_to_tile_8_18_1),
		.in_wire_1_2(vertical_tile_9_18_to_tile_8_18_2),
		.in_wire_1_3(vertical_tile_9_18_to_tile_8_18_3),
		.out_wire_2_0(horizontal_tile_8_18_to_tile_8_17_0),
		.out_wire_2_1(horizontal_tile_8_18_to_tile_8_17_1),
		.out_wire_2_2(horizontal_tile_8_18_to_tile_8_17_2),
		.out_wire_2_3(horizontal_tile_8_18_to_tile_8_17_3),
		.in_wire_2_0(horizontal_tile_8_17_to_tile_8_18_0),
		.in_wire_2_1(horizontal_tile_8_17_to_tile_8_18_1),
		.in_wire_2_2(horizontal_tile_8_17_to_tile_8_18_2),
		.in_wire_2_3(horizontal_tile_8_17_to_tile_8_18_3),
		.out_wire_0_0(horizontal_tile_8_18_to_tile_8_19_0),
		.out_wire_0_1(horizontal_tile_8_18_to_tile_8_19_1),
		.out_wire_0_2(horizontal_tile_8_18_to_tile_8_19_2),
		.out_wire_0_3(horizontal_tile_8_18_to_tile_8_19_3),
		.in_wire_0_0(horizontal_tile_8_19_to_tile_8_18_0),
		.in_wire_0_1(horizontal_tile_8_19_to_tile_8_18_1),
		.in_wire_0_2(horizontal_tile_8_19_to_tile_8_18_2),
		.in_wire_0_3(horizontal_tile_8_19_to_tile_8_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(275)
	);

	pe_tile pe_tile_8_19(
		.out_wire_3_0(vertical_tile_8_19_to_tile_7_19_0),
		.out_wire_3_1(vertical_tile_8_19_to_tile_7_19_1),
		.out_wire_3_2(vertical_tile_8_19_to_tile_7_19_2),
		.out_wire_3_3(vertical_tile_8_19_to_tile_7_19_3),
		.in_wire_3_0(vertical_tile_7_19_to_tile_8_19_0),
		.in_wire_3_1(vertical_tile_7_19_to_tile_8_19_1),
		.in_wire_3_2(vertical_tile_7_19_to_tile_8_19_2),
		.in_wire_3_3(vertical_tile_7_19_to_tile_8_19_3),
		.out_wire_1_0(vertical_tile_8_19_to_tile_9_19_0),
		.out_wire_1_1(vertical_tile_8_19_to_tile_9_19_1),
		.out_wire_1_2(vertical_tile_8_19_to_tile_9_19_2),
		.out_wire_1_3(vertical_tile_8_19_to_tile_9_19_3),
		.in_wire_1_0(vertical_tile_9_19_to_tile_8_19_0),
		.in_wire_1_1(vertical_tile_9_19_to_tile_8_19_1),
		.in_wire_1_2(vertical_tile_9_19_to_tile_8_19_2),
		.in_wire_1_3(vertical_tile_9_19_to_tile_8_19_3),
		.out_wire_2_0(horizontal_tile_8_19_to_tile_8_18_0),
		.out_wire_2_1(horizontal_tile_8_19_to_tile_8_18_1),
		.out_wire_2_2(horizontal_tile_8_19_to_tile_8_18_2),
		.out_wire_2_3(horizontal_tile_8_19_to_tile_8_18_3),
		.in_wire_2_0(horizontal_tile_8_18_to_tile_8_19_0),
		.in_wire_2_1(horizontal_tile_8_18_to_tile_8_19_1),
		.in_wire_2_2(horizontal_tile_8_18_to_tile_8_19_2),
		.in_wire_2_3(horizontal_tile_8_18_to_tile_8_19_3),
		.out_wire_0_0(horizontal_tile_8_19_to_tile_8_20_0),
		.out_wire_0_1(horizontal_tile_8_19_to_tile_8_20_1),
		.out_wire_0_2(horizontal_tile_8_19_to_tile_8_20_2),
		.out_wire_0_3(horizontal_tile_8_19_to_tile_8_20_3),
		.in_wire_0_0(horizontal_tile_8_20_to_tile_8_19_0),
		.in_wire_0_1(horizontal_tile_8_20_to_tile_8_19_1),
		.in_wire_0_2(horizontal_tile_8_20_to_tile_8_19_2),
		.in_wire_0_3(horizontal_tile_8_20_to_tile_8_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(276)
	);

	pe_tile pe_tile_8_20(
		.out_wire_3_0(vertical_tile_8_20_to_tile_7_20_0),
		.out_wire_3_1(vertical_tile_8_20_to_tile_7_20_1),
		.out_wire_3_2(vertical_tile_8_20_to_tile_7_20_2),
		.out_wire_3_3(vertical_tile_8_20_to_tile_7_20_3),
		.in_wire_3_0(vertical_tile_7_20_to_tile_8_20_0),
		.in_wire_3_1(vertical_tile_7_20_to_tile_8_20_1),
		.in_wire_3_2(vertical_tile_7_20_to_tile_8_20_2),
		.in_wire_3_3(vertical_tile_7_20_to_tile_8_20_3),
		.out_wire_1_0(vertical_tile_8_20_to_tile_9_20_0),
		.out_wire_1_1(vertical_tile_8_20_to_tile_9_20_1),
		.out_wire_1_2(vertical_tile_8_20_to_tile_9_20_2),
		.out_wire_1_3(vertical_tile_8_20_to_tile_9_20_3),
		.in_wire_1_0(vertical_tile_9_20_to_tile_8_20_0),
		.in_wire_1_1(vertical_tile_9_20_to_tile_8_20_1),
		.in_wire_1_2(vertical_tile_9_20_to_tile_8_20_2),
		.in_wire_1_3(vertical_tile_9_20_to_tile_8_20_3),
		.out_wire_2_0(horizontal_tile_8_20_to_tile_8_19_0),
		.out_wire_2_1(horizontal_tile_8_20_to_tile_8_19_1),
		.out_wire_2_2(horizontal_tile_8_20_to_tile_8_19_2),
		.out_wire_2_3(horizontal_tile_8_20_to_tile_8_19_3),
		.in_wire_2_0(horizontal_tile_8_19_to_tile_8_20_0),
		.in_wire_2_1(horizontal_tile_8_19_to_tile_8_20_1),
		.in_wire_2_2(horizontal_tile_8_19_to_tile_8_20_2),
		.in_wire_2_3(horizontal_tile_8_19_to_tile_8_20_3),
		.out_wire_0_0(horizontal_tile_8_20_to_tile_8_21_0),
		.out_wire_0_1(horizontal_tile_8_20_to_tile_8_21_1),
		.out_wire_0_2(horizontal_tile_8_20_to_tile_8_21_2),
		.out_wire_0_3(horizontal_tile_8_20_to_tile_8_21_3),
		.in_wire_0_0(horizontal_tile_8_21_to_tile_8_20_0),
		.in_wire_0_1(horizontal_tile_8_21_to_tile_8_20_1),
		.in_wire_0_2(horizontal_tile_8_21_to_tile_8_20_2),
		.in_wire_0_3(horizontal_tile_8_21_to_tile_8_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(277)
	);

	pe_tile pe_tile_8_21(
		.out_wire_3_0(vertical_tile_8_21_to_tile_7_21_0),
		.out_wire_3_1(vertical_tile_8_21_to_tile_7_21_1),
		.out_wire_3_2(vertical_tile_8_21_to_tile_7_21_2),
		.out_wire_3_3(vertical_tile_8_21_to_tile_7_21_3),
		.in_wire_3_0(vertical_tile_7_21_to_tile_8_21_0),
		.in_wire_3_1(vertical_tile_7_21_to_tile_8_21_1),
		.in_wire_3_2(vertical_tile_7_21_to_tile_8_21_2),
		.in_wire_3_3(vertical_tile_7_21_to_tile_8_21_3),
		.out_wire_1_0(vertical_tile_8_21_to_tile_9_21_0),
		.out_wire_1_1(vertical_tile_8_21_to_tile_9_21_1),
		.out_wire_1_2(vertical_tile_8_21_to_tile_9_21_2),
		.out_wire_1_3(vertical_tile_8_21_to_tile_9_21_3),
		.in_wire_1_0(vertical_tile_9_21_to_tile_8_21_0),
		.in_wire_1_1(vertical_tile_9_21_to_tile_8_21_1),
		.in_wire_1_2(vertical_tile_9_21_to_tile_8_21_2),
		.in_wire_1_3(vertical_tile_9_21_to_tile_8_21_3),
		.out_wire_2_0(horizontal_tile_8_21_to_tile_8_20_0),
		.out_wire_2_1(horizontal_tile_8_21_to_tile_8_20_1),
		.out_wire_2_2(horizontal_tile_8_21_to_tile_8_20_2),
		.out_wire_2_3(horizontal_tile_8_21_to_tile_8_20_3),
		.in_wire_2_0(horizontal_tile_8_20_to_tile_8_21_0),
		.in_wire_2_1(horizontal_tile_8_20_to_tile_8_21_1),
		.in_wire_2_2(horizontal_tile_8_20_to_tile_8_21_2),
		.in_wire_2_3(horizontal_tile_8_20_to_tile_8_21_3),
		.out_wire_0_0(horizontal_tile_8_21_to_tile_8_22_0),
		.out_wire_0_1(horizontal_tile_8_21_to_tile_8_22_1),
		.out_wire_0_2(horizontal_tile_8_21_to_tile_8_22_2),
		.out_wire_0_3(horizontal_tile_8_21_to_tile_8_22_3),
		.in_wire_0_0(horizontal_tile_8_22_to_tile_8_21_0),
		.in_wire_0_1(horizontal_tile_8_22_to_tile_8_21_1),
		.in_wire_0_2(horizontal_tile_8_22_to_tile_8_21_2),
		.in_wire_0_3(horizontal_tile_8_22_to_tile_8_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(278)
	);

	pe_tile pe_tile_8_22(
		.out_wire_3_0(vertical_tile_8_22_to_tile_7_22_0),
		.out_wire_3_1(vertical_tile_8_22_to_tile_7_22_1),
		.out_wire_3_2(vertical_tile_8_22_to_tile_7_22_2),
		.out_wire_3_3(vertical_tile_8_22_to_tile_7_22_3),
		.in_wire_3_0(vertical_tile_7_22_to_tile_8_22_0),
		.in_wire_3_1(vertical_tile_7_22_to_tile_8_22_1),
		.in_wire_3_2(vertical_tile_7_22_to_tile_8_22_2),
		.in_wire_3_3(vertical_tile_7_22_to_tile_8_22_3),
		.out_wire_1_0(vertical_tile_8_22_to_tile_9_22_0),
		.out_wire_1_1(vertical_tile_8_22_to_tile_9_22_1),
		.out_wire_1_2(vertical_tile_8_22_to_tile_9_22_2),
		.out_wire_1_3(vertical_tile_8_22_to_tile_9_22_3),
		.in_wire_1_0(vertical_tile_9_22_to_tile_8_22_0),
		.in_wire_1_1(vertical_tile_9_22_to_tile_8_22_1),
		.in_wire_1_2(vertical_tile_9_22_to_tile_8_22_2),
		.in_wire_1_3(vertical_tile_9_22_to_tile_8_22_3),
		.out_wire_2_0(horizontal_tile_8_22_to_tile_8_21_0),
		.out_wire_2_1(horizontal_tile_8_22_to_tile_8_21_1),
		.out_wire_2_2(horizontal_tile_8_22_to_tile_8_21_2),
		.out_wire_2_3(horizontal_tile_8_22_to_tile_8_21_3),
		.in_wire_2_0(horizontal_tile_8_21_to_tile_8_22_0),
		.in_wire_2_1(horizontal_tile_8_21_to_tile_8_22_1),
		.in_wire_2_2(horizontal_tile_8_21_to_tile_8_22_2),
		.in_wire_2_3(horizontal_tile_8_21_to_tile_8_22_3),
		.out_wire_0_0(horizontal_tile_8_22_to_tile_8_23_0),
		.out_wire_0_1(horizontal_tile_8_22_to_tile_8_23_1),
		.out_wire_0_2(horizontal_tile_8_22_to_tile_8_23_2),
		.out_wire_0_3(horizontal_tile_8_22_to_tile_8_23_3),
		.in_wire_0_0(horizontal_tile_8_23_to_tile_8_22_0),
		.in_wire_0_1(horizontal_tile_8_23_to_tile_8_22_1),
		.in_wire_0_2(horizontal_tile_8_23_to_tile_8_22_2),
		.in_wire_0_3(horizontal_tile_8_23_to_tile_8_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(279)
	);

	pe_tile pe_tile_8_23(
		.out_wire_3_0(vertical_tile_8_23_to_tile_7_23_0),
		.out_wire_3_1(vertical_tile_8_23_to_tile_7_23_1),
		.out_wire_3_2(vertical_tile_8_23_to_tile_7_23_2),
		.out_wire_3_3(vertical_tile_8_23_to_tile_7_23_3),
		.in_wire_3_0(vertical_tile_7_23_to_tile_8_23_0),
		.in_wire_3_1(vertical_tile_7_23_to_tile_8_23_1),
		.in_wire_3_2(vertical_tile_7_23_to_tile_8_23_2),
		.in_wire_3_3(vertical_tile_7_23_to_tile_8_23_3),
		.out_wire_1_0(vertical_tile_8_23_to_tile_9_23_0),
		.out_wire_1_1(vertical_tile_8_23_to_tile_9_23_1),
		.out_wire_1_2(vertical_tile_8_23_to_tile_9_23_2),
		.out_wire_1_3(vertical_tile_8_23_to_tile_9_23_3),
		.in_wire_1_0(vertical_tile_9_23_to_tile_8_23_0),
		.in_wire_1_1(vertical_tile_9_23_to_tile_8_23_1),
		.in_wire_1_2(vertical_tile_9_23_to_tile_8_23_2),
		.in_wire_1_3(vertical_tile_9_23_to_tile_8_23_3),
		.out_wire_2_0(horizontal_tile_8_23_to_tile_8_22_0),
		.out_wire_2_1(horizontal_tile_8_23_to_tile_8_22_1),
		.out_wire_2_2(horizontal_tile_8_23_to_tile_8_22_2),
		.out_wire_2_3(horizontal_tile_8_23_to_tile_8_22_3),
		.in_wire_2_0(horizontal_tile_8_22_to_tile_8_23_0),
		.in_wire_2_1(horizontal_tile_8_22_to_tile_8_23_1),
		.in_wire_2_2(horizontal_tile_8_22_to_tile_8_23_2),
		.in_wire_2_3(horizontal_tile_8_22_to_tile_8_23_3),
		.out_wire_0_0(horizontal_tile_8_23_to_tile_8_24_0),
		.out_wire_0_1(horizontal_tile_8_23_to_tile_8_24_1),
		.out_wire_0_2(horizontal_tile_8_23_to_tile_8_24_2),
		.out_wire_0_3(horizontal_tile_8_23_to_tile_8_24_3),
		.in_wire_0_0(horizontal_tile_8_24_to_tile_8_23_0),
		.in_wire_0_1(horizontal_tile_8_24_to_tile_8_23_1),
		.in_wire_0_2(horizontal_tile_8_24_to_tile_8_23_2),
		.in_wire_0_3(horizontal_tile_8_24_to_tile_8_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(280)
	);

	pe_tile pe_tile_8_24(
		.out_wire_3_0(vertical_tile_8_24_to_tile_7_24_0),
		.out_wire_3_1(vertical_tile_8_24_to_tile_7_24_1),
		.out_wire_3_2(vertical_tile_8_24_to_tile_7_24_2),
		.out_wire_3_3(vertical_tile_8_24_to_tile_7_24_3),
		.in_wire_3_0(vertical_tile_7_24_to_tile_8_24_0),
		.in_wire_3_1(vertical_tile_7_24_to_tile_8_24_1),
		.in_wire_3_2(vertical_tile_7_24_to_tile_8_24_2),
		.in_wire_3_3(vertical_tile_7_24_to_tile_8_24_3),
		.out_wire_1_0(vertical_tile_8_24_to_tile_9_24_0),
		.out_wire_1_1(vertical_tile_8_24_to_tile_9_24_1),
		.out_wire_1_2(vertical_tile_8_24_to_tile_9_24_2),
		.out_wire_1_3(vertical_tile_8_24_to_tile_9_24_3),
		.in_wire_1_0(vertical_tile_9_24_to_tile_8_24_0),
		.in_wire_1_1(vertical_tile_9_24_to_tile_8_24_1),
		.in_wire_1_2(vertical_tile_9_24_to_tile_8_24_2),
		.in_wire_1_3(vertical_tile_9_24_to_tile_8_24_3),
		.out_wire_2_0(horizontal_tile_8_24_to_tile_8_23_0),
		.out_wire_2_1(horizontal_tile_8_24_to_tile_8_23_1),
		.out_wire_2_2(horizontal_tile_8_24_to_tile_8_23_2),
		.out_wire_2_3(horizontal_tile_8_24_to_tile_8_23_3),
		.in_wire_2_0(horizontal_tile_8_23_to_tile_8_24_0),
		.in_wire_2_1(horizontal_tile_8_23_to_tile_8_24_1),
		.in_wire_2_2(horizontal_tile_8_23_to_tile_8_24_2),
		.in_wire_2_3(horizontal_tile_8_23_to_tile_8_24_3),
		.out_wire_0_0(horizontal_tile_8_24_to_tile_8_25_0),
		.out_wire_0_1(horizontal_tile_8_24_to_tile_8_25_1),
		.out_wire_0_2(horizontal_tile_8_24_to_tile_8_25_2),
		.out_wire_0_3(horizontal_tile_8_24_to_tile_8_25_3),
		.in_wire_0_0(horizontal_tile_8_25_to_tile_8_24_0),
		.in_wire_0_1(horizontal_tile_8_25_to_tile_8_24_1),
		.in_wire_0_2(horizontal_tile_8_25_to_tile_8_24_2),
		.in_wire_0_3(horizontal_tile_8_25_to_tile_8_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(281)
	);

	pe_tile pe_tile_8_25(
		.out_wire_3_0(vertical_tile_8_25_to_tile_7_25_0),
		.out_wire_3_1(vertical_tile_8_25_to_tile_7_25_1),
		.out_wire_3_2(vertical_tile_8_25_to_tile_7_25_2),
		.out_wire_3_3(vertical_tile_8_25_to_tile_7_25_3),
		.in_wire_3_0(vertical_tile_7_25_to_tile_8_25_0),
		.in_wire_3_1(vertical_tile_7_25_to_tile_8_25_1),
		.in_wire_3_2(vertical_tile_7_25_to_tile_8_25_2),
		.in_wire_3_3(vertical_tile_7_25_to_tile_8_25_3),
		.out_wire_1_0(vertical_tile_8_25_to_tile_9_25_0),
		.out_wire_1_1(vertical_tile_8_25_to_tile_9_25_1),
		.out_wire_1_2(vertical_tile_8_25_to_tile_9_25_2),
		.out_wire_1_3(vertical_tile_8_25_to_tile_9_25_3),
		.in_wire_1_0(vertical_tile_9_25_to_tile_8_25_0),
		.in_wire_1_1(vertical_tile_9_25_to_tile_8_25_1),
		.in_wire_1_2(vertical_tile_9_25_to_tile_8_25_2),
		.in_wire_1_3(vertical_tile_9_25_to_tile_8_25_3),
		.out_wire_2_0(horizontal_tile_8_25_to_tile_8_24_0),
		.out_wire_2_1(horizontal_tile_8_25_to_tile_8_24_1),
		.out_wire_2_2(horizontal_tile_8_25_to_tile_8_24_2),
		.out_wire_2_3(horizontal_tile_8_25_to_tile_8_24_3),
		.in_wire_2_0(horizontal_tile_8_24_to_tile_8_25_0),
		.in_wire_2_1(horizontal_tile_8_24_to_tile_8_25_1),
		.in_wire_2_2(horizontal_tile_8_24_to_tile_8_25_2),
		.in_wire_2_3(horizontal_tile_8_24_to_tile_8_25_3),
		.out_wire_0_0(horizontal_tile_8_25_to_tile_8_26_0),
		.out_wire_0_1(horizontal_tile_8_25_to_tile_8_26_1),
		.out_wire_0_2(horizontal_tile_8_25_to_tile_8_26_2),
		.out_wire_0_3(horizontal_tile_8_25_to_tile_8_26_3),
		.in_wire_0_0(horizontal_tile_8_26_to_tile_8_25_0),
		.in_wire_0_1(horizontal_tile_8_26_to_tile_8_25_1),
		.in_wire_0_2(horizontal_tile_8_26_to_tile_8_25_2),
		.in_wire_0_3(horizontal_tile_8_26_to_tile_8_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(282)
	);

	pe_tile pe_tile_8_26(
		.out_wire_3_0(vertical_tile_8_26_to_tile_7_26_0),
		.out_wire_3_1(vertical_tile_8_26_to_tile_7_26_1),
		.out_wire_3_2(vertical_tile_8_26_to_tile_7_26_2),
		.out_wire_3_3(vertical_tile_8_26_to_tile_7_26_3),
		.in_wire_3_0(vertical_tile_7_26_to_tile_8_26_0),
		.in_wire_3_1(vertical_tile_7_26_to_tile_8_26_1),
		.in_wire_3_2(vertical_tile_7_26_to_tile_8_26_2),
		.in_wire_3_3(vertical_tile_7_26_to_tile_8_26_3),
		.out_wire_1_0(vertical_tile_8_26_to_tile_9_26_0),
		.out_wire_1_1(vertical_tile_8_26_to_tile_9_26_1),
		.out_wire_1_2(vertical_tile_8_26_to_tile_9_26_2),
		.out_wire_1_3(vertical_tile_8_26_to_tile_9_26_3),
		.in_wire_1_0(vertical_tile_9_26_to_tile_8_26_0),
		.in_wire_1_1(vertical_tile_9_26_to_tile_8_26_1),
		.in_wire_1_2(vertical_tile_9_26_to_tile_8_26_2),
		.in_wire_1_3(vertical_tile_9_26_to_tile_8_26_3),
		.out_wire_2_0(horizontal_tile_8_26_to_tile_8_25_0),
		.out_wire_2_1(horizontal_tile_8_26_to_tile_8_25_1),
		.out_wire_2_2(horizontal_tile_8_26_to_tile_8_25_2),
		.out_wire_2_3(horizontal_tile_8_26_to_tile_8_25_3),
		.in_wire_2_0(horizontal_tile_8_25_to_tile_8_26_0),
		.in_wire_2_1(horizontal_tile_8_25_to_tile_8_26_1),
		.in_wire_2_2(horizontal_tile_8_25_to_tile_8_26_2),
		.in_wire_2_3(horizontal_tile_8_25_to_tile_8_26_3),
		.out_wire_0_0(horizontal_tile_8_26_to_tile_8_27_0),
		.out_wire_0_1(horizontal_tile_8_26_to_tile_8_27_1),
		.out_wire_0_2(horizontal_tile_8_26_to_tile_8_27_2),
		.out_wire_0_3(horizontal_tile_8_26_to_tile_8_27_3),
		.in_wire_0_0(horizontal_tile_8_27_to_tile_8_26_0),
		.in_wire_0_1(horizontal_tile_8_27_to_tile_8_26_1),
		.in_wire_0_2(horizontal_tile_8_27_to_tile_8_26_2),
		.in_wire_0_3(horizontal_tile_8_27_to_tile_8_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(283)
	);

	pe_tile pe_tile_8_27(
		.out_wire_3_0(vertical_tile_8_27_to_tile_7_27_0),
		.out_wire_3_1(vertical_tile_8_27_to_tile_7_27_1),
		.out_wire_3_2(vertical_tile_8_27_to_tile_7_27_2),
		.out_wire_3_3(vertical_tile_8_27_to_tile_7_27_3),
		.in_wire_3_0(vertical_tile_7_27_to_tile_8_27_0),
		.in_wire_3_1(vertical_tile_7_27_to_tile_8_27_1),
		.in_wire_3_2(vertical_tile_7_27_to_tile_8_27_2),
		.in_wire_3_3(vertical_tile_7_27_to_tile_8_27_3),
		.out_wire_1_0(vertical_tile_8_27_to_tile_9_27_0),
		.out_wire_1_1(vertical_tile_8_27_to_tile_9_27_1),
		.out_wire_1_2(vertical_tile_8_27_to_tile_9_27_2),
		.out_wire_1_3(vertical_tile_8_27_to_tile_9_27_3),
		.in_wire_1_0(vertical_tile_9_27_to_tile_8_27_0),
		.in_wire_1_1(vertical_tile_9_27_to_tile_8_27_1),
		.in_wire_1_2(vertical_tile_9_27_to_tile_8_27_2),
		.in_wire_1_3(vertical_tile_9_27_to_tile_8_27_3),
		.out_wire_2_0(horizontal_tile_8_27_to_tile_8_26_0),
		.out_wire_2_1(horizontal_tile_8_27_to_tile_8_26_1),
		.out_wire_2_2(horizontal_tile_8_27_to_tile_8_26_2),
		.out_wire_2_3(horizontal_tile_8_27_to_tile_8_26_3),
		.in_wire_2_0(horizontal_tile_8_26_to_tile_8_27_0),
		.in_wire_2_1(horizontal_tile_8_26_to_tile_8_27_1),
		.in_wire_2_2(horizontal_tile_8_26_to_tile_8_27_2),
		.in_wire_2_3(horizontal_tile_8_26_to_tile_8_27_3),
		.out_wire_0_0(horizontal_tile_8_27_to_tile_8_28_0),
		.out_wire_0_1(horizontal_tile_8_27_to_tile_8_28_1),
		.out_wire_0_2(horizontal_tile_8_27_to_tile_8_28_2),
		.out_wire_0_3(horizontal_tile_8_27_to_tile_8_28_3),
		.in_wire_0_0(horizontal_tile_8_28_to_tile_8_27_0),
		.in_wire_0_1(horizontal_tile_8_28_to_tile_8_27_1),
		.in_wire_0_2(horizontal_tile_8_28_to_tile_8_27_2),
		.in_wire_0_3(horizontal_tile_8_28_to_tile_8_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(284)
	);

	pe_tile pe_tile_8_28(
		.out_wire_3_0(vertical_tile_8_28_to_tile_7_28_0),
		.out_wire_3_1(vertical_tile_8_28_to_tile_7_28_1),
		.out_wire_3_2(vertical_tile_8_28_to_tile_7_28_2),
		.out_wire_3_3(vertical_tile_8_28_to_tile_7_28_3),
		.in_wire_3_0(vertical_tile_7_28_to_tile_8_28_0),
		.in_wire_3_1(vertical_tile_7_28_to_tile_8_28_1),
		.in_wire_3_2(vertical_tile_7_28_to_tile_8_28_2),
		.in_wire_3_3(vertical_tile_7_28_to_tile_8_28_3),
		.out_wire_1_0(vertical_tile_8_28_to_tile_9_28_0),
		.out_wire_1_1(vertical_tile_8_28_to_tile_9_28_1),
		.out_wire_1_2(vertical_tile_8_28_to_tile_9_28_2),
		.out_wire_1_3(vertical_tile_8_28_to_tile_9_28_3),
		.in_wire_1_0(vertical_tile_9_28_to_tile_8_28_0),
		.in_wire_1_1(vertical_tile_9_28_to_tile_8_28_1),
		.in_wire_1_2(vertical_tile_9_28_to_tile_8_28_2),
		.in_wire_1_3(vertical_tile_9_28_to_tile_8_28_3),
		.out_wire_2_0(horizontal_tile_8_28_to_tile_8_27_0),
		.out_wire_2_1(horizontal_tile_8_28_to_tile_8_27_1),
		.out_wire_2_2(horizontal_tile_8_28_to_tile_8_27_2),
		.out_wire_2_3(horizontal_tile_8_28_to_tile_8_27_3),
		.in_wire_2_0(horizontal_tile_8_27_to_tile_8_28_0),
		.in_wire_2_1(horizontal_tile_8_27_to_tile_8_28_1),
		.in_wire_2_2(horizontal_tile_8_27_to_tile_8_28_2),
		.in_wire_2_3(horizontal_tile_8_27_to_tile_8_28_3),
		.out_wire_0_0(horizontal_tile_8_28_to_tile_8_29_0),
		.out_wire_0_1(horizontal_tile_8_28_to_tile_8_29_1),
		.out_wire_0_2(horizontal_tile_8_28_to_tile_8_29_2),
		.out_wire_0_3(horizontal_tile_8_28_to_tile_8_29_3),
		.in_wire_0_0(horizontal_tile_8_29_to_tile_8_28_0),
		.in_wire_0_1(horizontal_tile_8_29_to_tile_8_28_1),
		.in_wire_0_2(horizontal_tile_8_29_to_tile_8_28_2),
		.in_wire_0_3(horizontal_tile_8_29_to_tile_8_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(285)
	);

	pe_tile pe_tile_8_29(
		.out_wire_3_0(vertical_tile_8_29_to_tile_7_29_0),
		.out_wire_3_1(vertical_tile_8_29_to_tile_7_29_1),
		.out_wire_3_2(vertical_tile_8_29_to_tile_7_29_2),
		.out_wire_3_3(vertical_tile_8_29_to_tile_7_29_3),
		.in_wire_3_0(vertical_tile_7_29_to_tile_8_29_0),
		.in_wire_3_1(vertical_tile_7_29_to_tile_8_29_1),
		.in_wire_3_2(vertical_tile_7_29_to_tile_8_29_2),
		.in_wire_3_3(vertical_tile_7_29_to_tile_8_29_3),
		.out_wire_1_0(vertical_tile_8_29_to_tile_9_29_0),
		.out_wire_1_1(vertical_tile_8_29_to_tile_9_29_1),
		.out_wire_1_2(vertical_tile_8_29_to_tile_9_29_2),
		.out_wire_1_3(vertical_tile_8_29_to_tile_9_29_3),
		.in_wire_1_0(vertical_tile_9_29_to_tile_8_29_0),
		.in_wire_1_1(vertical_tile_9_29_to_tile_8_29_1),
		.in_wire_1_2(vertical_tile_9_29_to_tile_8_29_2),
		.in_wire_1_3(vertical_tile_9_29_to_tile_8_29_3),
		.out_wire_2_0(horizontal_tile_8_29_to_tile_8_28_0),
		.out_wire_2_1(horizontal_tile_8_29_to_tile_8_28_1),
		.out_wire_2_2(horizontal_tile_8_29_to_tile_8_28_2),
		.out_wire_2_3(horizontal_tile_8_29_to_tile_8_28_3),
		.in_wire_2_0(horizontal_tile_8_28_to_tile_8_29_0),
		.in_wire_2_1(horizontal_tile_8_28_to_tile_8_29_1),
		.in_wire_2_2(horizontal_tile_8_28_to_tile_8_29_2),
		.in_wire_2_3(horizontal_tile_8_28_to_tile_8_29_3),
		.out_wire_0_0(horizontal_tile_8_29_to_tile_8_30_0),
		.out_wire_0_1(horizontal_tile_8_29_to_tile_8_30_1),
		.out_wire_0_2(horizontal_tile_8_29_to_tile_8_30_2),
		.out_wire_0_3(horizontal_tile_8_29_to_tile_8_30_3),
		.in_wire_0_0(horizontal_tile_8_30_to_tile_8_29_0),
		.in_wire_0_1(horizontal_tile_8_30_to_tile_8_29_1),
		.in_wire_0_2(horizontal_tile_8_30_to_tile_8_29_2),
		.in_wire_0_3(horizontal_tile_8_30_to_tile_8_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(286)
	);

	pe_tile pe_tile_8_30(
		.out_wire_3_0(vertical_tile_8_30_to_tile_7_30_0),
		.out_wire_3_1(vertical_tile_8_30_to_tile_7_30_1),
		.out_wire_3_2(vertical_tile_8_30_to_tile_7_30_2),
		.out_wire_3_3(vertical_tile_8_30_to_tile_7_30_3),
		.in_wire_3_0(vertical_tile_7_30_to_tile_8_30_0),
		.in_wire_3_1(vertical_tile_7_30_to_tile_8_30_1),
		.in_wire_3_2(vertical_tile_7_30_to_tile_8_30_2),
		.in_wire_3_3(vertical_tile_7_30_to_tile_8_30_3),
		.out_wire_1_0(vertical_tile_8_30_to_tile_9_30_0),
		.out_wire_1_1(vertical_tile_8_30_to_tile_9_30_1),
		.out_wire_1_2(vertical_tile_8_30_to_tile_9_30_2),
		.out_wire_1_3(vertical_tile_8_30_to_tile_9_30_3),
		.in_wire_1_0(vertical_tile_9_30_to_tile_8_30_0),
		.in_wire_1_1(vertical_tile_9_30_to_tile_8_30_1),
		.in_wire_1_2(vertical_tile_9_30_to_tile_8_30_2),
		.in_wire_1_3(vertical_tile_9_30_to_tile_8_30_3),
		.out_wire_2_0(horizontal_tile_8_30_to_tile_8_29_0),
		.out_wire_2_1(horizontal_tile_8_30_to_tile_8_29_1),
		.out_wire_2_2(horizontal_tile_8_30_to_tile_8_29_2),
		.out_wire_2_3(horizontal_tile_8_30_to_tile_8_29_3),
		.in_wire_2_0(horizontal_tile_8_29_to_tile_8_30_0),
		.in_wire_2_1(horizontal_tile_8_29_to_tile_8_30_1),
		.in_wire_2_2(horizontal_tile_8_29_to_tile_8_30_2),
		.in_wire_2_3(horizontal_tile_8_29_to_tile_8_30_3),
		.out_wire_0_0(horizontal_tile_8_30_to_tile_8_31_0),
		.out_wire_0_1(horizontal_tile_8_30_to_tile_8_31_1),
		.out_wire_0_2(horizontal_tile_8_30_to_tile_8_31_2),
		.out_wire_0_3(horizontal_tile_8_30_to_tile_8_31_3),
		.in_wire_0_0(horizontal_tile_8_31_to_tile_8_30_0),
		.in_wire_0_1(horizontal_tile_8_31_to_tile_8_30_1),
		.in_wire_0_2(horizontal_tile_8_31_to_tile_8_30_2),
		.in_wire_0_3(horizontal_tile_8_31_to_tile_8_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(287)
	);

	pe_tile_right pe_tile_8_31(
		.out_wire_3_0(vertical_tile_8_31_to_tile_7_31_0),
		.out_wire_3_1(vertical_tile_8_31_to_tile_7_31_1),
		.out_wire_3_2(vertical_tile_8_31_to_tile_7_31_2),
		.out_wire_3_3(vertical_tile_8_31_to_tile_7_31_3),
		.in_wire_3_0(vertical_tile_7_31_to_tile_8_31_0),
		.in_wire_3_1(vertical_tile_7_31_to_tile_8_31_1),
		.in_wire_3_2(vertical_tile_7_31_to_tile_8_31_2),
		.in_wire_3_3(vertical_tile_7_31_to_tile_8_31_3),
		.out_wire_1_0(vertical_tile_8_31_to_tile_9_31_0),
		.out_wire_1_1(vertical_tile_8_31_to_tile_9_31_1),
		.out_wire_1_2(vertical_tile_8_31_to_tile_9_31_2),
		.out_wire_1_3(vertical_tile_8_31_to_tile_9_31_3),
		.in_wire_1_0(vertical_tile_9_31_to_tile_8_31_0),
		.in_wire_1_1(vertical_tile_9_31_to_tile_8_31_1),
		.in_wire_1_2(vertical_tile_9_31_to_tile_8_31_2),
		.in_wire_1_3(vertical_tile_9_31_to_tile_8_31_3),
		.out_wire_2_0(horizontal_tile_8_31_to_tile_8_30_0),
		.out_wire_2_1(horizontal_tile_8_31_to_tile_8_30_1),
		.out_wire_2_2(horizontal_tile_8_31_to_tile_8_30_2),
		.out_wire_2_3(horizontal_tile_8_31_to_tile_8_30_3),
		.in_wire_2_0(horizontal_tile_8_30_to_tile_8_31_0),
		.in_wire_2_1(horizontal_tile_8_30_to_tile_8_31_1),
		.in_wire_2_2(horizontal_tile_8_30_to_tile_8_31_2),
		.in_wire_2_3(horizontal_tile_8_30_to_tile_8_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(288)
	);

	pe_tile_left pe_tile_9_0(
		.out_wire_3_0(vertical_tile_9_0_to_tile_8_0_0),
		.out_wire_3_1(vertical_tile_9_0_to_tile_8_0_1),
		.out_wire_3_2(vertical_tile_9_0_to_tile_8_0_2),
		.out_wire_3_3(vertical_tile_9_0_to_tile_8_0_3),
		.in_wire_3_0(vertical_tile_8_0_to_tile_9_0_0),
		.in_wire_3_1(vertical_tile_8_0_to_tile_9_0_1),
		.in_wire_3_2(vertical_tile_8_0_to_tile_9_0_2),
		.in_wire_3_3(vertical_tile_8_0_to_tile_9_0_3),
		.out_wire_1_0(vertical_tile_9_0_to_tile_10_0_0),
		.out_wire_1_1(vertical_tile_9_0_to_tile_10_0_1),
		.out_wire_1_2(vertical_tile_9_0_to_tile_10_0_2),
		.out_wire_1_3(vertical_tile_9_0_to_tile_10_0_3),
		.in_wire_1_0(vertical_tile_10_0_to_tile_9_0_0),
		.in_wire_1_1(vertical_tile_10_0_to_tile_9_0_1),
		.in_wire_1_2(vertical_tile_10_0_to_tile_9_0_2),
		.in_wire_1_3(vertical_tile_10_0_to_tile_9_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_9_0_to_tile_9_1_0),
		.out_wire_0_1(horizontal_tile_9_0_to_tile_9_1_1),
		.out_wire_0_2(horizontal_tile_9_0_to_tile_9_1_2),
		.out_wire_0_3(horizontal_tile_9_0_to_tile_9_1_3),
		.in_wire_0_0(horizontal_tile_9_1_to_tile_9_0_0),
		.in_wire_0_1(horizontal_tile_9_1_to_tile_9_0_1),
		.in_wire_0_2(horizontal_tile_9_1_to_tile_9_0_2),
		.in_wire_0_3(horizontal_tile_9_1_to_tile_9_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(289)
	);

	pe_tile pe_tile_9_1(
		.out_wire_3_0(vertical_tile_9_1_to_tile_8_1_0),
		.out_wire_3_1(vertical_tile_9_1_to_tile_8_1_1),
		.out_wire_3_2(vertical_tile_9_1_to_tile_8_1_2),
		.out_wire_3_3(vertical_tile_9_1_to_tile_8_1_3),
		.in_wire_3_0(vertical_tile_8_1_to_tile_9_1_0),
		.in_wire_3_1(vertical_tile_8_1_to_tile_9_1_1),
		.in_wire_3_2(vertical_tile_8_1_to_tile_9_1_2),
		.in_wire_3_3(vertical_tile_8_1_to_tile_9_1_3),
		.out_wire_1_0(vertical_tile_9_1_to_tile_10_1_0),
		.out_wire_1_1(vertical_tile_9_1_to_tile_10_1_1),
		.out_wire_1_2(vertical_tile_9_1_to_tile_10_1_2),
		.out_wire_1_3(vertical_tile_9_1_to_tile_10_1_3),
		.in_wire_1_0(vertical_tile_10_1_to_tile_9_1_0),
		.in_wire_1_1(vertical_tile_10_1_to_tile_9_1_1),
		.in_wire_1_2(vertical_tile_10_1_to_tile_9_1_2),
		.in_wire_1_3(vertical_tile_10_1_to_tile_9_1_3),
		.out_wire_2_0(horizontal_tile_9_1_to_tile_9_0_0),
		.out_wire_2_1(horizontal_tile_9_1_to_tile_9_0_1),
		.out_wire_2_2(horizontal_tile_9_1_to_tile_9_0_2),
		.out_wire_2_3(horizontal_tile_9_1_to_tile_9_0_3),
		.in_wire_2_0(horizontal_tile_9_0_to_tile_9_1_0),
		.in_wire_2_1(horizontal_tile_9_0_to_tile_9_1_1),
		.in_wire_2_2(horizontal_tile_9_0_to_tile_9_1_2),
		.in_wire_2_3(horizontal_tile_9_0_to_tile_9_1_3),
		.out_wire_0_0(horizontal_tile_9_1_to_tile_9_2_0),
		.out_wire_0_1(horizontal_tile_9_1_to_tile_9_2_1),
		.out_wire_0_2(horizontal_tile_9_1_to_tile_9_2_2),
		.out_wire_0_3(horizontal_tile_9_1_to_tile_9_2_3),
		.in_wire_0_0(horizontal_tile_9_2_to_tile_9_1_0),
		.in_wire_0_1(horizontal_tile_9_2_to_tile_9_1_1),
		.in_wire_0_2(horizontal_tile_9_2_to_tile_9_1_2),
		.in_wire_0_3(horizontal_tile_9_2_to_tile_9_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(290)
	);

	pe_tile pe_tile_9_2(
		.out_wire_3_0(vertical_tile_9_2_to_tile_8_2_0),
		.out_wire_3_1(vertical_tile_9_2_to_tile_8_2_1),
		.out_wire_3_2(vertical_tile_9_2_to_tile_8_2_2),
		.out_wire_3_3(vertical_tile_9_2_to_tile_8_2_3),
		.in_wire_3_0(vertical_tile_8_2_to_tile_9_2_0),
		.in_wire_3_1(vertical_tile_8_2_to_tile_9_2_1),
		.in_wire_3_2(vertical_tile_8_2_to_tile_9_2_2),
		.in_wire_3_3(vertical_tile_8_2_to_tile_9_2_3),
		.out_wire_1_0(vertical_tile_9_2_to_tile_10_2_0),
		.out_wire_1_1(vertical_tile_9_2_to_tile_10_2_1),
		.out_wire_1_2(vertical_tile_9_2_to_tile_10_2_2),
		.out_wire_1_3(vertical_tile_9_2_to_tile_10_2_3),
		.in_wire_1_0(vertical_tile_10_2_to_tile_9_2_0),
		.in_wire_1_1(vertical_tile_10_2_to_tile_9_2_1),
		.in_wire_1_2(vertical_tile_10_2_to_tile_9_2_2),
		.in_wire_1_3(vertical_tile_10_2_to_tile_9_2_3),
		.out_wire_2_0(horizontal_tile_9_2_to_tile_9_1_0),
		.out_wire_2_1(horizontal_tile_9_2_to_tile_9_1_1),
		.out_wire_2_2(horizontal_tile_9_2_to_tile_9_1_2),
		.out_wire_2_3(horizontal_tile_9_2_to_tile_9_1_3),
		.in_wire_2_0(horizontal_tile_9_1_to_tile_9_2_0),
		.in_wire_2_1(horizontal_tile_9_1_to_tile_9_2_1),
		.in_wire_2_2(horizontal_tile_9_1_to_tile_9_2_2),
		.in_wire_2_3(horizontal_tile_9_1_to_tile_9_2_3),
		.out_wire_0_0(horizontal_tile_9_2_to_tile_9_3_0),
		.out_wire_0_1(horizontal_tile_9_2_to_tile_9_3_1),
		.out_wire_0_2(horizontal_tile_9_2_to_tile_9_3_2),
		.out_wire_0_3(horizontal_tile_9_2_to_tile_9_3_3),
		.in_wire_0_0(horizontal_tile_9_3_to_tile_9_2_0),
		.in_wire_0_1(horizontal_tile_9_3_to_tile_9_2_1),
		.in_wire_0_2(horizontal_tile_9_3_to_tile_9_2_2),
		.in_wire_0_3(horizontal_tile_9_3_to_tile_9_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(291)
	);

	pe_tile pe_tile_9_3(
		.out_wire_3_0(vertical_tile_9_3_to_tile_8_3_0),
		.out_wire_3_1(vertical_tile_9_3_to_tile_8_3_1),
		.out_wire_3_2(vertical_tile_9_3_to_tile_8_3_2),
		.out_wire_3_3(vertical_tile_9_3_to_tile_8_3_3),
		.in_wire_3_0(vertical_tile_8_3_to_tile_9_3_0),
		.in_wire_3_1(vertical_tile_8_3_to_tile_9_3_1),
		.in_wire_3_2(vertical_tile_8_3_to_tile_9_3_2),
		.in_wire_3_3(vertical_tile_8_3_to_tile_9_3_3),
		.out_wire_1_0(vertical_tile_9_3_to_tile_10_3_0),
		.out_wire_1_1(vertical_tile_9_3_to_tile_10_3_1),
		.out_wire_1_2(vertical_tile_9_3_to_tile_10_3_2),
		.out_wire_1_3(vertical_tile_9_3_to_tile_10_3_3),
		.in_wire_1_0(vertical_tile_10_3_to_tile_9_3_0),
		.in_wire_1_1(vertical_tile_10_3_to_tile_9_3_1),
		.in_wire_1_2(vertical_tile_10_3_to_tile_9_3_2),
		.in_wire_1_3(vertical_tile_10_3_to_tile_9_3_3),
		.out_wire_2_0(horizontal_tile_9_3_to_tile_9_2_0),
		.out_wire_2_1(horizontal_tile_9_3_to_tile_9_2_1),
		.out_wire_2_2(horizontal_tile_9_3_to_tile_9_2_2),
		.out_wire_2_3(horizontal_tile_9_3_to_tile_9_2_3),
		.in_wire_2_0(horizontal_tile_9_2_to_tile_9_3_0),
		.in_wire_2_1(horizontal_tile_9_2_to_tile_9_3_1),
		.in_wire_2_2(horizontal_tile_9_2_to_tile_9_3_2),
		.in_wire_2_3(horizontal_tile_9_2_to_tile_9_3_3),
		.out_wire_0_0(horizontal_tile_9_3_to_tile_9_4_0),
		.out_wire_0_1(horizontal_tile_9_3_to_tile_9_4_1),
		.out_wire_0_2(horizontal_tile_9_3_to_tile_9_4_2),
		.out_wire_0_3(horizontal_tile_9_3_to_tile_9_4_3),
		.in_wire_0_0(horizontal_tile_9_4_to_tile_9_3_0),
		.in_wire_0_1(horizontal_tile_9_4_to_tile_9_3_1),
		.in_wire_0_2(horizontal_tile_9_4_to_tile_9_3_2),
		.in_wire_0_3(horizontal_tile_9_4_to_tile_9_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(292)
	);

	pe_tile pe_tile_9_4(
		.out_wire_3_0(vertical_tile_9_4_to_tile_8_4_0),
		.out_wire_3_1(vertical_tile_9_4_to_tile_8_4_1),
		.out_wire_3_2(vertical_tile_9_4_to_tile_8_4_2),
		.out_wire_3_3(vertical_tile_9_4_to_tile_8_4_3),
		.in_wire_3_0(vertical_tile_8_4_to_tile_9_4_0),
		.in_wire_3_1(vertical_tile_8_4_to_tile_9_4_1),
		.in_wire_3_2(vertical_tile_8_4_to_tile_9_4_2),
		.in_wire_3_3(vertical_tile_8_4_to_tile_9_4_3),
		.out_wire_1_0(vertical_tile_9_4_to_tile_10_4_0),
		.out_wire_1_1(vertical_tile_9_4_to_tile_10_4_1),
		.out_wire_1_2(vertical_tile_9_4_to_tile_10_4_2),
		.out_wire_1_3(vertical_tile_9_4_to_tile_10_4_3),
		.in_wire_1_0(vertical_tile_10_4_to_tile_9_4_0),
		.in_wire_1_1(vertical_tile_10_4_to_tile_9_4_1),
		.in_wire_1_2(vertical_tile_10_4_to_tile_9_4_2),
		.in_wire_1_3(vertical_tile_10_4_to_tile_9_4_3),
		.out_wire_2_0(horizontal_tile_9_4_to_tile_9_3_0),
		.out_wire_2_1(horizontal_tile_9_4_to_tile_9_3_1),
		.out_wire_2_2(horizontal_tile_9_4_to_tile_9_3_2),
		.out_wire_2_3(horizontal_tile_9_4_to_tile_9_3_3),
		.in_wire_2_0(horizontal_tile_9_3_to_tile_9_4_0),
		.in_wire_2_1(horizontal_tile_9_3_to_tile_9_4_1),
		.in_wire_2_2(horizontal_tile_9_3_to_tile_9_4_2),
		.in_wire_2_3(horizontal_tile_9_3_to_tile_9_4_3),
		.out_wire_0_0(horizontal_tile_9_4_to_tile_9_5_0),
		.out_wire_0_1(horizontal_tile_9_4_to_tile_9_5_1),
		.out_wire_0_2(horizontal_tile_9_4_to_tile_9_5_2),
		.out_wire_0_3(horizontal_tile_9_4_to_tile_9_5_3),
		.in_wire_0_0(horizontal_tile_9_5_to_tile_9_4_0),
		.in_wire_0_1(horizontal_tile_9_5_to_tile_9_4_1),
		.in_wire_0_2(horizontal_tile_9_5_to_tile_9_4_2),
		.in_wire_0_3(horizontal_tile_9_5_to_tile_9_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(293)
	);

	pe_tile pe_tile_9_5(
		.out_wire_3_0(vertical_tile_9_5_to_tile_8_5_0),
		.out_wire_3_1(vertical_tile_9_5_to_tile_8_5_1),
		.out_wire_3_2(vertical_tile_9_5_to_tile_8_5_2),
		.out_wire_3_3(vertical_tile_9_5_to_tile_8_5_3),
		.in_wire_3_0(vertical_tile_8_5_to_tile_9_5_0),
		.in_wire_3_1(vertical_tile_8_5_to_tile_9_5_1),
		.in_wire_3_2(vertical_tile_8_5_to_tile_9_5_2),
		.in_wire_3_3(vertical_tile_8_5_to_tile_9_5_3),
		.out_wire_1_0(vertical_tile_9_5_to_tile_10_5_0),
		.out_wire_1_1(vertical_tile_9_5_to_tile_10_5_1),
		.out_wire_1_2(vertical_tile_9_5_to_tile_10_5_2),
		.out_wire_1_3(vertical_tile_9_5_to_tile_10_5_3),
		.in_wire_1_0(vertical_tile_10_5_to_tile_9_5_0),
		.in_wire_1_1(vertical_tile_10_5_to_tile_9_5_1),
		.in_wire_1_2(vertical_tile_10_5_to_tile_9_5_2),
		.in_wire_1_3(vertical_tile_10_5_to_tile_9_5_3),
		.out_wire_2_0(horizontal_tile_9_5_to_tile_9_4_0),
		.out_wire_2_1(horizontal_tile_9_5_to_tile_9_4_1),
		.out_wire_2_2(horizontal_tile_9_5_to_tile_9_4_2),
		.out_wire_2_3(horizontal_tile_9_5_to_tile_9_4_3),
		.in_wire_2_0(horizontal_tile_9_4_to_tile_9_5_0),
		.in_wire_2_1(horizontal_tile_9_4_to_tile_9_5_1),
		.in_wire_2_2(horizontal_tile_9_4_to_tile_9_5_2),
		.in_wire_2_3(horizontal_tile_9_4_to_tile_9_5_3),
		.out_wire_0_0(horizontal_tile_9_5_to_tile_9_6_0),
		.out_wire_0_1(horizontal_tile_9_5_to_tile_9_6_1),
		.out_wire_0_2(horizontal_tile_9_5_to_tile_9_6_2),
		.out_wire_0_3(horizontal_tile_9_5_to_tile_9_6_3),
		.in_wire_0_0(horizontal_tile_9_6_to_tile_9_5_0),
		.in_wire_0_1(horizontal_tile_9_6_to_tile_9_5_1),
		.in_wire_0_2(horizontal_tile_9_6_to_tile_9_5_2),
		.in_wire_0_3(horizontal_tile_9_6_to_tile_9_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(294)
	);

	pe_tile pe_tile_9_6(
		.out_wire_3_0(vertical_tile_9_6_to_tile_8_6_0),
		.out_wire_3_1(vertical_tile_9_6_to_tile_8_6_1),
		.out_wire_3_2(vertical_tile_9_6_to_tile_8_6_2),
		.out_wire_3_3(vertical_tile_9_6_to_tile_8_6_3),
		.in_wire_3_0(vertical_tile_8_6_to_tile_9_6_0),
		.in_wire_3_1(vertical_tile_8_6_to_tile_9_6_1),
		.in_wire_3_2(vertical_tile_8_6_to_tile_9_6_2),
		.in_wire_3_3(vertical_tile_8_6_to_tile_9_6_3),
		.out_wire_1_0(vertical_tile_9_6_to_tile_10_6_0),
		.out_wire_1_1(vertical_tile_9_6_to_tile_10_6_1),
		.out_wire_1_2(vertical_tile_9_6_to_tile_10_6_2),
		.out_wire_1_3(vertical_tile_9_6_to_tile_10_6_3),
		.in_wire_1_0(vertical_tile_10_6_to_tile_9_6_0),
		.in_wire_1_1(vertical_tile_10_6_to_tile_9_6_1),
		.in_wire_1_2(vertical_tile_10_6_to_tile_9_6_2),
		.in_wire_1_3(vertical_tile_10_6_to_tile_9_6_3),
		.out_wire_2_0(horizontal_tile_9_6_to_tile_9_5_0),
		.out_wire_2_1(horizontal_tile_9_6_to_tile_9_5_1),
		.out_wire_2_2(horizontal_tile_9_6_to_tile_9_5_2),
		.out_wire_2_3(horizontal_tile_9_6_to_tile_9_5_3),
		.in_wire_2_0(horizontal_tile_9_5_to_tile_9_6_0),
		.in_wire_2_1(horizontal_tile_9_5_to_tile_9_6_1),
		.in_wire_2_2(horizontal_tile_9_5_to_tile_9_6_2),
		.in_wire_2_3(horizontal_tile_9_5_to_tile_9_6_3),
		.out_wire_0_0(horizontal_tile_9_6_to_tile_9_7_0),
		.out_wire_0_1(horizontal_tile_9_6_to_tile_9_7_1),
		.out_wire_0_2(horizontal_tile_9_6_to_tile_9_7_2),
		.out_wire_0_3(horizontal_tile_9_6_to_tile_9_7_3),
		.in_wire_0_0(horizontal_tile_9_7_to_tile_9_6_0),
		.in_wire_0_1(horizontal_tile_9_7_to_tile_9_6_1),
		.in_wire_0_2(horizontal_tile_9_7_to_tile_9_6_2),
		.in_wire_0_3(horizontal_tile_9_7_to_tile_9_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(295)
	);

	pe_tile pe_tile_9_7(
		.out_wire_3_0(vertical_tile_9_7_to_tile_8_7_0),
		.out_wire_3_1(vertical_tile_9_7_to_tile_8_7_1),
		.out_wire_3_2(vertical_tile_9_7_to_tile_8_7_2),
		.out_wire_3_3(vertical_tile_9_7_to_tile_8_7_3),
		.in_wire_3_0(vertical_tile_8_7_to_tile_9_7_0),
		.in_wire_3_1(vertical_tile_8_7_to_tile_9_7_1),
		.in_wire_3_2(vertical_tile_8_7_to_tile_9_7_2),
		.in_wire_3_3(vertical_tile_8_7_to_tile_9_7_3),
		.out_wire_1_0(vertical_tile_9_7_to_tile_10_7_0),
		.out_wire_1_1(vertical_tile_9_7_to_tile_10_7_1),
		.out_wire_1_2(vertical_tile_9_7_to_tile_10_7_2),
		.out_wire_1_3(vertical_tile_9_7_to_tile_10_7_3),
		.in_wire_1_0(vertical_tile_10_7_to_tile_9_7_0),
		.in_wire_1_1(vertical_tile_10_7_to_tile_9_7_1),
		.in_wire_1_2(vertical_tile_10_7_to_tile_9_7_2),
		.in_wire_1_3(vertical_tile_10_7_to_tile_9_7_3),
		.out_wire_2_0(horizontal_tile_9_7_to_tile_9_6_0),
		.out_wire_2_1(horizontal_tile_9_7_to_tile_9_6_1),
		.out_wire_2_2(horizontal_tile_9_7_to_tile_9_6_2),
		.out_wire_2_3(horizontal_tile_9_7_to_tile_9_6_3),
		.in_wire_2_0(horizontal_tile_9_6_to_tile_9_7_0),
		.in_wire_2_1(horizontal_tile_9_6_to_tile_9_7_1),
		.in_wire_2_2(horizontal_tile_9_6_to_tile_9_7_2),
		.in_wire_2_3(horizontal_tile_9_6_to_tile_9_7_3),
		.out_wire_0_0(horizontal_tile_9_7_to_tile_9_8_0),
		.out_wire_0_1(horizontal_tile_9_7_to_tile_9_8_1),
		.out_wire_0_2(horizontal_tile_9_7_to_tile_9_8_2),
		.out_wire_0_3(horizontal_tile_9_7_to_tile_9_8_3),
		.in_wire_0_0(horizontal_tile_9_8_to_tile_9_7_0),
		.in_wire_0_1(horizontal_tile_9_8_to_tile_9_7_1),
		.in_wire_0_2(horizontal_tile_9_8_to_tile_9_7_2),
		.in_wire_0_3(horizontal_tile_9_8_to_tile_9_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(296)
	);

	pe_tile pe_tile_9_8(
		.out_wire_3_0(vertical_tile_9_8_to_tile_8_8_0),
		.out_wire_3_1(vertical_tile_9_8_to_tile_8_8_1),
		.out_wire_3_2(vertical_tile_9_8_to_tile_8_8_2),
		.out_wire_3_3(vertical_tile_9_8_to_tile_8_8_3),
		.in_wire_3_0(vertical_tile_8_8_to_tile_9_8_0),
		.in_wire_3_1(vertical_tile_8_8_to_tile_9_8_1),
		.in_wire_3_2(vertical_tile_8_8_to_tile_9_8_2),
		.in_wire_3_3(vertical_tile_8_8_to_tile_9_8_3),
		.out_wire_1_0(vertical_tile_9_8_to_tile_10_8_0),
		.out_wire_1_1(vertical_tile_9_8_to_tile_10_8_1),
		.out_wire_1_2(vertical_tile_9_8_to_tile_10_8_2),
		.out_wire_1_3(vertical_tile_9_8_to_tile_10_8_3),
		.in_wire_1_0(vertical_tile_10_8_to_tile_9_8_0),
		.in_wire_1_1(vertical_tile_10_8_to_tile_9_8_1),
		.in_wire_1_2(vertical_tile_10_8_to_tile_9_8_2),
		.in_wire_1_3(vertical_tile_10_8_to_tile_9_8_3),
		.out_wire_2_0(horizontal_tile_9_8_to_tile_9_7_0),
		.out_wire_2_1(horizontal_tile_9_8_to_tile_9_7_1),
		.out_wire_2_2(horizontal_tile_9_8_to_tile_9_7_2),
		.out_wire_2_3(horizontal_tile_9_8_to_tile_9_7_3),
		.in_wire_2_0(horizontal_tile_9_7_to_tile_9_8_0),
		.in_wire_2_1(horizontal_tile_9_7_to_tile_9_8_1),
		.in_wire_2_2(horizontal_tile_9_7_to_tile_9_8_2),
		.in_wire_2_3(horizontal_tile_9_7_to_tile_9_8_3),
		.out_wire_0_0(horizontal_tile_9_8_to_tile_9_9_0),
		.out_wire_0_1(horizontal_tile_9_8_to_tile_9_9_1),
		.out_wire_0_2(horizontal_tile_9_8_to_tile_9_9_2),
		.out_wire_0_3(horizontal_tile_9_8_to_tile_9_9_3),
		.in_wire_0_0(horizontal_tile_9_9_to_tile_9_8_0),
		.in_wire_0_1(horizontal_tile_9_9_to_tile_9_8_1),
		.in_wire_0_2(horizontal_tile_9_9_to_tile_9_8_2),
		.in_wire_0_3(horizontal_tile_9_9_to_tile_9_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(297)
	);

	pe_tile pe_tile_9_9(
		.out_wire_3_0(vertical_tile_9_9_to_tile_8_9_0),
		.out_wire_3_1(vertical_tile_9_9_to_tile_8_9_1),
		.out_wire_3_2(vertical_tile_9_9_to_tile_8_9_2),
		.out_wire_3_3(vertical_tile_9_9_to_tile_8_9_3),
		.in_wire_3_0(vertical_tile_8_9_to_tile_9_9_0),
		.in_wire_3_1(vertical_tile_8_9_to_tile_9_9_1),
		.in_wire_3_2(vertical_tile_8_9_to_tile_9_9_2),
		.in_wire_3_3(vertical_tile_8_9_to_tile_9_9_3),
		.out_wire_1_0(vertical_tile_9_9_to_tile_10_9_0),
		.out_wire_1_1(vertical_tile_9_9_to_tile_10_9_1),
		.out_wire_1_2(vertical_tile_9_9_to_tile_10_9_2),
		.out_wire_1_3(vertical_tile_9_9_to_tile_10_9_3),
		.in_wire_1_0(vertical_tile_10_9_to_tile_9_9_0),
		.in_wire_1_1(vertical_tile_10_9_to_tile_9_9_1),
		.in_wire_1_2(vertical_tile_10_9_to_tile_9_9_2),
		.in_wire_1_3(vertical_tile_10_9_to_tile_9_9_3),
		.out_wire_2_0(horizontal_tile_9_9_to_tile_9_8_0),
		.out_wire_2_1(horizontal_tile_9_9_to_tile_9_8_1),
		.out_wire_2_2(horizontal_tile_9_9_to_tile_9_8_2),
		.out_wire_2_3(horizontal_tile_9_9_to_tile_9_8_3),
		.in_wire_2_0(horizontal_tile_9_8_to_tile_9_9_0),
		.in_wire_2_1(horizontal_tile_9_8_to_tile_9_9_1),
		.in_wire_2_2(horizontal_tile_9_8_to_tile_9_9_2),
		.in_wire_2_3(horizontal_tile_9_8_to_tile_9_9_3),
		.out_wire_0_0(horizontal_tile_9_9_to_tile_9_10_0),
		.out_wire_0_1(horizontal_tile_9_9_to_tile_9_10_1),
		.out_wire_0_2(horizontal_tile_9_9_to_tile_9_10_2),
		.out_wire_0_3(horizontal_tile_9_9_to_tile_9_10_3),
		.in_wire_0_0(horizontal_tile_9_10_to_tile_9_9_0),
		.in_wire_0_1(horizontal_tile_9_10_to_tile_9_9_1),
		.in_wire_0_2(horizontal_tile_9_10_to_tile_9_9_2),
		.in_wire_0_3(horizontal_tile_9_10_to_tile_9_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(298)
	);

	pe_tile pe_tile_9_10(
		.out_wire_3_0(vertical_tile_9_10_to_tile_8_10_0),
		.out_wire_3_1(vertical_tile_9_10_to_tile_8_10_1),
		.out_wire_3_2(vertical_tile_9_10_to_tile_8_10_2),
		.out_wire_3_3(vertical_tile_9_10_to_tile_8_10_3),
		.in_wire_3_0(vertical_tile_8_10_to_tile_9_10_0),
		.in_wire_3_1(vertical_tile_8_10_to_tile_9_10_1),
		.in_wire_3_2(vertical_tile_8_10_to_tile_9_10_2),
		.in_wire_3_3(vertical_tile_8_10_to_tile_9_10_3),
		.out_wire_1_0(vertical_tile_9_10_to_tile_10_10_0),
		.out_wire_1_1(vertical_tile_9_10_to_tile_10_10_1),
		.out_wire_1_2(vertical_tile_9_10_to_tile_10_10_2),
		.out_wire_1_3(vertical_tile_9_10_to_tile_10_10_3),
		.in_wire_1_0(vertical_tile_10_10_to_tile_9_10_0),
		.in_wire_1_1(vertical_tile_10_10_to_tile_9_10_1),
		.in_wire_1_2(vertical_tile_10_10_to_tile_9_10_2),
		.in_wire_1_3(vertical_tile_10_10_to_tile_9_10_3),
		.out_wire_2_0(horizontal_tile_9_10_to_tile_9_9_0),
		.out_wire_2_1(horizontal_tile_9_10_to_tile_9_9_1),
		.out_wire_2_2(horizontal_tile_9_10_to_tile_9_9_2),
		.out_wire_2_3(horizontal_tile_9_10_to_tile_9_9_3),
		.in_wire_2_0(horizontal_tile_9_9_to_tile_9_10_0),
		.in_wire_2_1(horizontal_tile_9_9_to_tile_9_10_1),
		.in_wire_2_2(horizontal_tile_9_9_to_tile_9_10_2),
		.in_wire_2_3(horizontal_tile_9_9_to_tile_9_10_3),
		.out_wire_0_0(horizontal_tile_9_10_to_tile_9_11_0),
		.out_wire_0_1(horizontal_tile_9_10_to_tile_9_11_1),
		.out_wire_0_2(horizontal_tile_9_10_to_tile_9_11_2),
		.out_wire_0_3(horizontal_tile_9_10_to_tile_9_11_3),
		.in_wire_0_0(horizontal_tile_9_11_to_tile_9_10_0),
		.in_wire_0_1(horizontal_tile_9_11_to_tile_9_10_1),
		.in_wire_0_2(horizontal_tile_9_11_to_tile_9_10_2),
		.in_wire_0_3(horizontal_tile_9_11_to_tile_9_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(299)
	);

	pe_tile pe_tile_9_11(
		.out_wire_3_0(vertical_tile_9_11_to_tile_8_11_0),
		.out_wire_3_1(vertical_tile_9_11_to_tile_8_11_1),
		.out_wire_3_2(vertical_tile_9_11_to_tile_8_11_2),
		.out_wire_3_3(vertical_tile_9_11_to_tile_8_11_3),
		.in_wire_3_0(vertical_tile_8_11_to_tile_9_11_0),
		.in_wire_3_1(vertical_tile_8_11_to_tile_9_11_1),
		.in_wire_3_2(vertical_tile_8_11_to_tile_9_11_2),
		.in_wire_3_3(vertical_tile_8_11_to_tile_9_11_3),
		.out_wire_1_0(vertical_tile_9_11_to_tile_10_11_0),
		.out_wire_1_1(vertical_tile_9_11_to_tile_10_11_1),
		.out_wire_1_2(vertical_tile_9_11_to_tile_10_11_2),
		.out_wire_1_3(vertical_tile_9_11_to_tile_10_11_3),
		.in_wire_1_0(vertical_tile_10_11_to_tile_9_11_0),
		.in_wire_1_1(vertical_tile_10_11_to_tile_9_11_1),
		.in_wire_1_2(vertical_tile_10_11_to_tile_9_11_2),
		.in_wire_1_3(vertical_tile_10_11_to_tile_9_11_3),
		.out_wire_2_0(horizontal_tile_9_11_to_tile_9_10_0),
		.out_wire_2_1(horizontal_tile_9_11_to_tile_9_10_1),
		.out_wire_2_2(horizontal_tile_9_11_to_tile_9_10_2),
		.out_wire_2_3(horizontal_tile_9_11_to_tile_9_10_3),
		.in_wire_2_0(horizontal_tile_9_10_to_tile_9_11_0),
		.in_wire_2_1(horizontal_tile_9_10_to_tile_9_11_1),
		.in_wire_2_2(horizontal_tile_9_10_to_tile_9_11_2),
		.in_wire_2_3(horizontal_tile_9_10_to_tile_9_11_3),
		.out_wire_0_0(horizontal_tile_9_11_to_tile_9_12_0),
		.out_wire_0_1(horizontal_tile_9_11_to_tile_9_12_1),
		.out_wire_0_2(horizontal_tile_9_11_to_tile_9_12_2),
		.out_wire_0_3(horizontal_tile_9_11_to_tile_9_12_3),
		.in_wire_0_0(horizontal_tile_9_12_to_tile_9_11_0),
		.in_wire_0_1(horizontal_tile_9_12_to_tile_9_11_1),
		.in_wire_0_2(horizontal_tile_9_12_to_tile_9_11_2),
		.in_wire_0_3(horizontal_tile_9_12_to_tile_9_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(300)
	);

	pe_tile pe_tile_9_12(
		.out_wire_3_0(vertical_tile_9_12_to_tile_8_12_0),
		.out_wire_3_1(vertical_tile_9_12_to_tile_8_12_1),
		.out_wire_3_2(vertical_tile_9_12_to_tile_8_12_2),
		.out_wire_3_3(vertical_tile_9_12_to_tile_8_12_3),
		.in_wire_3_0(vertical_tile_8_12_to_tile_9_12_0),
		.in_wire_3_1(vertical_tile_8_12_to_tile_9_12_1),
		.in_wire_3_2(vertical_tile_8_12_to_tile_9_12_2),
		.in_wire_3_3(vertical_tile_8_12_to_tile_9_12_3),
		.out_wire_1_0(vertical_tile_9_12_to_tile_10_12_0),
		.out_wire_1_1(vertical_tile_9_12_to_tile_10_12_1),
		.out_wire_1_2(vertical_tile_9_12_to_tile_10_12_2),
		.out_wire_1_3(vertical_tile_9_12_to_tile_10_12_3),
		.in_wire_1_0(vertical_tile_10_12_to_tile_9_12_0),
		.in_wire_1_1(vertical_tile_10_12_to_tile_9_12_1),
		.in_wire_1_2(vertical_tile_10_12_to_tile_9_12_2),
		.in_wire_1_3(vertical_tile_10_12_to_tile_9_12_3),
		.out_wire_2_0(horizontal_tile_9_12_to_tile_9_11_0),
		.out_wire_2_1(horizontal_tile_9_12_to_tile_9_11_1),
		.out_wire_2_2(horizontal_tile_9_12_to_tile_9_11_2),
		.out_wire_2_3(horizontal_tile_9_12_to_tile_9_11_3),
		.in_wire_2_0(horizontal_tile_9_11_to_tile_9_12_0),
		.in_wire_2_1(horizontal_tile_9_11_to_tile_9_12_1),
		.in_wire_2_2(horizontal_tile_9_11_to_tile_9_12_2),
		.in_wire_2_3(horizontal_tile_9_11_to_tile_9_12_3),
		.out_wire_0_0(horizontal_tile_9_12_to_tile_9_13_0),
		.out_wire_0_1(horizontal_tile_9_12_to_tile_9_13_1),
		.out_wire_0_2(horizontal_tile_9_12_to_tile_9_13_2),
		.out_wire_0_3(horizontal_tile_9_12_to_tile_9_13_3),
		.in_wire_0_0(horizontal_tile_9_13_to_tile_9_12_0),
		.in_wire_0_1(horizontal_tile_9_13_to_tile_9_12_1),
		.in_wire_0_2(horizontal_tile_9_13_to_tile_9_12_2),
		.in_wire_0_3(horizontal_tile_9_13_to_tile_9_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(301)
	);

	pe_tile pe_tile_9_13(
		.out_wire_3_0(vertical_tile_9_13_to_tile_8_13_0),
		.out_wire_3_1(vertical_tile_9_13_to_tile_8_13_1),
		.out_wire_3_2(vertical_tile_9_13_to_tile_8_13_2),
		.out_wire_3_3(vertical_tile_9_13_to_tile_8_13_3),
		.in_wire_3_0(vertical_tile_8_13_to_tile_9_13_0),
		.in_wire_3_1(vertical_tile_8_13_to_tile_9_13_1),
		.in_wire_3_2(vertical_tile_8_13_to_tile_9_13_2),
		.in_wire_3_3(vertical_tile_8_13_to_tile_9_13_3),
		.out_wire_1_0(vertical_tile_9_13_to_tile_10_13_0),
		.out_wire_1_1(vertical_tile_9_13_to_tile_10_13_1),
		.out_wire_1_2(vertical_tile_9_13_to_tile_10_13_2),
		.out_wire_1_3(vertical_tile_9_13_to_tile_10_13_3),
		.in_wire_1_0(vertical_tile_10_13_to_tile_9_13_0),
		.in_wire_1_1(vertical_tile_10_13_to_tile_9_13_1),
		.in_wire_1_2(vertical_tile_10_13_to_tile_9_13_2),
		.in_wire_1_3(vertical_tile_10_13_to_tile_9_13_3),
		.out_wire_2_0(horizontal_tile_9_13_to_tile_9_12_0),
		.out_wire_2_1(horizontal_tile_9_13_to_tile_9_12_1),
		.out_wire_2_2(horizontal_tile_9_13_to_tile_9_12_2),
		.out_wire_2_3(horizontal_tile_9_13_to_tile_9_12_3),
		.in_wire_2_0(horizontal_tile_9_12_to_tile_9_13_0),
		.in_wire_2_1(horizontal_tile_9_12_to_tile_9_13_1),
		.in_wire_2_2(horizontal_tile_9_12_to_tile_9_13_2),
		.in_wire_2_3(horizontal_tile_9_12_to_tile_9_13_3),
		.out_wire_0_0(horizontal_tile_9_13_to_tile_9_14_0),
		.out_wire_0_1(horizontal_tile_9_13_to_tile_9_14_1),
		.out_wire_0_2(horizontal_tile_9_13_to_tile_9_14_2),
		.out_wire_0_3(horizontal_tile_9_13_to_tile_9_14_3),
		.in_wire_0_0(horizontal_tile_9_14_to_tile_9_13_0),
		.in_wire_0_1(horizontal_tile_9_14_to_tile_9_13_1),
		.in_wire_0_2(horizontal_tile_9_14_to_tile_9_13_2),
		.in_wire_0_3(horizontal_tile_9_14_to_tile_9_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(302)
	);

	pe_tile pe_tile_9_14(
		.out_wire_3_0(vertical_tile_9_14_to_tile_8_14_0),
		.out_wire_3_1(vertical_tile_9_14_to_tile_8_14_1),
		.out_wire_3_2(vertical_tile_9_14_to_tile_8_14_2),
		.out_wire_3_3(vertical_tile_9_14_to_tile_8_14_3),
		.in_wire_3_0(vertical_tile_8_14_to_tile_9_14_0),
		.in_wire_3_1(vertical_tile_8_14_to_tile_9_14_1),
		.in_wire_3_2(vertical_tile_8_14_to_tile_9_14_2),
		.in_wire_3_3(vertical_tile_8_14_to_tile_9_14_3),
		.out_wire_1_0(vertical_tile_9_14_to_tile_10_14_0),
		.out_wire_1_1(vertical_tile_9_14_to_tile_10_14_1),
		.out_wire_1_2(vertical_tile_9_14_to_tile_10_14_2),
		.out_wire_1_3(vertical_tile_9_14_to_tile_10_14_3),
		.in_wire_1_0(vertical_tile_10_14_to_tile_9_14_0),
		.in_wire_1_1(vertical_tile_10_14_to_tile_9_14_1),
		.in_wire_1_2(vertical_tile_10_14_to_tile_9_14_2),
		.in_wire_1_3(vertical_tile_10_14_to_tile_9_14_3),
		.out_wire_2_0(horizontal_tile_9_14_to_tile_9_13_0),
		.out_wire_2_1(horizontal_tile_9_14_to_tile_9_13_1),
		.out_wire_2_2(horizontal_tile_9_14_to_tile_9_13_2),
		.out_wire_2_3(horizontal_tile_9_14_to_tile_9_13_3),
		.in_wire_2_0(horizontal_tile_9_13_to_tile_9_14_0),
		.in_wire_2_1(horizontal_tile_9_13_to_tile_9_14_1),
		.in_wire_2_2(horizontal_tile_9_13_to_tile_9_14_2),
		.in_wire_2_3(horizontal_tile_9_13_to_tile_9_14_3),
		.out_wire_0_0(horizontal_tile_9_14_to_tile_9_15_0),
		.out_wire_0_1(horizontal_tile_9_14_to_tile_9_15_1),
		.out_wire_0_2(horizontal_tile_9_14_to_tile_9_15_2),
		.out_wire_0_3(horizontal_tile_9_14_to_tile_9_15_3),
		.in_wire_0_0(horizontal_tile_9_15_to_tile_9_14_0),
		.in_wire_0_1(horizontal_tile_9_15_to_tile_9_14_1),
		.in_wire_0_2(horizontal_tile_9_15_to_tile_9_14_2),
		.in_wire_0_3(horizontal_tile_9_15_to_tile_9_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(303)
	);

	pe_tile pe_tile_9_15(
		.out_wire_3_0(vertical_tile_9_15_to_tile_8_15_0),
		.out_wire_3_1(vertical_tile_9_15_to_tile_8_15_1),
		.out_wire_3_2(vertical_tile_9_15_to_tile_8_15_2),
		.out_wire_3_3(vertical_tile_9_15_to_tile_8_15_3),
		.in_wire_3_0(vertical_tile_8_15_to_tile_9_15_0),
		.in_wire_3_1(vertical_tile_8_15_to_tile_9_15_1),
		.in_wire_3_2(vertical_tile_8_15_to_tile_9_15_2),
		.in_wire_3_3(vertical_tile_8_15_to_tile_9_15_3),
		.out_wire_1_0(vertical_tile_9_15_to_tile_10_15_0),
		.out_wire_1_1(vertical_tile_9_15_to_tile_10_15_1),
		.out_wire_1_2(vertical_tile_9_15_to_tile_10_15_2),
		.out_wire_1_3(vertical_tile_9_15_to_tile_10_15_3),
		.in_wire_1_0(vertical_tile_10_15_to_tile_9_15_0),
		.in_wire_1_1(vertical_tile_10_15_to_tile_9_15_1),
		.in_wire_1_2(vertical_tile_10_15_to_tile_9_15_2),
		.in_wire_1_3(vertical_tile_10_15_to_tile_9_15_3),
		.out_wire_2_0(horizontal_tile_9_15_to_tile_9_14_0),
		.out_wire_2_1(horizontal_tile_9_15_to_tile_9_14_1),
		.out_wire_2_2(horizontal_tile_9_15_to_tile_9_14_2),
		.out_wire_2_3(horizontal_tile_9_15_to_tile_9_14_3),
		.in_wire_2_0(horizontal_tile_9_14_to_tile_9_15_0),
		.in_wire_2_1(horizontal_tile_9_14_to_tile_9_15_1),
		.in_wire_2_2(horizontal_tile_9_14_to_tile_9_15_2),
		.in_wire_2_3(horizontal_tile_9_14_to_tile_9_15_3),
		.out_wire_0_0(horizontal_tile_9_15_to_tile_9_16_0),
		.out_wire_0_1(horizontal_tile_9_15_to_tile_9_16_1),
		.out_wire_0_2(horizontal_tile_9_15_to_tile_9_16_2),
		.out_wire_0_3(horizontal_tile_9_15_to_tile_9_16_3),
		.in_wire_0_0(horizontal_tile_9_16_to_tile_9_15_0),
		.in_wire_0_1(horizontal_tile_9_16_to_tile_9_15_1),
		.in_wire_0_2(horizontal_tile_9_16_to_tile_9_15_2),
		.in_wire_0_3(horizontal_tile_9_16_to_tile_9_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(304)
	);

	pe_tile pe_tile_9_16(
		.out_wire_3_0(vertical_tile_9_16_to_tile_8_16_0),
		.out_wire_3_1(vertical_tile_9_16_to_tile_8_16_1),
		.out_wire_3_2(vertical_tile_9_16_to_tile_8_16_2),
		.out_wire_3_3(vertical_tile_9_16_to_tile_8_16_3),
		.in_wire_3_0(vertical_tile_8_16_to_tile_9_16_0),
		.in_wire_3_1(vertical_tile_8_16_to_tile_9_16_1),
		.in_wire_3_2(vertical_tile_8_16_to_tile_9_16_2),
		.in_wire_3_3(vertical_tile_8_16_to_tile_9_16_3),
		.out_wire_1_0(vertical_tile_9_16_to_tile_10_16_0),
		.out_wire_1_1(vertical_tile_9_16_to_tile_10_16_1),
		.out_wire_1_2(vertical_tile_9_16_to_tile_10_16_2),
		.out_wire_1_3(vertical_tile_9_16_to_tile_10_16_3),
		.in_wire_1_0(vertical_tile_10_16_to_tile_9_16_0),
		.in_wire_1_1(vertical_tile_10_16_to_tile_9_16_1),
		.in_wire_1_2(vertical_tile_10_16_to_tile_9_16_2),
		.in_wire_1_3(vertical_tile_10_16_to_tile_9_16_3),
		.out_wire_2_0(horizontal_tile_9_16_to_tile_9_15_0),
		.out_wire_2_1(horizontal_tile_9_16_to_tile_9_15_1),
		.out_wire_2_2(horizontal_tile_9_16_to_tile_9_15_2),
		.out_wire_2_3(horizontal_tile_9_16_to_tile_9_15_3),
		.in_wire_2_0(horizontal_tile_9_15_to_tile_9_16_0),
		.in_wire_2_1(horizontal_tile_9_15_to_tile_9_16_1),
		.in_wire_2_2(horizontal_tile_9_15_to_tile_9_16_2),
		.in_wire_2_3(horizontal_tile_9_15_to_tile_9_16_3),
		.out_wire_0_0(horizontal_tile_9_16_to_tile_9_17_0),
		.out_wire_0_1(horizontal_tile_9_16_to_tile_9_17_1),
		.out_wire_0_2(horizontal_tile_9_16_to_tile_9_17_2),
		.out_wire_0_3(horizontal_tile_9_16_to_tile_9_17_3),
		.in_wire_0_0(horizontal_tile_9_17_to_tile_9_16_0),
		.in_wire_0_1(horizontal_tile_9_17_to_tile_9_16_1),
		.in_wire_0_2(horizontal_tile_9_17_to_tile_9_16_2),
		.in_wire_0_3(horizontal_tile_9_17_to_tile_9_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(305)
	);

	pe_tile pe_tile_9_17(
		.out_wire_3_0(vertical_tile_9_17_to_tile_8_17_0),
		.out_wire_3_1(vertical_tile_9_17_to_tile_8_17_1),
		.out_wire_3_2(vertical_tile_9_17_to_tile_8_17_2),
		.out_wire_3_3(vertical_tile_9_17_to_tile_8_17_3),
		.in_wire_3_0(vertical_tile_8_17_to_tile_9_17_0),
		.in_wire_3_1(vertical_tile_8_17_to_tile_9_17_1),
		.in_wire_3_2(vertical_tile_8_17_to_tile_9_17_2),
		.in_wire_3_3(vertical_tile_8_17_to_tile_9_17_3),
		.out_wire_1_0(vertical_tile_9_17_to_tile_10_17_0),
		.out_wire_1_1(vertical_tile_9_17_to_tile_10_17_1),
		.out_wire_1_2(vertical_tile_9_17_to_tile_10_17_2),
		.out_wire_1_3(vertical_tile_9_17_to_tile_10_17_3),
		.in_wire_1_0(vertical_tile_10_17_to_tile_9_17_0),
		.in_wire_1_1(vertical_tile_10_17_to_tile_9_17_1),
		.in_wire_1_2(vertical_tile_10_17_to_tile_9_17_2),
		.in_wire_1_3(vertical_tile_10_17_to_tile_9_17_3),
		.out_wire_2_0(horizontal_tile_9_17_to_tile_9_16_0),
		.out_wire_2_1(horizontal_tile_9_17_to_tile_9_16_1),
		.out_wire_2_2(horizontal_tile_9_17_to_tile_9_16_2),
		.out_wire_2_3(horizontal_tile_9_17_to_tile_9_16_3),
		.in_wire_2_0(horizontal_tile_9_16_to_tile_9_17_0),
		.in_wire_2_1(horizontal_tile_9_16_to_tile_9_17_1),
		.in_wire_2_2(horizontal_tile_9_16_to_tile_9_17_2),
		.in_wire_2_3(horizontal_tile_9_16_to_tile_9_17_3),
		.out_wire_0_0(horizontal_tile_9_17_to_tile_9_18_0),
		.out_wire_0_1(horizontal_tile_9_17_to_tile_9_18_1),
		.out_wire_0_2(horizontal_tile_9_17_to_tile_9_18_2),
		.out_wire_0_3(horizontal_tile_9_17_to_tile_9_18_3),
		.in_wire_0_0(horizontal_tile_9_18_to_tile_9_17_0),
		.in_wire_0_1(horizontal_tile_9_18_to_tile_9_17_1),
		.in_wire_0_2(horizontal_tile_9_18_to_tile_9_17_2),
		.in_wire_0_3(horizontal_tile_9_18_to_tile_9_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(306)
	);

	pe_tile pe_tile_9_18(
		.out_wire_3_0(vertical_tile_9_18_to_tile_8_18_0),
		.out_wire_3_1(vertical_tile_9_18_to_tile_8_18_1),
		.out_wire_3_2(vertical_tile_9_18_to_tile_8_18_2),
		.out_wire_3_3(vertical_tile_9_18_to_tile_8_18_3),
		.in_wire_3_0(vertical_tile_8_18_to_tile_9_18_0),
		.in_wire_3_1(vertical_tile_8_18_to_tile_9_18_1),
		.in_wire_3_2(vertical_tile_8_18_to_tile_9_18_2),
		.in_wire_3_3(vertical_tile_8_18_to_tile_9_18_3),
		.out_wire_1_0(vertical_tile_9_18_to_tile_10_18_0),
		.out_wire_1_1(vertical_tile_9_18_to_tile_10_18_1),
		.out_wire_1_2(vertical_tile_9_18_to_tile_10_18_2),
		.out_wire_1_3(vertical_tile_9_18_to_tile_10_18_3),
		.in_wire_1_0(vertical_tile_10_18_to_tile_9_18_0),
		.in_wire_1_1(vertical_tile_10_18_to_tile_9_18_1),
		.in_wire_1_2(vertical_tile_10_18_to_tile_9_18_2),
		.in_wire_1_3(vertical_tile_10_18_to_tile_9_18_3),
		.out_wire_2_0(horizontal_tile_9_18_to_tile_9_17_0),
		.out_wire_2_1(horizontal_tile_9_18_to_tile_9_17_1),
		.out_wire_2_2(horizontal_tile_9_18_to_tile_9_17_2),
		.out_wire_2_3(horizontal_tile_9_18_to_tile_9_17_3),
		.in_wire_2_0(horizontal_tile_9_17_to_tile_9_18_0),
		.in_wire_2_1(horizontal_tile_9_17_to_tile_9_18_1),
		.in_wire_2_2(horizontal_tile_9_17_to_tile_9_18_2),
		.in_wire_2_3(horizontal_tile_9_17_to_tile_9_18_3),
		.out_wire_0_0(horizontal_tile_9_18_to_tile_9_19_0),
		.out_wire_0_1(horizontal_tile_9_18_to_tile_9_19_1),
		.out_wire_0_2(horizontal_tile_9_18_to_tile_9_19_2),
		.out_wire_0_3(horizontal_tile_9_18_to_tile_9_19_3),
		.in_wire_0_0(horizontal_tile_9_19_to_tile_9_18_0),
		.in_wire_0_1(horizontal_tile_9_19_to_tile_9_18_1),
		.in_wire_0_2(horizontal_tile_9_19_to_tile_9_18_2),
		.in_wire_0_3(horizontal_tile_9_19_to_tile_9_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(307)
	);

	pe_tile pe_tile_9_19(
		.out_wire_3_0(vertical_tile_9_19_to_tile_8_19_0),
		.out_wire_3_1(vertical_tile_9_19_to_tile_8_19_1),
		.out_wire_3_2(vertical_tile_9_19_to_tile_8_19_2),
		.out_wire_3_3(vertical_tile_9_19_to_tile_8_19_3),
		.in_wire_3_0(vertical_tile_8_19_to_tile_9_19_0),
		.in_wire_3_1(vertical_tile_8_19_to_tile_9_19_1),
		.in_wire_3_2(vertical_tile_8_19_to_tile_9_19_2),
		.in_wire_3_3(vertical_tile_8_19_to_tile_9_19_3),
		.out_wire_1_0(vertical_tile_9_19_to_tile_10_19_0),
		.out_wire_1_1(vertical_tile_9_19_to_tile_10_19_1),
		.out_wire_1_2(vertical_tile_9_19_to_tile_10_19_2),
		.out_wire_1_3(vertical_tile_9_19_to_tile_10_19_3),
		.in_wire_1_0(vertical_tile_10_19_to_tile_9_19_0),
		.in_wire_1_1(vertical_tile_10_19_to_tile_9_19_1),
		.in_wire_1_2(vertical_tile_10_19_to_tile_9_19_2),
		.in_wire_1_3(vertical_tile_10_19_to_tile_9_19_3),
		.out_wire_2_0(horizontal_tile_9_19_to_tile_9_18_0),
		.out_wire_2_1(horizontal_tile_9_19_to_tile_9_18_1),
		.out_wire_2_2(horizontal_tile_9_19_to_tile_9_18_2),
		.out_wire_2_3(horizontal_tile_9_19_to_tile_9_18_3),
		.in_wire_2_0(horizontal_tile_9_18_to_tile_9_19_0),
		.in_wire_2_1(horizontal_tile_9_18_to_tile_9_19_1),
		.in_wire_2_2(horizontal_tile_9_18_to_tile_9_19_2),
		.in_wire_2_3(horizontal_tile_9_18_to_tile_9_19_3),
		.out_wire_0_0(horizontal_tile_9_19_to_tile_9_20_0),
		.out_wire_0_1(horizontal_tile_9_19_to_tile_9_20_1),
		.out_wire_0_2(horizontal_tile_9_19_to_tile_9_20_2),
		.out_wire_0_3(horizontal_tile_9_19_to_tile_9_20_3),
		.in_wire_0_0(horizontal_tile_9_20_to_tile_9_19_0),
		.in_wire_0_1(horizontal_tile_9_20_to_tile_9_19_1),
		.in_wire_0_2(horizontal_tile_9_20_to_tile_9_19_2),
		.in_wire_0_3(horizontal_tile_9_20_to_tile_9_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(308)
	);

	pe_tile pe_tile_9_20(
		.out_wire_3_0(vertical_tile_9_20_to_tile_8_20_0),
		.out_wire_3_1(vertical_tile_9_20_to_tile_8_20_1),
		.out_wire_3_2(vertical_tile_9_20_to_tile_8_20_2),
		.out_wire_3_3(vertical_tile_9_20_to_tile_8_20_3),
		.in_wire_3_0(vertical_tile_8_20_to_tile_9_20_0),
		.in_wire_3_1(vertical_tile_8_20_to_tile_9_20_1),
		.in_wire_3_2(vertical_tile_8_20_to_tile_9_20_2),
		.in_wire_3_3(vertical_tile_8_20_to_tile_9_20_3),
		.out_wire_1_0(vertical_tile_9_20_to_tile_10_20_0),
		.out_wire_1_1(vertical_tile_9_20_to_tile_10_20_1),
		.out_wire_1_2(vertical_tile_9_20_to_tile_10_20_2),
		.out_wire_1_3(vertical_tile_9_20_to_tile_10_20_3),
		.in_wire_1_0(vertical_tile_10_20_to_tile_9_20_0),
		.in_wire_1_1(vertical_tile_10_20_to_tile_9_20_1),
		.in_wire_1_2(vertical_tile_10_20_to_tile_9_20_2),
		.in_wire_1_3(vertical_tile_10_20_to_tile_9_20_3),
		.out_wire_2_0(horizontal_tile_9_20_to_tile_9_19_0),
		.out_wire_2_1(horizontal_tile_9_20_to_tile_9_19_1),
		.out_wire_2_2(horizontal_tile_9_20_to_tile_9_19_2),
		.out_wire_2_3(horizontal_tile_9_20_to_tile_9_19_3),
		.in_wire_2_0(horizontal_tile_9_19_to_tile_9_20_0),
		.in_wire_2_1(horizontal_tile_9_19_to_tile_9_20_1),
		.in_wire_2_2(horizontal_tile_9_19_to_tile_9_20_2),
		.in_wire_2_3(horizontal_tile_9_19_to_tile_9_20_3),
		.out_wire_0_0(horizontal_tile_9_20_to_tile_9_21_0),
		.out_wire_0_1(horizontal_tile_9_20_to_tile_9_21_1),
		.out_wire_0_2(horizontal_tile_9_20_to_tile_9_21_2),
		.out_wire_0_3(horizontal_tile_9_20_to_tile_9_21_3),
		.in_wire_0_0(horizontal_tile_9_21_to_tile_9_20_0),
		.in_wire_0_1(horizontal_tile_9_21_to_tile_9_20_1),
		.in_wire_0_2(horizontal_tile_9_21_to_tile_9_20_2),
		.in_wire_0_3(horizontal_tile_9_21_to_tile_9_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(309)
	);

	pe_tile pe_tile_9_21(
		.out_wire_3_0(vertical_tile_9_21_to_tile_8_21_0),
		.out_wire_3_1(vertical_tile_9_21_to_tile_8_21_1),
		.out_wire_3_2(vertical_tile_9_21_to_tile_8_21_2),
		.out_wire_3_3(vertical_tile_9_21_to_tile_8_21_3),
		.in_wire_3_0(vertical_tile_8_21_to_tile_9_21_0),
		.in_wire_3_1(vertical_tile_8_21_to_tile_9_21_1),
		.in_wire_3_2(vertical_tile_8_21_to_tile_9_21_2),
		.in_wire_3_3(vertical_tile_8_21_to_tile_9_21_3),
		.out_wire_1_0(vertical_tile_9_21_to_tile_10_21_0),
		.out_wire_1_1(vertical_tile_9_21_to_tile_10_21_1),
		.out_wire_1_2(vertical_tile_9_21_to_tile_10_21_2),
		.out_wire_1_3(vertical_tile_9_21_to_tile_10_21_3),
		.in_wire_1_0(vertical_tile_10_21_to_tile_9_21_0),
		.in_wire_1_1(vertical_tile_10_21_to_tile_9_21_1),
		.in_wire_1_2(vertical_tile_10_21_to_tile_9_21_2),
		.in_wire_1_3(vertical_tile_10_21_to_tile_9_21_3),
		.out_wire_2_0(horizontal_tile_9_21_to_tile_9_20_0),
		.out_wire_2_1(horizontal_tile_9_21_to_tile_9_20_1),
		.out_wire_2_2(horizontal_tile_9_21_to_tile_9_20_2),
		.out_wire_2_3(horizontal_tile_9_21_to_tile_9_20_3),
		.in_wire_2_0(horizontal_tile_9_20_to_tile_9_21_0),
		.in_wire_2_1(horizontal_tile_9_20_to_tile_9_21_1),
		.in_wire_2_2(horizontal_tile_9_20_to_tile_9_21_2),
		.in_wire_2_3(horizontal_tile_9_20_to_tile_9_21_3),
		.out_wire_0_0(horizontal_tile_9_21_to_tile_9_22_0),
		.out_wire_0_1(horizontal_tile_9_21_to_tile_9_22_1),
		.out_wire_0_2(horizontal_tile_9_21_to_tile_9_22_2),
		.out_wire_0_3(horizontal_tile_9_21_to_tile_9_22_3),
		.in_wire_0_0(horizontal_tile_9_22_to_tile_9_21_0),
		.in_wire_0_1(horizontal_tile_9_22_to_tile_9_21_1),
		.in_wire_0_2(horizontal_tile_9_22_to_tile_9_21_2),
		.in_wire_0_3(horizontal_tile_9_22_to_tile_9_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(310)
	);

	pe_tile pe_tile_9_22(
		.out_wire_3_0(vertical_tile_9_22_to_tile_8_22_0),
		.out_wire_3_1(vertical_tile_9_22_to_tile_8_22_1),
		.out_wire_3_2(vertical_tile_9_22_to_tile_8_22_2),
		.out_wire_3_3(vertical_tile_9_22_to_tile_8_22_3),
		.in_wire_3_0(vertical_tile_8_22_to_tile_9_22_0),
		.in_wire_3_1(vertical_tile_8_22_to_tile_9_22_1),
		.in_wire_3_2(vertical_tile_8_22_to_tile_9_22_2),
		.in_wire_3_3(vertical_tile_8_22_to_tile_9_22_3),
		.out_wire_1_0(vertical_tile_9_22_to_tile_10_22_0),
		.out_wire_1_1(vertical_tile_9_22_to_tile_10_22_1),
		.out_wire_1_2(vertical_tile_9_22_to_tile_10_22_2),
		.out_wire_1_3(vertical_tile_9_22_to_tile_10_22_3),
		.in_wire_1_0(vertical_tile_10_22_to_tile_9_22_0),
		.in_wire_1_1(vertical_tile_10_22_to_tile_9_22_1),
		.in_wire_1_2(vertical_tile_10_22_to_tile_9_22_2),
		.in_wire_1_3(vertical_tile_10_22_to_tile_9_22_3),
		.out_wire_2_0(horizontal_tile_9_22_to_tile_9_21_0),
		.out_wire_2_1(horizontal_tile_9_22_to_tile_9_21_1),
		.out_wire_2_2(horizontal_tile_9_22_to_tile_9_21_2),
		.out_wire_2_3(horizontal_tile_9_22_to_tile_9_21_3),
		.in_wire_2_0(horizontal_tile_9_21_to_tile_9_22_0),
		.in_wire_2_1(horizontal_tile_9_21_to_tile_9_22_1),
		.in_wire_2_2(horizontal_tile_9_21_to_tile_9_22_2),
		.in_wire_2_3(horizontal_tile_9_21_to_tile_9_22_3),
		.out_wire_0_0(horizontal_tile_9_22_to_tile_9_23_0),
		.out_wire_0_1(horizontal_tile_9_22_to_tile_9_23_1),
		.out_wire_0_2(horizontal_tile_9_22_to_tile_9_23_2),
		.out_wire_0_3(horizontal_tile_9_22_to_tile_9_23_3),
		.in_wire_0_0(horizontal_tile_9_23_to_tile_9_22_0),
		.in_wire_0_1(horizontal_tile_9_23_to_tile_9_22_1),
		.in_wire_0_2(horizontal_tile_9_23_to_tile_9_22_2),
		.in_wire_0_3(horizontal_tile_9_23_to_tile_9_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(311)
	);

	pe_tile pe_tile_9_23(
		.out_wire_3_0(vertical_tile_9_23_to_tile_8_23_0),
		.out_wire_3_1(vertical_tile_9_23_to_tile_8_23_1),
		.out_wire_3_2(vertical_tile_9_23_to_tile_8_23_2),
		.out_wire_3_3(vertical_tile_9_23_to_tile_8_23_3),
		.in_wire_3_0(vertical_tile_8_23_to_tile_9_23_0),
		.in_wire_3_1(vertical_tile_8_23_to_tile_9_23_1),
		.in_wire_3_2(vertical_tile_8_23_to_tile_9_23_2),
		.in_wire_3_3(vertical_tile_8_23_to_tile_9_23_3),
		.out_wire_1_0(vertical_tile_9_23_to_tile_10_23_0),
		.out_wire_1_1(vertical_tile_9_23_to_tile_10_23_1),
		.out_wire_1_2(vertical_tile_9_23_to_tile_10_23_2),
		.out_wire_1_3(vertical_tile_9_23_to_tile_10_23_3),
		.in_wire_1_0(vertical_tile_10_23_to_tile_9_23_0),
		.in_wire_1_1(vertical_tile_10_23_to_tile_9_23_1),
		.in_wire_1_2(vertical_tile_10_23_to_tile_9_23_2),
		.in_wire_1_3(vertical_tile_10_23_to_tile_9_23_3),
		.out_wire_2_0(horizontal_tile_9_23_to_tile_9_22_0),
		.out_wire_2_1(horizontal_tile_9_23_to_tile_9_22_1),
		.out_wire_2_2(horizontal_tile_9_23_to_tile_9_22_2),
		.out_wire_2_3(horizontal_tile_9_23_to_tile_9_22_3),
		.in_wire_2_0(horizontal_tile_9_22_to_tile_9_23_0),
		.in_wire_2_1(horizontal_tile_9_22_to_tile_9_23_1),
		.in_wire_2_2(horizontal_tile_9_22_to_tile_9_23_2),
		.in_wire_2_3(horizontal_tile_9_22_to_tile_9_23_3),
		.out_wire_0_0(horizontal_tile_9_23_to_tile_9_24_0),
		.out_wire_0_1(horizontal_tile_9_23_to_tile_9_24_1),
		.out_wire_0_2(horizontal_tile_9_23_to_tile_9_24_2),
		.out_wire_0_3(horizontal_tile_9_23_to_tile_9_24_3),
		.in_wire_0_0(horizontal_tile_9_24_to_tile_9_23_0),
		.in_wire_0_1(horizontal_tile_9_24_to_tile_9_23_1),
		.in_wire_0_2(horizontal_tile_9_24_to_tile_9_23_2),
		.in_wire_0_3(horizontal_tile_9_24_to_tile_9_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(312)
	);

	pe_tile pe_tile_9_24(
		.out_wire_3_0(vertical_tile_9_24_to_tile_8_24_0),
		.out_wire_3_1(vertical_tile_9_24_to_tile_8_24_1),
		.out_wire_3_2(vertical_tile_9_24_to_tile_8_24_2),
		.out_wire_3_3(vertical_tile_9_24_to_tile_8_24_3),
		.in_wire_3_0(vertical_tile_8_24_to_tile_9_24_0),
		.in_wire_3_1(vertical_tile_8_24_to_tile_9_24_1),
		.in_wire_3_2(vertical_tile_8_24_to_tile_9_24_2),
		.in_wire_3_3(vertical_tile_8_24_to_tile_9_24_3),
		.out_wire_1_0(vertical_tile_9_24_to_tile_10_24_0),
		.out_wire_1_1(vertical_tile_9_24_to_tile_10_24_1),
		.out_wire_1_2(vertical_tile_9_24_to_tile_10_24_2),
		.out_wire_1_3(vertical_tile_9_24_to_tile_10_24_3),
		.in_wire_1_0(vertical_tile_10_24_to_tile_9_24_0),
		.in_wire_1_1(vertical_tile_10_24_to_tile_9_24_1),
		.in_wire_1_2(vertical_tile_10_24_to_tile_9_24_2),
		.in_wire_1_3(vertical_tile_10_24_to_tile_9_24_3),
		.out_wire_2_0(horizontal_tile_9_24_to_tile_9_23_0),
		.out_wire_2_1(horizontal_tile_9_24_to_tile_9_23_1),
		.out_wire_2_2(horizontal_tile_9_24_to_tile_9_23_2),
		.out_wire_2_3(horizontal_tile_9_24_to_tile_9_23_3),
		.in_wire_2_0(horizontal_tile_9_23_to_tile_9_24_0),
		.in_wire_2_1(horizontal_tile_9_23_to_tile_9_24_1),
		.in_wire_2_2(horizontal_tile_9_23_to_tile_9_24_2),
		.in_wire_2_3(horizontal_tile_9_23_to_tile_9_24_3),
		.out_wire_0_0(horizontal_tile_9_24_to_tile_9_25_0),
		.out_wire_0_1(horizontal_tile_9_24_to_tile_9_25_1),
		.out_wire_0_2(horizontal_tile_9_24_to_tile_9_25_2),
		.out_wire_0_3(horizontal_tile_9_24_to_tile_9_25_3),
		.in_wire_0_0(horizontal_tile_9_25_to_tile_9_24_0),
		.in_wire_0_1(horizontal_tile_9_25_to_tile_9_24_1),
		.in_wire_0_2(horizontal_tile_9_25_to_tile_9_24_2),
		.in_wire_0_3(horizontal_tile_9_25_to_tile_9_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(313)
	);

	pe_tile pe_tile_9_25(
		.out_wire_3_0(vertical_tile_9_25_to_tile_8_25_0),
		.out_wire_3_1(vertical_tile_9_25_to_tile_8_25_1),
		.out_wire_3_2(vertical_tile_9_25_to_tile_8_25_2),
		.out_wire_3_3(vertical_tile_9_25_to_tile_8_25_3),
		.in_wire_3_0(vertical_tile_8_25_to_tile_9_25_0),
		.in_wire_3_1(vertical_tile_8_25_to_tile_9_25_1),
		.in_wire_3_2(vertical_tile_8_25_to_tile_9_25_2),
		.in_wire_3_3(vertical_tile_8_25_to_tile_9_25_3),
		.out_wire_1_0(vertical_tile_9_25_to_tile_10_25_0),
		.out_wire_1_1(vertical_tile_9_25_to_tile_10_25_1),
		.out_wire_1_2(vertical_tile_9_25_to_tile_10_25_2),
		.out_wire_1_3(vertical_tile_9_25_to_tile_10_25_3),
		.in_wire_1_0(vertical_tile_10_25_to_tile_9_25_0),
		.in_wire_1_1(vertical_tile_10_25_to_tile_9_25_1),
		.in_wire_1_2(vertical_tile_10_25_to_tile_9_25_2),
		.in_wire_1_3(vertical_tile_10_25_to_tile_9_25_3),
		.out_wire_2_0(horizontal_tile_9_25_to_tile_9_24_0),
		.out_wire_2_1(horizontal_tile_9_25_to_tile_9_24_1),
		.out_wire_2_2(horizontal_tile_9_25_to_tile_9_24_2),
		.out_wire_2_3(horizontal_tile_9_25_to_tile_9_24_3),
		.in_wire_2_0(horizontal_tile_9_24_to_tile_9_25_0),
		.in_wire_2_1(horizontal_tile_9_24_to_tile_9_25_1),
		.in_wire_2_2(horizontal_tile_9_24_to_tile_9_25_2),
		.in_wire_2_3(horizontal_tile_9_24_to_tile_9_25_3),
		.out_wire_0_0(horizontal_tile_9_25_to_tile_9_26_0),
		.out_wire_0_1(horizontal_tile_9_25_to_tile_9_26_1),
		.out_wire_0_2(horizontal_tile_9_25_to_tile_9_26_2),
		.out_wire_0_3(horizontal_tile_9_25_to_tile_9_26_3),
		.in_wire_0_0(horizontal_tile_9_26_to_tile_9_25_0),
		.in_wire_0_1(horizontal_tile_9_26_to_tile_9_25_1),
		.in_wire_0_2(horizontal_tile_9_26_to_tile_9_25_2),
		.in_wire_0_3(horizontal_tile_9_26_to_tile_9_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(314)
	);

	pe_tile pe_tile_9_26(
		.out_wire_3_0(vertical_tile_9_26_to_tile_8_26_0),
		.out_wire_3_1(vertical_tile_9_26_to_tile_8_26_1),
		.out_wire_3_2(vertical_tile_9_26_to_tile_8_26_2),
		.out_wire_3_3(vertical_tile_9_26_to_tile_8_26_3),
		.in_wire_3_0(vertical_tile_8_26_to_tile_9_26_0),
		.in_wire_3_1(vertical_tile_8_26_to_tile_9_26_1),
		.in_wire_3_2(vertical_tile_8_26_to_tile_9_26_2),
		.in_wire_3_3(vertical_tile_8_26_to_tile_9_26_3),
		.out_wire_1_0(vertical_tile_9_26_to_tile_10_26_0),
		.out_wire_1_1(vertical_tile_9_26_to_tile_10_26_1),
		.out_wire_1_2(vertical_tile_9_26_to_tile_10_26_2),
		.out_wire_1_3(vertical_tile_9_26_to_tile_10_26_3),
		.in_wire_1_0(vertical_tile_10_26_to_tile_9_26_0),
		.in_wire_1_1(vertical_tile_10_26_to_tile_9_26_1),
		.in_wire_1_2(vertical_tile_10_26_to_tile_9_26_2),
		.in_wire_1_3(vertical_tile_10_26_to_tile_9_26_3),
		.out_wire_2_0(horizontal_tile_9_26_to_tile_9_25_0),
		.out_wire_2_1(horizontal_tile_9_26_to_tile_9_25_1),
		.out_wire_2_2(horizontal_tile_9_26_to_tile_9_25_2),
		.out_wire_2_3(horizontal_tile_9_26_to_tile_9_25_3),
		.in_wire_2_0(horizontal_tile_9_25_to_tile_9_26_0),
		.in_wire_2_1(horizontal_tile_9_25_to_tile_9_26_1),
		.in_wire_2_2(horizontal_tile_9_25_to_tile_9_26_2),
		.in_wire_2_3(horizontal_tile_9_25_to_tile_9_26_3),
		.out_wire_0_0(horizontal_tile_9_26_to_tile_9_27_0),
		.out_wire_0_1(horizontal_tile_9_26_to_tile_9_27_1),
		.out_wire_0_2(horizontal_tile_9_26_to_tile_9_27_2),
		.out_wire_0_3(horizontal_tile_9_26_to_tile_9_27_3),
		.in_wire_0_0(horizontal_tile_9_27_to_tile_9_26_0),
		.in_wire_0_1(horizontal_tile_9_27_to_tile_9_26_1),
		.in_wire_0_2(horizontal_tile_9_27_to_tile_9_26_2),
		.in_wire_0_3(horizontal_tile_9_27_to_tile_9_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(315)
	);

	pe_tile pe_tile_9_27(
		.out_wire_3_0(vertical_tile_9_27_to_tile_8_27_0),
		.out_wire_3_1(vertical_tile_9_27_to_tile_8_27_1),
		.out_wire_3_2(vertical_tile_9_27_to_tile_8_27_2),
		.out_wire_3_3(vertical_tile_9_27_to_tile_8_27_3),
		.in_wire_3_0(vertical_tile_8_27_to_tile_9_27_0),
		.in_wire_3_1(vertical_tile_8_27_to_tile_9_27_1),
		.in_wire_3_2(vertical_tile_8_27_to_tile_9_27_2),
		.in_wire_3_3(vertical_tile_8_27_to_tile_9_27_3),
		.out_wire_1_0(vertical_tile_9_27_to_tile_10_27_0),
		.out_wire_1_1(vertical_tile_9_27_to_tile_10_27_1),
		.out_wire_1_2(vertical_tile_9_27_to_tile_10_27_2),
		.out_wire_1_3(vertical_tile_9_27_to_tile_10_27_3),
		.in_wire_1_0(vertical_tile_10_27_to_tile_9_27_0),
		.in_wire_1_1(vertical_tile_10_27_to_tile_9_27_1),
		.in_wire_1_2(vertical_tile_10_27_to_tile_9_27_2),
		.in_wire_1_3(vertical_tile_10_27_to_tile_9_27_3),
		.out_wire_2_0(horizontal_tile_9_27_to_tile_9_26_0),
		.out_wire_2_1(horizontal_tile_9_27_to_tile_9_26_1),
		.out_wire_2_2(horizontal_tile_9_27_to_tile_9_26_2),
		.out_wire_2_3(horizontal_tile_9_27_to_tile_9_26_3),
		.in_wire_2_0(horizontal_tile_9_26_to_tile_9_27_0),
		.in_wire_2_1(horizontal_tile_9_26_to_tile_9_27_1),
		.in_wire_2_2(horizontal_tile_9_26_to_tile_9_27_2),
		.in_wire_2_3(horizontal_tile_9_26_to_tile_9_27_3),
		.out_wire_0_0(horizontal_tile_9_27_to_tile_9_28_0),
		.out_wire_0_1(horizontal_tile_9_27_to_tile_9_28_1),
		.out_wire_0_2(horizontal_tile_9_27_to_tile_9_28_2),
		.out_wire_0_3(horizontal_tile_9_27_to_tile_9_28_3),
		.in_wire_0_0(horizontal_tile_9_28_to_tile_9_27_0),
		.in_wire_0_1(horizontal_tile_9_28_to_tile_9_27_1),
		.in_wire_0_2(horizontal_tile_9_28_to_tile_9_27_2),
		.in_wire_0_3(horizontal_tile_9_28_to_tile_9_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(316)
	);

	pe_tile pe_tile_9_28(
		.out_wire_3_0(vertical_tile_9_28_to_tile_8_28_0),
		.out_wire_3_1(vertical_tile_9_28_to_tile_8_28_1),
		.out_wire_3_2(vertical_tile_9_28_to_tile_8_28_2),
		.out_wire_3_3(vertical_tile_9_28_to_tile_8_28_3),
		.in_wire_3_0(vertical_tile_8_28_to_tile_9_28_0),
		.in_wire_3_1(vertical_tile_8_28_to_tile_9_28_1),
		.in_wire_3_2(vertical_tile_8_28_to_tile_9_28_2),
		.in_wire_3_3(vertical_tile_8_28_to_tile_9_28_3),
		.out_wire_1_0(vertical_tile_9_28_to_tile_10_28_0),
		.out_wire_1_1(vertical_tile_9_28_to_tile_10_28_1),
		.out_wire_1_2(vertical_tile_9_28_to_tile_10_28_2),
		.out_wire_1_3(vertical_tile_9_28_to_tile_10_28_3),
		.in_wire_1_0(vertical_tile_10_28_to_tile_9_28_0),
		.in_wire_1_1(vertical_tile_10_28_to_tile_9_28_1),
		.in_wire_1_2(vertical_tile_10_28_to_tile_9_28_2),
		.in_wire_1_3(vertical_tile_10_28_to_tile_9_28_3),
		.out_wire_2_0(horizontal_tile_9_28_to_tile_9_27_0),
		.out_wire_2_1(horizontal_tile_9_28_to_tile_9_27_1),
		.out_wire_2_2(horizontal_tile_9_28_to_tile_9_27_2),
		.out_wire_2_3(horizontal_tile_9_28_to_tile_9_27_3),
		.in_wire_2_0(horizontal_tile_9_27_to_tile_9_28_0),
		.in_wire_2_1(horizontal_tile_9_27_to_tile_9_28_1),
		.in_wire_2_2(horizontal_tile_9_27_to_tile_9_28_2),
		.in_wire_2_3(horizontal_tile_9_27_to_tile_9_28_3),
		.out_wire_0_0(horizontal_tile_9_28_to_tile_9_29_0),
		.out_wire_0_1(horizontal_tile_9_28_to_tile_9_29_1),
		.out_wire_0_2(horizontal_tile_9_28_to_tile_9_29_2),
		.out_wire_0_3(horizontal_tile_9_28_to_tile_9_29_3),
		.in_wire_0_0(horizontal_tile_9_29_to_tile_9_28_0),
		.in_wire_0_1(horizontal_tile_9_29_to_tile_9_28_1),
		.in_wire_0_2(horizontal_tile_9_29_to_tile_9_28_2),
		.in_wire_0_3(horizontal_tile_9_29_to_tile_9_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(317)
	);

	pe_tile pe_tile_9_29(
		.out_wire_3_0(vertical_tile_9_29_to_tile_8_29_0),
		.out_wire_3_1(vertical_tile_9_29_to_tile_8_29_1),
		.out_wire_3_2(vertical_tile_9_29_to_tile_8_29_2),
		.out_wire_3_3(vertical_tile_9_29_to_tile_8_29_3),
		.in_wire_3_0(vertical_tile_8_29_to_tile_9_29_0),
		.in_wire_3_1(vertical_tile_8_29_to_tile_9_29_1),
		.in_wire_3_2(vertical_tile_8_29_to_tile_9_29_2),
		.in_wire_3_3(vertical_tile_8_29_to_tile_9_29_3),
		.out_wire_1_0(vertical_tile_9_29_to_tile_10_29_0),
		.out_wire_1_1(vertical_tile_9_29_to_tile_10_29_1),
		.out_wire_1_2(vertical_tile_9_29_to_tile_10_29_2),
		.out_wire_1_3(vertical_tile_9_29_to_tile_10_29_3),
		.in_wire_1_0(vertical_tile_10_29_to_tile_9_29_0),
		.in_wire_1_1(vertical_tile_10_29_to_tile_9_29_1),
		.in_wire_1_2(vertical_tile_10_29_to_tile_9_29_2),
		.in_wire_1_3(vertical_tile_10_29_to_tile_9_29_3),
		.out_wire_2_0(horizontal_tile_9_29_to_tile_9_28_0),
		.out_wire_2_1(horizontal_tile_9_29_to_tile_9_28_1),
		.out_wire_2_2(horizontal_tile_9_29_to_tile_9_28_2),
		.out_wire_2_3(horizontal_tile_9_29_to_tile_9_28_3),
		.in_wire_2_0(horizontal_tile_9_28_to_tile_9_29_0),
		.in_wire_2_1(horizontal_tile_9_28_to_tile_9_29_1),
		.in_wire_2_2(horizontal_tile_9_28_to_tile_9_29_2),
		.in_wire_2_3(horizontal_tile_9_28_to_tile_9_29_3),
		.out_wire_0_0(horizontal_tile_9_29_to_tile_9_30_0),
		.out_wire_0_1(horizontal_tile_9_29_to_tile_9_30_1),
		.out_wire_0_2(horizontal_tile_9_29_to_tile_9_30_2),
		.out_wire_0_3(horizontal_tile_9_29_to_tile_9_30_3),
		.in_wire_0_0(horizontal_tile_9_30_to_tile_9_29_0),
		.in_wire_0_1(horizontal_tile_9_30_to_tile_9_29_1),
		.in_wire_0_2(horizontal_tile_9_30_to_tile_9_29_2),
		.in_wire_0_3(horizontal_tile_9_30_to_tile_9_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(318)
	);

	pe_tile pe_tile_9_30(
		.out_wire_3_0(vertical_tile_9_30_to_tile_8_30_0),
		.out_wire_3_1(vertical_tile_9_30_to_tile_8_30_1),
		.out_wire_3_2(vertical_tile_9_30_to_tile_8_30_2),
		.out_wire_3_3(vertical_tile_9_30_to_tile_8_30_3),
		.in_wire_3_0(vertical_tile_8_30_to_tile_9_30_0),
		.in_wire_3_1(vertical_tile_8_30_to_tile_9_30_1),
		.in_wire_3_2(vertical_tile_8_30_to_tile_9_30_2),
		.in_wire_3_3(vertical_tile_8_30_to_tile_9_30_3),
		.out_wire_1_0(vertical_tile_9_30_to_tile_10_30_0),
		.out_wire_1_1(vertical_tile_9_30_to_tile_10_30_1),
		.out_wire_1_2(vertical_tile_9_30_to_tile_10_30_2),
		.out_wire_1_3(vertical_tile_9_30_to_tile_10_30_3),
		.in_wire_1_0(vertical_tile_10_30_to_tile_9_30_0),
		.in_wire_1_1(vertical_tile_10_30_to_tile_9_30_1),
		.in_wire_1_2(vertical_tile_10_30_to_tile_9_30_2),
		.in_wire_1_3(vertical_tile_10_30_to_tile_9_30_3),
		.out_wire_2_0(horizontal_tile_9_30_to_tile_9_29_0),
		.out_wire_2_1(horizontal_tile_9_30_to_tile_9_29_1),
		.out_wire_2_2(horizontal_tile_9_30_to_tile_9_29_2),
		.out_wire_2_3(horizontal_tile_9_30_to_tile_9_29_3),
		.in_wire_2_0(horizontal_tile_9_29_to_tile_9_30_0),
		.in_wire_2_1(horizontal_tile_9_29_to_tile_9_30_1),
		.in_wire_2_2(horizontal_tile_9_29_to_tile_9_30_2),
		.in_wire_2_3(horizontal_tile_9_29_to_tile_9_30_3),
		.out_wire_0_0(horizontal_tile_9_30_to_tile_9_31_0),
		.out_wire_0_1(horizontal_tile_9_30_to_tile_9_31_1),
		.out_wire_0_2(horizontal_tile_9_30_to_tile_9_31_2),
		.out_wire_0_3(horizontal_tile_9_30_to_tile_9_31_3),
		.in_wire_0_0(horizontal_tile_9_31_to_tile_9_30_0),
		.in_wire_0_1(horizontal_tile_9_31_to_tile_9_30_1),
		.in_wire_0_2(horizontal_tile_9_31_to_tile_9_30_2),
		.in_wire_0_3(horizontal_tile_9_31_to_tile_9_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(319)
	);

	pe_tile_right pe_tile_9_31(
		.out_wire_3_0(vertical_tile_9_31_to_tile_8_31_0),
		.out_wire_3_1(vertical_tile_9_31_to_tile_8_31_1),
		.out_wire_3_2(vertical_tile_9_31_to_tile_8_31_2),
		.out_wire_3_3(vertical_tile_9_31_to_tile_8_31_3),
		.in_wire_3_0(vertical_tile_8_31_to_tile_9_31_0),
		.in_wire_3_1(vertical_tile_8_31_to_tile_9_31_1),
		.in_wire_3_2(vertical_tile_8_31_to_tile_9_31_2),
		.in_wire_3_3(vertical_tile_8_31_to_tile_9_31_3),
		.out_wire_1_0(vertical_tile_9_31_to_tile_10_31_0),
		.out_wire_1_1(vertical_tile_9_31_to_tile_10_31_1),
		.out_wire_1_2(vertical_tile_9_31_to_tile_10_31_2),
		.out_wire_1_3(vertical_tile_9_31_to_tile_10_31_3),
		.in_wire_1_0(vertical_tile_10_31_to_tile_9_31_0),
		.in_wire_1_1(vertical_tile_10_31_to_tile_9_31_1),
		.in_wire_1_2(vertical_tile_10_31_to_tile_9_31_2),
		.in_wire_1_3(vertical_tile_10_31_to_tile_9_31_3),
		.out_wire_2_0(horizontal_tile_9_31_to_tile_9_30_0),
		.out_wire_2_1(horizontal_tile_9_31_to_tile_9_30_1),
		.out_wire_2_2(horizontal_tile_9_31_to_tile_9_30_2),
		.out_wire_2_3(horizontal_tile_9_31_to_tile_9_30_3),
		.in_wire_2_0(horizontal_tile_9_30_to_tile_9_31_0),
		.in_wire_2_1(horizontal_tile_9_30_to_tile_9_31_1),
		.in_wire_2_2(horizontal_tile_9_30_to_tile_9_31_2),
		.in_wire_2_3(horizontal_tile_9_30_to_tile_9_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(320)
	);

	pe_tile_left pe_tile_10_0(
		.out_wire_3_0(vertical_tile_10_0_to_tile_9_0_0),
		.out_wire_3_1(vertical_tile_10_0_to_tile_9_0_1),
		.out_wire_3_2(vertical_tile_10_0_to_tile_9_0_2),
		.out_wire_3_3(vertical_tile_10_0_to_tile_9_0_3),
		.in_wire_3_0(vertical_tile_9_0_to_tile_10_0_0),
		.in_wire_3_1(vertical_tile_9_0_to_tile_10_0_1),
		.in_wire_3_2(vertical_tile_9_0_to_tile_10_0_2),
		.in_wire_3_3(vertical_tile_9_0_to_tile_10_0_3),
		.out_wire_1_0(vertical_tile_10_0_to_tile_11_0_0),
		.out_wire_1_1(vertical_tile_10_0_to_tile_11_0_1),
		.out_wire_1_2(vertical_tile_10_0_to_tile_11_0_2),
		.out_wire_1_3(vertical_tile_10_0_to_tile_11_0_3),
		.in_wire_1_0(vertical_tile_11_0_to_tile_10_0_0),
		.in_wire_1_1(vertical_tile_11_0_to_tile_10_0_1),
		.in_wire_1_2(vertical_tile_11_0_to_tile_10_0_2),
		.in_wire_1_3(vertical_tile_11_0_to_tile_10_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_10_0_to_tile_10_1_0),
		.out_wire_0_1(horizontal_tile_10_0_to_tile_10_1_1),
		.out_wire_0_2(horizontal_tile_10_0_to_tile_10_1_2),
		.out_wire_0_3(horizontal_tile_10_0_to_tile_10_1_3),
		.in_wire_0_0(horizontal_tile_10_1_to_tile_10_0_0),
		.in_wire_0_1(horizontal_tile_10_1_to_tile_10_0_1),
		.in_wire_0_2(horizontal_tile_10_1_to_tile_10_0_2),
		.in_wire_0_3(horizontal_tile_10_1_to_tile_10_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(321)
	);

	pe_tile pe_tile_10_1(
		.out_wire_3_0(vertical_tile_10_1_to_tile_9_1_0),
		.out_wire_3_1(vertical_tile_10_1_to_tile_9_1_1),
		.out_wire_3_2(vertical_tile_10_1_to_tile_9_1_2),
		.out_wire_3_3(vertical_tile_10_1_to_tile_9_1_3),
		.in_wire_3_0(vertical_tile_9_1_to_tile_10_1_0),
		.in_wire_3_1(vertical_tile_9_1_to_tile_10_1_1),
		.in_wire_3_2(vertical_tile_9_1_to_tile_10_1_2),
		.in_wire_3_3(vertical_tile_9_1_to_tile_10_1_3),
		.out_wire_1_0(vertical_tile_10_1_to_tile_11_1_0),
		.out_wire_1_1(vertical_tile_10_1_to_tile_11_1_1),
		.out_wire_1_2(vertical_tile_10_1_to_tile_11_1_2),
		.out_wire_1_3(vertical_tile_10_1_to_tile_11_1_3),
		.in_wire_1_0(vertical_tile_11_1_to_tile_10_1_0),
		.in_wire_1_1(vertical_tile_11_1_to_tile_10_1_1),
		.in_wire_1_2(vertical_tile_11_1_to_tile_10_1_2),
		.in_wire_1_3(vertical_tile_11_1_to_tile_10_1_3),
		.out_wire_2_0(horizontal_tile_10_1_to_tile_10_0_0),
		.out_wire_2_1(horizontal_tile_10_1_to_tile_10_0_1),
		.out_wire_2_2(horizontal_tile_10_1_to_tile_10_0_2),
		.out_wire_2_3(horizontal_tile_10_1_to_tile_10_0_3),
		.in_wire_2_0(horizontal_tile_10_0_to_tile_10_1_0),
		.in_wire_2_1(horizontal_tile_10_0_to_tile_10_1_1),
		.in_wire_2_2(horizontal_tile_10_0_to_tile_10_1_2),
		.in_wire_2_3(horizontal_tile_10_0_to_tile_10_1_3),
		.out_wire_0_0(horizontal_tile_10_1_to_tile_10_2_0),
		.out_wire_0_1(horizontal_tile_10_1_to_tile_10_2_1),
		.out_wire_0_2(horizontal_tile_10_1_to_tile_10_2_2),
		.out_wire_0_3(horizontal_tile_10_1_to_tile_10_2_3),
		.in_wire_0_0(horizontal_tile_10_2_to_tile_10_1_0),
		.in_wire_0_1(horizontal_tile_10_2_to_tile_10_1_1),
		.in_wire_0_2(horizontal_tile_10_2_to_tile_10_1_2),
		.in_wire_0_3(horizontal_tile_10_2_to_tile_10_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(322)
	);

	pe_tile pe_tile_10_2(
		.out_wire_3_0(vertical_tile_10_2_to_tile_9_2_0),
		.out_wire_3_1(vertical_tile_10_2_to_tile_9_2_1),
		.out_wire_3_2(vertical_tile_10_2_to_tile_9_2_2),
		.out_wire_3_3(vertical_tile_10_2_to_tile_9_2_3),
		.in_wire_3_0(vertical_tile_9_2_to_tile_10_2_0),
		.in_wire_3_1(vertical_tile_9_2_to_tile_10_2_1),
		.in_wire_3_2(vertical_tile_9_2_to_tile_10_2_2),
		.in_wire_3_3(vertical_tile_9_2_to_tile_10_2_3),
		.out_wire_1_0(vertical_tile_10_2_to_tile_11_2_0),
		.out_wire_1_1(vertical_tile_10_2_to_tile_11_2_1),
		.out_wire_1_2(vertical_tile_10_2_to_tile_11_2_2),
		.out_wire_1_3(vertical_tile_10_2_to_tile_11_2_3),
		.in_wire_1_0(vertical_tile_11_2_to_tile_10_2_0),
		.in_wire_1_1(vertical_tile_11_2_to_tile_10_2_1),
		.in_wire_1_2(vertical_tile_11_2_to_tile_10_2_2),
		.in_wire_1_3(vertical_tile_11_2_to_tile_10_2_3),
		.out_wire_2_0(horizontal_tile_10_2_to_tile_10_1_0),
		.out_wire_2_1(horizontal_tile_10_2_to_tile_10_1_1),
		.out_wire_2_2(horizontal_tile_10_2_to_tile_10_1_2),
		.out_wire_2_3(horizontal_tile_10_2_to_tile_10_1_3),
		.in_wire_2_0(horizontal_tile_10_1_to_tile_10_2_0),
		.in_wire_2_1(horizontal_tile_10_1_to_tile_10_2_1),
		.in_wire_2_2(horizontal_tile_10_1_to_tile_10_2_2),
		.in_wire_2_3(horizontal_tile_10_1_to_tile_10_2_3),
		.out_wire_0_0(horizontal_tile_10_2_to_tile_10_3_0),
		.out_wire_0_1(horizontal_tile_10_2_to_tile_10_3_1),
		.out_wire_0_2(horizontal_tile_10_2_to_tile_10_3_2),
		.out_wire_0_3(horizontal_tile_10_2_to_tile_10_3_3),
		.in_wire_0_0(horizontal_tile_10_3_to_tile_10_2_0),
		.in_wire_0_1(horizontal_tile_10_3_to_tile_10_2_1),
		.in_wire_0_2(horizontal_tile_10_3_to_tile_10_2_2),
		.in_wire_0_3(horizontal_tile_10_3_to_tile_10_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(323)
	);

	pe_tile pe_tile_10_3(
		.out_wire_3_0(vertical_tile_10_3_to_tile_9_3_0),
		.out_wire_3_1(vertical_tile_10_3_to_tile_9_3_1),
		.out_wire_3_2(vertical_tile_10_3_to_tile_9_3_2),
		.out_wire_3_3(vertical_tile_10_3_to_tile_9_3_3),
		.in_wire_3_0(vertical_tile_9_3_to_tile_10_3_0),
		.in_wire_3_1(vertical_tile_9_3_to_tile_10_3_1),
		.in_wire_3_2(vertical_tile_9_3_to_tile_10_3_2),
		.in_wire_3_3(vertical_tile_9_3_to_tile_10_3_3),
		.out_wire_1_0(vertical_tile_10_3_to_tile_11_3_0),
		.out_wire_1_1(vertical_tile_10_3_to_tile_11_3_1),
		.out_wire_1_2(vertical_tile_10_3_to_tile_11_3_2),
		.out_wire_1_3(vertical_tile_10_3_to_tile_11_3_3),
		.in_wire_1_0(vertical_tile_11_3_to_tile_10_3_0),
		.in_wire_1_1(vertical_tile_11_3_to_tile_10_3_1),
		.in_wire_1_2(vertical_tile_11_3_to_tile_10_3_2),
		.in_wire_1_3(vertical_tile_11_3_to_tile_10_3_3),
		.out_wire_2_0(horizontal_tile_10_3_to_tile_10_2_0),
		.out_wire_2_1(horizontal_tile_10_3_to_tile_10_2_1),
		.out_wire_2_2(horizontal_tile_10_3_to_tile_10_2_2),
		.out_wire_2_3(horizontal_tile_10_3_to_tile_10_2_3),
		.in_wire_2_0(horizontal_tile_10_2_to_tile_10_3_0),
		.in_wire_2_1(horizontal_tile_10_2_to_tile_10_3_1),
		.in_wire_2_2(horizontal_tile_10_2_to_tile_10_3_2),
		.in_wire_2_3(horizontal_tile_10_2_to_tile_10_3_3),
		.out_wire_0_0(horizontal_tile_10_3_to_tile_10_4_0),
		.out_wire_0_1(horizontal_tile_10_3_to_tile_10_4_1),
		.out_wire_0_2(horizontal_tile_10_3_to_tile_10_4_2),
		.out_wire_0_3(horizontal_tile_10_3_to_tile_10_4_3),
		.in_wire_0_0(horizontal_tile_10_4_to_tile_10_3_0),
		.in_wire_0_1(horizontal_tile_10_4_to_tile_10_3_1),
		.in_wire_0_2(horizontal_tile_10_4_to_tile_10_3_2),
		.in_wire_0_3(horizontal_tile_10_4_to_tile_10_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(324)
	);

	pe_tile pe_tile_10_4(
		.out_wire_3_0(vertical_tile_10_4_to_tile_9_4_0),
		.out_wire_3_1(vertical_tile_10_4_to_tile_9_4_1),
		.out_wire_3_2(vertical_tile_10_4_to_tile_9_4_2),
		.out_wire_3_3(vertical_tile_10_4_to_tile_9_4_3),
		.in_wire_3_0(vertical_tile_9_4_to_tile_10_4_0),
		.in_wire_3_1(vertical_tile_9_4_to_tile_10_4_1),
		.in_wire_3_2(vertical_tile_9_4_to_tile_10_4_2),
		.in_wire_3_3(vertical_tile_9_4_to_tile_10_4_3),
		.out_wire_1_0(vertical_tile_10_4_to_tile_11_4_0),
		.out_wire_1_1(vertical_tile_10_4_to_tile_11_4_1),
		.out_wire_1_2(vertical_tile_10_4_to_tile_11_4_2),
		.out_wire_1_3(vertical_tile_10_4_to_tile_11_4_3),
		.in_wire_1_0(vertical_tile_11_4_to_tile_10_4_0),
		.in_wire_1_1(vertical_tile_11_4_to_tile_10_4_1),
		.in_wire_1_2(vertical_tile_11_4_to_tile_10_4_2),
		.in_wire_1_3(vertical_tile_11_4_to_tile_10_4_3),
		.out_wire_2_0(horizontal_tile_10_4_to_tile_10_3_0),
		.out_wire_2_1(horizontal_tile_10_4_to_tile_10_3_1),
		.out_wire_2_2(horizontal_tile_10_4_to_tile_10_3_2),
		.out_wire_2_3(horizontal_tile_10_4_to_tile_10_3_3),
		.in_wire_2_0(horizontal_tile_10_3_to_tile_10_4_0),
		.in_wire_2_1(horizontal_tile_10_3_to_tile_10_4_1),
		.in_wire_2_2(horizontal_tile_10_3_to_tile_10_4_2),
		.in_wire_2_3(horizontal_tile_10_3_to_tile_10_4_3),
		.out_wire_0_0(horizontal_tile_10_4_to_tile_10_5_0),
		.out_wire_0_1(horizontal_tile_10_4_to_tile_10_5_1),
		.out_wire_0_2(horizontal_tile_10_4_to_tile_10_5_2),
		.out_wire_0_3(horizontal_tile_10_4_to_tile_10_5_3),
		.in_wire_0_0(horizontal_tile_10_5_to_tile_10_4_0),
		.in_wire_0_1(horizontal_tile_10_5_to_tile_10_4_1),
		.in_wire_0_2(horizontal_tile_10_5_to_tile_10_4_2),
		.in_wire_0_3(horizontal_tile_10_5_to_tile_10_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(325)
	);

	pe_tile pe_tile_10_5(
		.out_wire_3_0(vertical_tile_10_5_to_tile_9_5_0),
		.out_wire_3_1(vertical_tile_10_5_to_tile_9_5_1),
		.out_wire_3_2(vertical_tile_10_5_to_tile_9_5_2),
		.out_wire_3_3(vertical_tile_10_5_to_tile_9_5_3),
		.in_wire_3_0(vertical_tile_9_5_to_tile_10_5_0),
		.in_wire_3_1(vertical_tile_9_5_to_tile_10_5_1),
		.in_wire_3_2(vertical_tile_9_5_to_tile_10_5_2),
		.in_wire_3_3(vertical_tile_9_5_to_tile_10_5_3),
		.out_wire_1_0(vertical_tile_10_5_to_tile_11_5_0),
		.out_wire_1_1(vertical_tile_10_5_to_tile_11_5_1),
		.out_wire_1_2(vertical_tile_10_5_to_tile_11_5_2),
		.out_wire_1_3(vertical_tile_10_5_to_tile_11_5_3),
		.in_wire_1_0(vertical_tile_11_5_to_tile_10_5_0),
		.in_wire_1_1(vertical_tile_11_5_to_tile_10_5_1),
		.in_wire_1_2(vertical_tile_11_5_to_tile_10_5_2),
		.in_wire_1_3(vertical_tile_11_5_to_tile_10_5_3),
		.out_wire_2_0(horizontal_tile_10_5_to_tile_10_4_0),
		.out_wire_2_1(horizontal_tile_10_5_to_tile_10_4_1),
		.out_wire_2_2(horizontal_tile_10_5_to_tile_10_4_2),
		.out_wire_2_3(horizontal_tile_10_5_to_tile_10_4_3),
		.in_wire_2_0(horizontal_tile_10_4_to_tile_10_5_0),
		.in_wire_2_1(horizontal_tile_10_4_to_tile_10_5_1),
		.in_wire_2_2(horizontal_tile_10_4_to_tile_10_5_2),
		.in_wire_2_3(horizontal_tile_10_4_to_tile_10_5_3),
		.out_wire_0_0(horizontal_tile_10_5_to_tile_10_6_0),
		.out_wire_0_1(horizontal_tile_10_5_to_tile_10_6_1),
		.out_wire_0_2(horizontal_tile_10_5_to_tile_10_6_2),
		.out_wire_0_3(horizontal_tile_10_5_to_tile_10_6_3),
		.in_wire_0_0(horizontal_tile_10_6_to_tile_10_5_0),
		.in_wire_0_1(horizontal_tile_10_6_to_tile_10_5_1),
		.in_wire_0_2(horizontal_tile_10_6_to_tile_10_5_2),
		.in_wire_0_3(horizontal_tile_10_6_to_tile_10_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(326)
	);

	pe_tile pe_tile_10_6(
		.out_wire_3_0(vertical_tile_10_6_to_tile_9_6_0),
		.out_wire_3_1(vertical_tile_10_6_to_tile_9_6_1),
		.out_wire_3_2(vertical_tile_10_6_to_tile_9_6_2),
		.out_wire_3_3(vertical_tile_10_6_to_tile_9_6_3),
		.in_wire_3_0(vertical_tile_9_6_to_tile_10_6_0),
		.in_wire_3_1(vertical_tile_9_6_to_tile_10_6_1),
		.in_wire_3_2(vertical_tile_9_6_to_tile_10_6_2),
		.in_wire_3_3(vertical_tile_9_6_to_tile_10_6_3),
		.out_wire_1_0(vertical_tile_10_6_to_tile_11_6_0),
		.out_wire_1_1(vertical_tile_10_6_to_tile_11_6_1),
		.out_wire_1_2(vertical_tile_10_6_to_tile_11_6_2),
		.out_wire_1_3(vertical_tile_10_6_to_tile_11_6_3),
		.in_wire_1_0(vertical_tile_11_6_to_tile_10_6_0),
		.in_wire_1_1(vertical_tile_11_6_to_tile_10_6_1),
		.in_wire_1_2(vertical_tile_11_6_to_tile_10_6_2),
		.in_wire_1_3(vertical_tile_11_6_to_tile_10_6_3),
		.out_wire_2_0(horizontal_tile_10_6_to_tile_10_5_0),
		.out_wire_2_1(horizontal_tile_10_6_to_tile_10_5_1),
		.out_wire_2_2(horizontal_tile_10_6_to_tile_10_5_2),
		.out_wire_2_3(horizontal_tile_10_6_to_tile_10_5_3),
		.in_wire_2_0(horizontal_tile_10_5_to_tile_10_6_0),
		.in_wire_2_1(horizontal_tile_10_5_to_tile_10_6_1),
		.in_wire_2_2(horizontal_tile_10_5_to_tile_10_6_2),
		.in_wire_2_3(horizontal_tile_10_5_to_tile_10_6_3),
		.out_wire_0_0(horizontal_tile_10_6_to_tile_10_7_0),
		.out_wire_0_1(horizontal_tile_10_6_to_tile_10_7_1),
		.out_wire_0_2(horizontal_tile_10_6_to_tile_10_7_2),
		.out_wire_0_3(horizontal_tile_10_6_to_tile_10_7_3),
		.in_wire_0_0(horizontal_tile_10_7_to_tile_10_6_0),
		.in_wire_0_1(horizontal_tile_10_7_to_tile_10_6_1),
		.in_wire_0_2(horizontal_tile_10_7_to_tile_10_6_2),
		.in_wire_0_3(horizontal_tile_10_7_to_tile_10_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(327)
	);

	pe_tile pe_tile_10_7(
		.out_wire_3_0(vertical_tile_10_7_to_tile_9_7_0),
		.out_wire_3_1(vertical_tile_10_7_to_tile_9_7_1),
		.out_wire_3_2(vertical_tile_10_7_to_tile_9_7_2),
		.out_wire_3_3(vertical_tile_10_7_to_tile_9_7_3),
		.in_wire_3_0(vertical_tile_9_7_to_tile_10_7_0),
		.in_wire_3_1(vertical_tile_9_7_to_tile_10_7_1),
		.in_wire_3_2(vertical_tile_9_7_to_tile_10_7_2),
		.in_wire_3_3(vertical_tile_9_7_to_tile_10_7_3),
		.out_wire_1_0(vertical_tile_10_7_to_tile_11_7_0),
		.out_wire_1_1(vertical_tile_10_7_to_tile_11_7_1),
		.out_wire_1_2(vertical_tile_10_7_to_tile_11_7_2),
		.out_wire_1_3(vertical_tile_10_7_to_tile_11_7_3),
		.in_wire_1_0(vertical_tile_11_7_to_tile_10_7_0),
		.in_wire_1_1(vertical_tile_11_7_to_tile_10_7_1),
		.in_wire_1_2(vertical_tile_11_7_to_tile_10_7_2),
		.in_wire_1_3(vertical_tile_11_7_to_tile_10_7_3),
		.out_wire_2_0(horizontal_tile_10_7_to_tile_10_6_0),
		.out_wire_2_1(horizontal_tile_10_7_to_tile_10_6_1),
		.out_wire_2_2(horizontal_tile_10_7_to_tile_10_6_2),
		.out_wire_2_3(horizontal_tile_10_7_to_tile_10_6_3),
		.in_wire_2_0(horizontal_tile_10_6_to_tile_10_7_0),
		.in_wire_2_1(horizontal_tile_10_6_to_tile_10_7_1),
		.in_wire_2_2(horizontal_tile_10_6_to_tile_10_7_2),
		.in_wire_2_3(horizontal_tile_10_6_to_tile_10_7_3),
		.out_wire_0_0(horizontal_tile_10_7_to_tile_10_8_0),
		.out_wire_0_1(horizontal_tile_10_7_to_tile_10_8_1),
		.out_wire_0_2(horizontal_tile_10_7_to_tile_10_8_2),
		.out_wire_0_3(horizontal_tile_10_7_to_tile_10_8_3),
		.in_wire_0_0(horizontal_tile_10_8_to_tile_10_7_0),
		.in_wire_0_1(horizontal_tile_10_8_to_tile_10_7_1),
		.in_wire_0_2(horizontal_tile_10_8_to_tile_10_7_2),
		.in_wire_0_3(horizontal_tile_10_8_to_tile_10_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(328)
	);

	pe_tile pe_tile_10_8(
		.out_wire_3_0(vertical_tile_10_8_to_tile_9_8_0),
		.out_wire_3_1(vertical_tile_10_8_to_tile_9_8_1),
		.out_wire_3_2(vertical_tile_10_8_to_tile_9_8_2),
		.out_wire_3_3(vertical_tile_10_8_to_tile_9_8_3),
		.in_wire_3_0(vertical_tile_9_8_to_tile_10_8_0),
		.in_wire_3_1(vertical_tile_9_8_to_tile_10_8_1),
		.in_wire_3_2(vertical_tile_9_8_to_tile_10_8_2),
		.in_wire_3_3(vertical_tile_9_8_to_tile_10_8_3),
		.out_wire_1_0(vertical_tile_10_8_to_tile_11_8_0),
		.out_wire_1_1(vertical_tile_10_8_to_tile_11_8_1),
		.out_wire_1_2(vertical_tile_10_8_to_tile_11_8_2),
		.out_wire_1_3(vertical_tile_10_8_to_tile_11_8_3),
		.in_wire_1_0(vertical_tile_11_8_to_tile_10_8_0),
		.in_wire_1_1(vertical_tile_11_8_to_tile_10_8_1),
		.in_wire_1_2(vertical_tile_11_8_to_tile_10_8_2),
		.in_wire_1_3(vertical_tile_11_8_to_tile_10_8_3),
		.out_wire_2_0(horizontal_tile_10_8_to_tile_10_7_0),
		.out_wire_2_1(horizontal_tile_10_8_to_tile_10_7_1),
		.out_wire_2_2(horizontal_tile_10_8_to_tile_10_7_2),
		.out_wire_2_3(horizontal_tile_10_8_to_tile_10_7_3),
		.in_wire_2_0(horizontal_tile_10_7_to_tile_10_8_0),
		.in_wire_2_1(horizontal_tile_10_7_to_tile_10_8_1),
		.in_wire_2_2(horizontal_tile_10_7_to_tile_10_8_2),
		.in_wire_2_3(horizontal_tile_10_7_to_tile_10_8_3),
		.out_wire_0_0(horizontal_tile_10_8_to_tile_10_9_0),
		.out_wire_0_1(horizontal_tile_10_8_to_tile_10_9_1),
		.out_wire_0_2(horizontal_tile_10_8_to_tile_10_9_2),
		.out_wire_0_3(horizontal_tile_10_8_to_tile_10_9_3),
		.in_wire_0_0(horizontal_tile_10_9_to_tile_10_8_0),
		.in_wire_0_1(horizontal_tile_10_9_to_tile_10_8_1),
		.in_wire_0_2(horizontal_tile_10_9_to_tile_10_8_2),
		.in_wire_0_3(horizontal_tile_10_9_to_tile_10_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(329)
	);

	pe_tile pe_tile_10_9(
		.out_wire_3_0(vertical_tile_10_9_to_tile_9_9_0),
		.out_wire_3_1(vertical_tile_10_9_to_tile_9_9_1),
		.out_wire_3_2(vertical_tile_10_9_to_tile_9_9_2),
		.out_wire_3_3(vertical_tile_10_9_to_tile_9_9_3),
		.in_wire_3_0(vertical_tile_9_9_to_tile_10_9_0),
		.in_wire_3_1(vertical_tile_9_9_to_tile_10_9_1),
		.in_wire_3_2(vertical_tile_9_9_to_tile_10_9_2),
		.in_wire_3_3(vertical_tile_9_9_to_tile_10_9_3),
		.out_wire_1_0(vertical_tile_10_9_to_tile_11_9_0),
		.out_wire_1_1(vertical_tile_10_9_to_tile_11_9_1),
		.out_wire_1_2(vertical_tile_10_9_to_tile_11_9_2),
		.out_wire_1_3(vertical_tile_10_9_to_tile_11_9_3),
		.in_wire_1_0(vertical_tile_11_9_to_tile_10_9_0),
		.in_wire_1_1(vertical_tile_11_9_to_tile_10_9_1),
		.in_wire_1_2(vertical_tile_11_9_to_tile_10_9_2),
		.in_wire_1_3(vertical_tile_11_9_to_tile_10_9_3),
		.out_wire_2_0(horizontal_tile_10_9_to_tile_10_8_0),
		.out_wire_2_1(horizontal_tile_10_9_to_tile_10_8_1),
		.out_wire_2_2(horizontal_tile_10_9_to_tile_10_8_2),
		.out_wire_2_3(horizontal_tile_10_9_to_tile_10_8_3),
		.in_wire_2_0(horizontal_tile_10_8_to_tile_10_9_0),
		.in_wire_2_1(horizontal_tile_10_8_to_tile_10_9_1),
		.in_wire_2_2(horizontal_tile_10_8_to_tile_10_9_2),
		.in_wire_2_3(horizontal_tile_10_8_to_tile_10_9_3),
		.out_wire_0_0(horizontal_tile_10_9_to_tile_10_10_0),
		.out_wire_0_1(horizontal_tile_10_9_to_tile_10_10_1),
		.out_wire_0_2(horizontal_tile_10_9_to_tile_10_10_2),
		.out_wire_0_3(horizontal_tile_10_9_to_tile_10_10_3),
		.in_wire_0_0(horizontal_tile_10_10_to_tile_10_9_0),
		.in_wire_0_1(horizontal_tile_10_10_to_tile_10_9_1),
		.in_wire_0_2(horizontal_tile_10_10_to_tile_10_9_2),
		.in_wire_0_3(horizontal_tile_10_10_to_tile_10_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(330)
	);

	pe_tile pe_tile_10_10(
		.out_wire_3_0(vertical_tile_10_10_to_tile_9_10_0),
		.out_wire_3_1(vertical_tile_10_10_to_tile_9_10_1),
		.out_wire_3_2(vertical_tile_10_10_to_tile_9_10_2),
		.out_wire_3_3(vertical_tile_10_10_to_tile_9_10_3),
		.in_wire_3_0(vertical_tile_9_10_to_tile_10_10_0),
		.in_wire_3_1(vertical_tile_9_10_to_tile_10_10_1),
		.in_wire_3_2(vertical_tile_9_10_to_tile_10_10_2),
		.in_wire_3_3(vertical_tile_9_10_to_tile_10_10_3),
		.out_wire_1_0(vertical_tile_10_10_to_tile_11_10_0),
		.out_wire_1_1(vertical_tile_10_10_to_tile_11_10_1),
		.out_wire_1_2(vertical_tile_10_10_to_tile_11_10_2),
		.out_wire_1_3(vertical_tile_10_10_to_tile_11_10_3),
		.in_wire_1_0(vertical_tile_11_10_to_tile_10_10_0),
		.in_wire_1_1(vertical_tile_11_10_to_tile_10_10_1),
		.in_wire_1_2(vertical_tile_11_10_to_tile_10_10_2),
		.in_wire_1_3(vertical_tile_11_10_to_tile_10_10_3),
		.out_wire_2_0(horizontal_tile_10_10_to_tile_10_9_0),
		.out_wire_2_1(horizontal_tile_10_10_to_tile_10_9_1),
		.out_wire_2_2(horizontal_tile_10_10_to_tile_10_9_2),
		.out_wire_2_3(horizontal_tile_10_10_to_tile_10_9_3),
		.in_wire_2_0(horizontal_tile_10_9_to_tile_10_10_0),
		.in_wire_2_1(horizontal_tile_10_9_to_tile_10_10_1),
		.in_wire_2_2(horizontal_tile_10_9_to_tile_10_10_2),
		.in_wire_2_3(horizontal_tile_10_9_to_tile_10_10_3),
		.out_wire_0_0(horizontal_tile_10_10_to_tile_10_11_0),
		.out_wire_0_1(horizontal_tile_10_10_to_tile_10_11_1),
		.out_wire_0_2(horizontal_tile_10_10_to_tile_10_11_2),
		.out_wire_0_3(horizontal_tile_10_10_to_tile_10_11_3),
		.in_wire_0_0(horizontal_tile_10_11_to_tile_10_10_0),
		.in_wire_0_1(horizontal_tile_10_11_to_tile_10_10_1),
		.in_wire_0_2(horizontal_tile_10_11_to_tile_10_10_2),
		.in_wire_0_3(horizontal_tile_10_11_to_tile_10_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(331)
	);

	pe_tile pe_tile_10_11(
		.out_wire_3_0(vertical_tile_10_11_to_tile_9_11_0),
		.out_wire_3_1(vertical_tile_10_11_to_tile_9_11_1),
		.out_wire_3_2(vertical_tile_10_11_to_tile_9_11_2),
		.out_wire_3_3(vertical_tile_10_11_to_tile_9_11_3),
		.in_wire_3_0(vertical_tile_9_11_to_tile_10_11_0),
		.in_wire_3_1(vertical_tile_9_11_to_tile_10_11_1),
		.in_wire_3_2(vertical_tile_9_11_to_tile_10_11_2),
		.in_wire_3_3(vertical_tile_9_11_to_tile_10_11_3),
		.out_wire_1_0(vertical_tile_10_11_to_tile_11_11_0),
		.out_wire_1_1(vertical_tile_10_11_to_tile_11_11_1),
		.out_wire_1_2(vertical_tile_10_11_to_tile_11_11_2),
		.out_wire_1_3(vertical_tile_10_11_to_tile_11_11_3),
		.in_wire_1_0(vertical_tile_11_11_to_tile_10_11_0),
		.in_wire_1_1(vertical_tile_11_11_to_tile_10_11_1),
		.in_wire_1_2(vertical_tile_11_11_to_tile_10_11_2),
		.in_wire_1_3(vertical_tile_11_11_to_tile_10_11_3),
		.out_wire_2_0(horizontal_tile_10_11_to_tile_10_10_0),
		.out_wire_2_1(horizontal_tile_10_11_to_tile_10_10_1),
		.out_wire_2_2(horizontal_tile_10_11_to_tile_10_10_2),
		.out_wire_2_3(horizontal_tile_10_11_to_tile_10_10_3),
		.in_wire_2_0(horizontal_tile_10_10_to_tile_10_11_0),
		.in_wire_2_1(horizontal_tile_10_10_to_tile_10_11_1),
		.in_wire_2_2(horizontal_tile_10_10_to_tile_10_11_2),
		.in_wire_2_3(horizontal_tile_10_10_to_tile_10_11_3),
		.out_wire_0_0(horizontal_tile_10_11_to_tile_10_12_0),
		.out_wire_0_1(horizontal_tile_10_11_to_tile_10_12_1),
		.out_wire_0_2(horizontal_tile_10_11_to_tile_10_12_2),
		.out_wire_0_3(horizontal_tile_10_11_to_tile_10_12_3),
		.in_wire_0_0(horizontal_tile_10_12_to_tile_10_11_0),
		.in_wire_0_1(horizontal_tile_10_12_to_tile_10_11_1),
		.in_wire_0_2(horizontal_tile_10_12_to_tile_10_11_2),
		.in_wire_0_3(horizontal_tile_10_12_to_tile_10_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(332)
	);

	pe_tile pe_tile_10_12(
		.out_wire_3_0(vertical_tile_10_12_to_tile_9_12_0),
		.out_wire_3_1(vertical_tile_10_12_to_tile_9_12_1),
		.out_wire_3_2(vertical_tile_10_12_to_tile_9_12_2),
		.out_wire_3_3(vertical_tile_10_12_to_tile_9_12_3),
		.in_wire_3_0(vertical_tile_9_12_to_tile_10_12_0),
		.in_wire_3_1(vertical_tile_9_12_to_tile_10_12_1),
		.in_wire_3_2(vertical_tile_9_12_to_tile_10_12_2),
		.in_wire_3_3(vertical_tile_9_12_to_tile_10_12_3),
		.out_wire_1_0(vertical_tile_10_12_to_tile_11_12_0),
		.out_wire_1_1(vertical_tile_10_12_to_tile_11_12_1),
		.out_wire_1_2(vertical_tile_10_12_to_tile_11_12_2),
		.out_wire_1_3(vertical_tile_10_12_to_tile_11_12_3),
		.in_wire_1_0(vertical_tile_11_12_to_tile_10_12_0),
		.in_wire_1_1(vertical_tile_11_12_to_tile_10_12_1),
		.in_wire_1_2(vertical_tile_11_12_to_tile_10_12_2),
		.in_wire_1_3(vertical_tile_11_12_to_tile_10_12_3),
		.out_wire_2_0(horizontal_tile_10_12_to_tile_10_11_0),
		.out_wire_2_1(horizontal_tile_10_12_to_tile_10_11_1),
		.out_wire_2_2(horizontal_tile_10_12_to_tile_10_11_2),
		.out_wire_2_3(horizontal_tile_10_12_to_tile_10_11_3),
		.in_wire_2_0(horizontal_tile_10_11_to_tile_10_12_0),
		.in_wire_2_1(horizontal_tile_10_11_to_tile_10_12_1),
		.in_wire_2_2(horizontal_tile_10_11_to_tile_10_12_2),
		.in_wire_2_3(horizontal_tile_10_11_to_tile_10_12_3),
		.out_wire_0_0(horizontal_tile_10_12_to_tile_10_13_0),
		.out_wire_0_1(horizontal_tile_10_12_to_tile_10_13_1),
		.out_wire_0_2(horizontal_tile_10_12_to_tile_10_13_2),
		.out_wire_0_3(horizontal_tile_10_12_to_tile_10_13_3),
		.in_wire_0_0(horizontal_tile_10_13_to_tile_10_12_0),
		.in_wire_0_1(horizontal_tile_10_13_to_tile_10_12_1),
		.in_wire_0_2(horizontal_tile_10_13_to_tile_10_12_2),
		.in_wire_0_3(horizontal_tile_10_13_to_tile_10_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(333)
	);

	pe_tile pe_tile_10_13(
		.out_wire_3_0(vertical_tile_10_13_to_tile_9_13_0),
		.out_wire_3_1(vertical_tile_10_13_to_tile_9_13_1),
		.out_wire_3_2(vertical_tile_10_13_to_tile_9_13_2),
		.out_wire_3_3(vertical_tile_10_13_to_tile_9_13_3),
		.in_wire_3_0(vertical_tile_9_13_to_tile_10_13_0),
		.in_wire_3_1(vertical_tile_9_13_to_tile_10_13_1),
		.in_wire_3_2(vertical_tile_9_13_to_tile_10_13_2),
		.in_wire_3_3(vertical_tile_9_13_to_tile_10_13_3),
		.out_wire_1_0(vertical_tile_10_13_to_tile_11_13_0),
		.out_wire_1_1(vertical_tile_10_13_to_tile_11_13_1),
		.out_wire_1_2(vertical_tile_10_13_to_tile_11_13_2),
		.out_wire_1_3(vertical_tile_10_13_to_tile_11_13_3),
		.in_wire_1_0(vertical_tile_11_13_to_tile_10_13_0),
		.in_wire_1_1(vertical_tile_11_13_to_tile_10_13_1),
		.in_wire_1_2(vertical_tile_11_13_to_tile_10_13_2),
		.in_wire_1_3(vertical_tile_11_13_to_tile_10_13_3),
		.out_wire_2_0(horizontal_tile_10_13_to_tile_10_12_0),
		.out_wire_2_1(horizontal_tile_10_13_to_tile_10_12_1),
		.out_wire_2_2(horizontal_tile_10_13_to_tile_10_12_2),
		.out_wire_2_3(horizontal_tile_10_13_to_tile_10_12_3),
		.in_wire_2_0(horizontal_tile_10_12_to_tile_10_13_0),
		.in_wire_2_1(horizontal_tile_10_12_to_tile_10_13_1),
		.in_wire_2_2(horizontal_tile_10_12_to_tile_10_13_2),
		.in_wire_2_3(horizontal_tile_10_12_to_tile_10_13_3),
		.out_wire_0_0(horizontal_tile_10_13_to_tile_10_14_0),
		.out_wire_0_1(horizontal_tile_10_13_to_tile_10_14_1),
		.out_wire_0_2(horizontal_tile_10_13_to_tile_10_14_2),
		.out_wire_0_3(horizontal_tile_10_13_to_tile_10_14_3),
		.in_wire_0_0(horizontal_tile_10_14_to_tile_10_13_0),
		.in_wire_0_1(horizontal_tile_10_14_to_tile_10_13_1),
		.in_wire_0_2(horizontal_tile_10_14_to_tile_10_13_2),
		.in_wire_0_3(horizontal_tile_10_14_to_tile_10_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(334)
	);

	pe_tile pe_tile_10_14(
		.out_wire_3_0(vertical_tile_10_14_to_tile_9_14_0),
		.out_wire_3_1(vertical_tile_10_14_to_tile_9_14_1),
		.out_wire_3_2(vertical_tile_10_14_to_tile_9_14_2),
		.out_wire_3_3(vertical_tile_10_14_to_tile_9_14_3),
		.in_wire_3_0(vertical_tile_9_14_to_tile_10_14_0),
		.in_wire_3_1(vertical_tile_9_14_to_tile_10_14_1),
		.in_wire_3_2(vertical_tile_9_14_to_tile_10_14_2),
		.in_wire_3_3(vertical_tile_9_14_to_tile_10_14_3),
		.out_wire_1_0(vertical_tile_10_14_to_tile_11_14_0),
		.out_wire_1_1(vertical_tile_10_14_to_tile_11_14_1),
		.out_wire_1_2(vertical_tile_10_14_to_tile_11_14_2),
		.out_wire_1_3(vertical_tile_10_14_to_tile_11_14_3),
		.in_wire_1_0(vertical_tile_11_14_to_tile_10_14_0),
		.in_wire_1_1(vertical_tile_11_14_to_tile_10_14_1),
		.in_wire_1_2(vertical_tile_11_14_to_tile_10_14_2),
		.in_wire_1_3(vertical_tile_11_14_to_tile_10_14_3),
		.out_wire_2_0(horizontal_tile_10_14_to_tile_10_13_0),
		.out_wire_2_1(horizontal_tile_10_14_to_tile_10_13_1),
		.out_wire_2_2(horizontal_tile_10_14_to_tile_10_13_2),
		.out_wire_2_3(horizontal_tile_10_14_to_tile_10_13_3),
		.in_wire_2_0(horizontal_tile_10_13_to_tile_10_14_0),
		.in_wire_2_1(horizontal_tile_10_13_to_tile_10_14_1),
		.in_wire_2_2(horizontal_tile_10_13_to_tile_10_14_2),
		.in_wire_2_3(horizontal_tile_10_13_to_tile_10_14_3),
		.out_wire_0_0(horizontal_tile_10_14_to_tile_10_15_0),
		.out_wire_0_1(horizontal_tile_10_14_to_tile_10_15_1),
		.out_wire_0_2(horizontal_tile_10_14_to_tile_10_15_2),
		.out_wire_0_3(horizontal_tile_10_14_to_tile_10_15_3),
		.in_wire_0_0(horizontal_tile_10_15_to_tile_10_14_0),
		.in_wire_0_1(horizontal_tile_10_15_to_tile_10_14_1),
		.in_wire_0_2(horizontal_tile_10_15_to_tile_10_14_2),
		.in_wire_0_3(horizontal_tile_10_15_to_tile_10_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(335)
	);

	pe_tile pe_tile_10_15(
		.out_wire_3_0(vertical_tile_10_15_to_tile_9_15_0),
		.out_wire_3_1(vertical_tile_10_15_to_tile_9_15_1),
		.out_wire_3_2(vertical_tile_10_15_to_tile_9_15_2),
		.out_wire_3_3(vertical_tile_10_15_to_tile_9_15_3),
		.in_wire_3_0(vertical_tile_9_15_to_tile_10_15_0),
		.in_wire_3_1(vertical_tile_9_15_to_tile_10_15_1),
		.in_wire_3_2(vertical_tile_9_15_to_tile_10_15_2),
		.in_wire_3_3(vertical_tile_9_15_to_tile_10_15_3),
		.out_wire_1_0(vertical_tile_10_15_to_tile_11_15_0),
		.out_wire_1_1(vertical_tile_10_15_to_tile_11_15_1),
		.out_wire_1_2(vertical_tile_10_15_to_tile_11_15_2),
		.out_wire_1_3(vertical_tile_10_15_to_tile_11_15_3),
		.in_wire_1_0(vertical_tile_11_15_to_tile_10_15_0),
		.in_wire_1_1(vertical_tile_11_15_to_tile_10_15_1),
		.in_wire_1_2(vertical_tile_11_15_to_tile_10_15_2),
		.in_wire_1_3(vertical_tile_11_15_to_tile_10_15_3),
		.out_wire_2_0(horizontal_tile_10_15_to_tile_10_14_0),
		.out_wire_2_1(horizontal_tile_10_15_to_tile_10_14_1),
		.out_wire_2_2(horizontal_tile_10_15_to_tile_10_14_2),
		.out_wire_2_3(horizontal_tile_10_15_to_tile_10_14_3),
		.in_wire_2_0(horizontal_tile_10_14_to_tile_10_15_0),
		.in_wire_2_1(horizontal_tile_10_14_to_tile_10_15_1),
		.in_wire_2_2(horizontal_tile_10_14_to_tile_10_15_2),
		.in_wire_2_3(horizontal_tile_10_14_to_tile_10_15_3),
		.out_wire_0_0(horizontal_tile_10_15_to_tile_10_16_0),
		.out_wire_0_1(horizontal_tile_10_15_to_tile_10_16_1),
		.out_wire_0_2(horizontal_tile_10_15_to_tile_10_16_2),
		.out_wire_0_3(horizontal_tile_10_15_to_tile_10_16_3),
		.in_wire_0_0(horizontal_tile_10_16_to_tile_10_15_0),
		.in_wire_0_1(horizontal_tile_10_16_to_tile_10_15_1),
		.in_wire_0_2(horizontal_tile_10_16_to_tile_10_15_2),
		.in_wire_0_3(horizontal_tile_10_16_to_tile_10_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(336)
	);

	pe_tile pe_tile_10_16(
		.out_wire_3_0(vertical_tile_10_16_to_tile_9_16_0),
		.out_wire_3_1(vertical_tile_10_16_to_tile_9_16_1),
		.out_wire_3_2(vertical_tile_10_16_to_tile_9_16_2),
		.out_wire_3_3(vertical_tile_10_16_to_tile_9_16_3),
		.in_wire_3_0(vertical_tile_9_16_to_tile_10_16_0),
		.in_wire_3_1(vertical_tile_9_16_to_tile_10_16_1),
		.in_wire_3_2(vertical_tile_9_16_to_tile_10_16_2),
		.in_wire_3_3(vertical_tile_9_16_to_tile_10_16_3),
		.out_wire_1_0(vertical_tile_10_16_to_tile_11_16_0),
		.out_wire_1_1(vertical_tile_10_16_to_tile_11_16_1),
		.out_wire_1_2(vertical_tile_10_16_to_tile_11_16_2),
		.out_wire_1_3(vertical_tile_10_16_to_tile_11_16_3),
		.in_wire_1_0(vertical_tile_11_16_to_tile_10_16_0),
		.in_wire_1_1(vertical_tile_11_16_to_tile_10_16_1),
		.in_wire_1_2(vertical_tile_11_16_to_tile_10_16_2),
		.in_wire_1_3(vertical_tile_11_16_to_tile_10_16_3),
		.out_wire_2_0(horizontal_tile_10_16_to_tile_10_15_0),
		.out_wire_2_1(horizontal_tile_10_16_to_tile_10_15_1),
		.out_wire_2_2(horizontal_tile_10_16_to_tile_10_15_2),
		.out_wire_2_3(horizontal_tile_10_16_to_tile_10_15_3),
		.in_wire_2_0(horizontal_tile_10_15_to_tile_10_16_0),
		.in_wire_2_1(horizontal_tile_10_15_to_tile_10_16_1),
		.in_wire_2_2(horizontal_tile_10_15_to_tile_10_16_2),
		.in_wire_2_3(horizontal_tile_10_15_to_tile_10_16_3),
		.out_wire_0_0(horizontal_tile_10_16_to_tile_10_17_0),
		.out_wire_0_1(horizontal_tile_10_16_to_tile_10_17_1),
		.out_wire_0_2(horizontal_tile_10_16_to_tile_10_17_2),
		.out_wire_0_3(horizontal_tile_10_16_to_tile_10_17_3),
		.in_wire_0_0(horizontal_tile_10_17_to_tile_10_16_0),
		.in_wire_0_1(horizontal_tile_10_17_to_tile_10_16_1),
		.in_wire_0_2(horizontal_tile_10_17_to_tile_10_16_2),
		.in_wire_0_3(horizontal_tile_10_17_to_tile_10_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(337)
	);

	pe_tile pe_tile_10_17(
		.out_wire_3_0(vertical_tile_10_17_to_tile_9_17_0),
		.out_wire_3_1(vertical_tile_10_17_to_tile_9_17_1),
		.out_wire_3_2(vertical_tile_10_17_to_tile_9_17_2),
		.out_wire_3_3(vertical_tile_10_17_to_tile_9_17_3),
		.in_wire_3_0(vertical_tile_9_17_to_tile_10_17_0),
		.in_wire_3_1(vertical_tile_9_17_to_tile_10_17_1),
		.in_wire_3_2(vertical_tile_9_17_to_tile_10_17_2),
		.in_wire_3_3(vertical_tile_9_17_to_tile_10_17_3),
		.out_wire_1_0(vertical_tile_10_17_to_tile_11_17_0),
		.out_wire_1_1(vertical_tile_10_17_to_tile_11_17_1),
		.out_wire_1_2(vertical_tile_10_17_to_tile_11_17_2),
		.out_wire_1_3(vertical_tile_10_17_to_tile_11_17_3),
		.in_wire_1_0(vertical_tile_11_17_to_tile_10_17_0),
		.in_wire_1_1(vertical_tile_11_17_to_tile_10_17_1),
		.in_wire_1_2(vertical_tile_11_17_to_tile_10_17_2),
		.in_wire_1_3(vertical_tile_11_17_to_tile_10_17_3),
		.out_wire_2_0(horizontal_tile_10_17_to_tile_10_16_0),
		.out_wire_2_1(horizontal_tile_10_17_to_tile_10_16_1),
		.out_wire_2_2(horizontal_tile_10_17_to_tile_10_16_2),
		.out_wire_2_3(horizontal_tile_10_17_to_tile_10_16_3),
		.in_wire_2_0(horizontal_tile_10_16_to_tile_10_17_0),
		.in_wire_2_1(horizontal_tile_10_16_to_tile_10_17_1),
		.in_wire_2_2(horizontal_tile_10_16_to_tile_10_17_2),
		.in_wire_2_3(horizontal_tile_10_16_to_tile_10_17_3),
		.out_wire_0_0(horizontal_tile_10_17_to_tile_10_18_0),
		.out_wire_0_1(horizontal_tile_10_17_to_tile_10_18_1),
		.out_wire_0_2(horizontal_tile_10_17_to_tile_10_18_2),
		.out_wire_0_3(horizontal_tile_10_17_to_tile_10_18_3),
		.in_wire_0_0(horizontal_tile_10_18_to_tile_10_17_0),
		.in_wire_0_1(horizontal_tile_10_18_to_tile_10_17_1),
		.in_wire_0_2(horizontal_tile_10_18_to_tile_10_17_2),
		.in_wire_0_3(horizontal_tile_10_18_to_tile_10_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(338)
	);

	pe_tile pe_tile_10_18(
		.out_wire_3_0(vertical_tile_10_18_to_tile_9_18_0),
		.out_wire_3_1(vertical_tile_10_18_to_tile_9_18_1),
		.out_wire_3_2(vertical_tile_10_18_to_tile_9_18_2),
		.out_wire_3_3(vertical_tile_10_18_to_tile_9_18_3),
		.in_wire_3_0(vertical_tile_9_18_to_tile_10_18_0),
		.in_wire_3_1(vertical_tile_9_18_to_tile_10_18_1),
		.in_wire_3_2(vertical_tile_9_18_to_tile_10_18_2),
		.in_wire_3_3(vertical_tile_9_18_to_tile_10_18_3),
		.out_wire_1_0(vertical_tile_10_18_to_tile_11_18_0),
		.out_wire_1_1(vertical_tile_10_18_to_tile_11_18_1),
		.out_wire_1_2(vertical_tile_10_18_to_tile_11_18_2),
		.out_wire_1_3(vertical_tile_10_18_to_tile_11_18_3),
		.in_wire_1_0(vertical_tile_11_18_to_tile_10_18_0),
		.in_wire_1_1(vertical_tile_11_18_to_tile_10_18_1),
		.in_wire_1_2(vertical_tile_11_18_to_tile_10_18_2),
		.in_wire_1_3(vertical_tile_11_18_to_tile_10_18_3),
		.out_wire_2_0(horizontal_tile_10_18_to_tile_10_17_0),
		.out_wire_2_1(horizontal_tile_10_18_to_tile_10_17_1),
		.out_wire_2_2(horizontal_tile_10_18_to_tile_10_17_2),
		.out_wire_2_3(horizontal_tile_10_18_to_tile_10_17_3),
		.in_wire_2_0(horizontal_tile_10_17_to_tile_10_18_0),
		.in_wire_2_1(horizontal_tile_10_17_to_tile_10_18_1),
		.in_wire_2_2(horizontal_tile_10_17_to_tile_10_18_2),
		.in_wire_2_3(horizontal_tile_10_17_to_tile_10_18_3),
		.out_wire_0_0(horizontal_tile_10_18_to_tile_10_19_0),
		.out_wire_0_1(horizontal_tile_10_18_to_tile_10_19_1),
		.out_wire_0_2(horizontal_tile_10_18_to_tile_10_19_2),
		.out_wire_0_3(horizontal_tile_10_18_to_tile_10_19_3),
		.in_wire_0_0(horizontal_tile_10_19_to_tile_10_18_0),
		.in_wire_0_1(horizontal_tile_10_19_to_tile_10_18_1),
		.in_wire_0_2(horizontal_tile_10_19_to_tile_10_18_2),
		.in_wire_0_3(horizontal_tile_10_19_to_tile_10_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(339)
	);

	pe_tile pe_tile_10_19(
		.out_wire_3_0(vertical_tile_10_19_to_tile_9_19_0),
		.out_wire_3_1(vertical_tile_10_19_to_tile_9_19_1),
		.out_wire_3_2(vertical_tile_10_19_to_tile_9_19_2),
		.out_wire_3_3(vertical_tile_10_19_to_tile_9_19_3),
		.in_wire_3_0(vertical_tile_9_19_to_tile_10_19_0),
		.in_wire_3_1(vertical_tile_9_19_to_tile_10_19_1),
		.in_wire_3_2(vertical_tile_9_19_to_tile_10_19_2),
		.in_wire_3_3(vertical_tile_9_19_to_tile_10_19_3),
		.out_wire_1_0(vertical_tile_10_19_to_tile_11_19_0),
		.out_wire_1_1(vertical_tile_10_19_to_tile_11_19_1),
		.out_wire_1_2(vertical_tile_10_19_to_tile_11_19_2),
		.out_wire_1_3(vertical_tile_10_19_to_tile_11_19_3),
		.in_wire_1_0(vertical_tile_11_19_to_tile_10_19_0),
		.in_wire_1_1(vertical_tile_11_19_to_tile_10_19_1),
		.in_wire_1_2(vertical_tile_11_19_to_tile_10_19_2),
		.in_wire_1_3(vertical_tile_11_19_to_tile_10_19_3),
		.out_wire_2_0(horizontal_tile_10_19_to_tile_10_18_0),
		.out_wire_2_1(horizontal_tile_10_19_to_tile_10_18_1),
		.out_wire_2_2(horizontal_tile_10_19_to_tile_10_18_2),
		.out_wire_2_3(horizontal_tile_10_19_to_tile_10_18_3),
		.in_wire_2_0(horizontal_tile_10_18_to_tile_10_19_0),
		.in_wire_2_1(horizontal_tile_10_18_to_tile_10_19_1),
		.in_wire_2_2(horizontal_tile_10_18_to_tile_10_19_2),
		.in_wire_2_3(horizontal_tile_10_18_to_tile_10_19_3),
		.out_wire_0_0(horizontal_tile_10_19_to_tile_10_20_0),
		.out_wire_0_1(horizontal_tile_10_19_to_tile_10_20_1),
		.out_wire_0_2(horizontal_tile_10_19_to_tile_10_20_2),
		.out_wire_0_3(horizontal_tile_10_19_to_tile_10_20_3),
		.in_wire_0_0(horizontal_tile_10_20_to_tile_10_19_0),
		.in_wire_0_1(horizontal_tile_10_20_to_tile_10_19_1),
		.in_wire_0_2(horizontal_tile_10_20_to_tile_10_19_2),
		.in_wire_0_3(horizontal_tile_10_20_to_tile_10_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(340)
	);

	pe_tile pe_tile_10_20(
		.out_wire_3_0(vertical_tile_10_20_to_tile_9_20_0),
		.out_wire_3_1(vertical_tile_10_20_to_tile_9_20_1),
		.out_wire_3_2(vertical_tile_10_20_to_tile_9_20_2),
		.out_wire_3_3(vertical_tile_10_20_to_tile_9_20_3),
		.in_wire_3_0(vertical_tile_9_20_to_tile_10_20_0),
		.in_wire_3_1(vertical_tile_9_20_to_tile_10_20_1),
		.in_wire_3_2(vertical_tile_9_20_to_tile_10_20_2),
		.in_wire_3_3(vertical_tile_9_20_to_tile_10_20_3),
		.out_wire_1_0(vertical_tile_10_20_to_tile_11_20_0),
		.out_wire_1_1(vertical_tile_10_20_to_tile_11_20_1),
		.out_wire_1_2(vertical_tile_10_20_to_tile_11_20_2),
		.out_wire_1_3(vertical_tile_10_20_to_tile_11_20_3),
		.in_wire_1_0(vertical_tile_11_20_to_tile_10_20_0),
		.in_wire_1_1(vertical_tile_11_20_to_tile_10_20_1),
		.in_wire_1_2(vertical_tile_11_20_to_tile_10_20_2),
		.in_wire_1_3(vertical_tile_11_20_to_tile_10_20_3),
		.out_wire_2_0(horizontal_tile_10_20_to_tile_10_19_0),
		.out_wire_2_1(horizontal_tile_10_20_to_tile_10_19_1),
		.out_wire_2_2(horizontal_tile_10_20_to_tile_10_19_2),
		.out_wire_2_3(horizontal_tile_10_20_to_tile_10_19_3),
		.in_wire_2_0(horizontal_tile_10_19_to_tile_10_20_0),
		.in_wire_2_1(horizontal_tile_10_19_to_tile_10_20_1),
		.in_wire_2_2(horizontal_tile_10_19_to_tile_10_20_2),
		.in_wire_2_3(horizontal_tile_10_19_to_tile_10_20_3),
		.out_wire_0_0(horizontal_tile_10_20_to_tile_10_21_0),
		.out_wire_0_1(horizontal_tile_10_20_to_tile_10_21_1),
		.out_wire_0_2(horizontal_tile_10_20_to_tile_10_21_2),
		.out_wire_0_3(horizontal_tile_10_20_to_tile_10_21_3),
		.in_wire_0_0(horizontal_tile_10_21_to_tile_10_20_0),
		.in_wire_0_1(horizontal_tile_10_21_to_tile_10_20_1),
		.in_wire_0_2(horizontal_tile_10_21_to_tile_10_20_2),
		.in_wire_0_3(horizontal_tile_10_21_to_tile_10_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(341)
	);

	pe_tile pe_tile_10_21(
		.out_wire_3_0(vertical_tile_10_21_to_tile_9_21_0),
		.out_wire_3_1(vertical_tile_10_21_to_tile_9_21_1),
		.out_wire_3_2(vertical_tile_10_21_to_tile_9_21_2),
		.out_wire_3_3(vertical_tile_10_21_to_tile_9_21_3),
		.in_wire_3_0(vertical_tile_9_21_to_tile_10_21_0),
		.in_wire_3_1(vertical_tile_9_21_to_tile_10_21_1),
		.in_wire_3_2(vertical_tile_9_21_to_tile_10_21_2),
		.in_wire_3_3(vertical_tile_9_21_to_tile_10_21_3),
		.out_wire_1_0(vertical_tile_10_21_to_tile_11_21_0),
		.out_wire_1_1(vertical_tile_10_21_to_tile_11_21_1),
		.out_wire_1_2(vertical_tile_10_21_to_tile_11_21_2),
		.out_wire_1_3(vertical_tile_10_21_to_tile_11_21_3),
		.in_wire_1_0(vertical_tile_11_21_to_tile_10_21_0),
		.in_wire_1_1(vertical_tile_11_21_to_tile_10_21_1),
		.in_wire_1_2(vertical_tile_11_21_to_tile_10_21_2),
		.in_wire_1_3(vertical_tile_11_21_to_tile_10_21_3),
		.out_wire_2_0(horizontal_tile_10_21_to_tile_10_20_0),
		.out_wire_2_1(horizontal_tile_10_21_to_tile_10_20_1),
		.out_wire_2_2(horizontal_tile_10_21_to_tile_10_20_2),
		.out_wire_2_3(horizontal_tile_10_21_to_tile_10_20_3),
		.in_wire_2_0(horizontal_tile_10_20_to_tile_10_21_0),
		.in_wire_2_1(horizontal_tile_10_20_to_tile_10_21_1),
		.in_wire_2_2(horizontal_tile_10_20_to_tile_10_21_2),
		.in_wire_2_3(horizontal_tile_10_20_to_tile_10_21_3),
		.out_wire_0_0(horizontal_tile_10_21_to_tile_10_22_0),
		.out_wire_0_1(horizontal_tile_10_21_to_tile_10_22_1),
		.out_wire_0_2(horizontal_tile_10_21_to_tile_10_22_2),
		.out_wire_0_3(horizontal_tile_10_21_to_tile_10_22_3),
		.in_wire_0_0(horizontal_tile_10_22_to_tile_10_21_0),
		.in_wire_0_1(horizontal_tile_10_22_to_tile_10_21_1),
		.in_wire_0_2(horizontal_tile_10_22_to_tile_10_21_2),
		.in_wire_0_3(horizontal_tile_10_22_to_tile_10_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(342)
	);

	pe_tile pe_tile_10_22(
		.out_wire_3_0(vertical_tile_10_22_to_tile_9_22_0),
		.out_wire_3_1(vertical_tile_10_22_to_tile_9_22_1),
		.out_wire_3_2(vertical_tile_10_22_to_tile_9_22_2),
		.out_wire_3_3(vertical_tile_10_22_to_tile_9_22_3),
		.in_wire_3_0(vertical_tile_9_22_to_tile_10_22_0),
		.in_wire_3_1(vertical_tile_9_22_to_tile_10_22_1),
		.in_wire_3_2(vertical_tile_9_22_to_tile_10_22_2),
		.in_wire_3_3(vertical_tile_9_22_to_tile_10_22_3),
		.out_wire_1_0(vertical_tile_10_22_to_tile_11_22_0),
		.out_wire_1_1(vertical_tile_10_22_to_tile_11_22_1),
		.out_wire_1_2(vertical_tile_10_22_to_tile_11_22_2),
		.out_wire_1_3(vertical_tile_10_22_to_tile_11_22_3),
		.in_wire_1_0(vertical_tile_11_22_to_tile_10_22_0),
		.in_wire_1_1(vertical_tile_11_22_to_tile_10_22_1),
		.in_wire_1_2(vertical_tile_11_22_to_tile_10_22_2),
		.in_wire_1_3(vertical_tile_11_22_to_tile_10_22_3),
		.out_wire_2_0(horizontal_tile_10_22_to_tile_10_21_0),
		.out_wire_2_1(horizontal_tile_10_22_to_tile_10_21_1),
		.out_wire_2_2(horizontal_tile_10_22_to_tile_10_21_2),
		.out_wire_2_3(horizontal_tile_10_22_to_tile_10_21_3),
		.in_wire_2_0(horizontal_tile_10_21_to_tile_10_22_0),
		.in_wire_2_1(horizontal_tile_10_21_to_tile_10_22_1),
		.in_wire_2_2(horizontal_tile_10_21_to_tile_10_22_2),
		.in_wire_2_3(horizontal_tile_10_21_to_tile_10_22_3),
		.out_wire_0_0(horizontal_tile_10_22_to_tile_10_23_0),
		.out_wire_0_1(horizontal_tile_10_22_to_tile_10_23_1),
		.out_wire_0_2(horizontal_tile_10_22_to_tile_10_23_2),
		.out_wire_0_3(horizontal_tile_10_22_to_tile_10_23_3),
		.in_wire_0_0(horizontal_tile_10_23_to_tile_10_22_0),
		.in_wire_0_1(horizontal_tile_10_23_to_tile_10_22_1),
		.in_wire_0_2(horizontal_tile_10_23_to_tile_10_22_2),
		.in_wire_0_3(horizontal_tile_10_23_to_tile_10_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(343)
	);

	pe_tile pe_tile_10_23(
		.out_wire_3_0(vertical_tile_10_23_to_tile_9_23_0),
		.out_wire_3_1(vertical_tile_10_23_to_tile_9_23_1),
		.out_wire_3_2(vertical_tile_10_23_to_tile_9_23_2),
		.out_wire_3_3(vertical_tile_10_23_to_tile_9_23_3),
		.in_wire_3_0(vertical_tile_9_23_to_tile_10_23_0),
		.in_wire_3_1(vertical_tile_9_23_to_tile_10_23_1),
		.in_wire_3_2(vertical_tile_9_23_to_tile_10_23_2),
		.in_wire_3_3(vertical_tile_9_23_to_tile_10_23_3),
		.out_wire_1_0(vertical_tile_10_23_to_tile_11_23_0),
		.out_wire_1_1(vertical_tile_10_23_to_tile_11_23_1),
		.out_wire_1_2(vertical_tile_10_23_to_tile_11_23_2),
		.out_wire_1_3(vertical_tile_10_23_to_tile_11_23_3),
		.in_wire_1_0(vertical_tile_11_23_to_tile_10_23_0),
		.in_wire_1_1(vertical_tile_11_23_to_tile_10_23_1),
		.in_wire_1_2(vertical_tile_11_23_to_tile_10_23_2),
		.in_wire_1_3(vertical_tile_11_23_to_tile_10_23_3),
		.out_wire_2_0(horizontal_tile_10_23_to_tile_10_22_0),
		.out_wire_2_1(horizontal_tile_10_23_to_tile_10_22_1),
		.out_wire_2_2(horizontal_tile_10_23_to_tile_10_22_2),
		.out_wire_2_3(horizontal_tile_10_23_to_tile_10_22_3),
		.in_wire_2_0(horizontal_tile_10_22_to_tile_10_23_0),
		.in_wire_2_1(horizontal_tile_10_22_to_tile_10_23_1),
		.in_wire_2_2(horizontal_tile_10_22_to_tile_10_23_2),
		.in_wire_2_3(horizontal_tile_10_22_to_tile_10_23_3),
		.out_wire_0_0(horizontal_tile_10_23_to_tile_10_24_0),
		.out_wire_0_1(horizontal_tile_10_23_to_tile_10_24_1),
		.out_wire_0_2(horizontal_tile_10_23_to_tile_10_24_2),
		.out_wire_0_3(horizontal_tile_10_23_to_tile_10_24_3),
		.in_wire_0_0(horizontal_tile_10_24_to_tile_10_23_0),
		.in_wire_0_1(horizontal_tile_10_24_to_tile_10_23_1),
		.in_wire_0_2(horizontal_tile_10_24_to_tile_10_23_2),
		.in_wire_0_3(horizontal_tile_10_24_to_tile_10_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(344)
	);

	pe_tile pe_tile_10_24(
		.out_wire_3_0(vertical_tile_10_24_to_tile_9_24_0),
		.out_wire_3_1(vertical_tile_10_24_to_tile_9_24_1),
		.out_wire_3_2(vertical_tile_10_24_to_tile_9_24_2),
		.out_wire_3_3(vertical_tile_10_24_to_tile_9_24_3),
		.in_wire_3_0(vertical_tile_9_24_to_tile_10_24_0),
		.in_wire_3_1(vertical_tile_9_24_to_tile_10_24_1),
		.in_wire_3_2(vertical_tile_9_24_to_tile_10_24_2),
		.in_wire_3_3(vertical_tile_9_24_to_tile_10_24_3),
		.out_wire_1_0(vertical_tile_10_24_to_tile_11_24_0),
		.out_wire_1_1(vertical_tile_10_24_to_tile_11_24_1),
		.out_wire_1_2(vertical_tile_10_24_to_tile_11_24_2),
		.out_wire_1_3(vertical_tile_10_24_to_tile_11_24_3),
		.in_wire_1_0(vertical_tile_11_24_to_tile_10_24_0),
		.in_wire_1_1(vertical_tile_11_24_to_tile_10_24_1),
		.in_wire_1_2(vertical_tile_11_24_to_tile_10_24_2),
		.in_wire_1_3(vertical_tile_11_24_to_tile_10_24_3),
		.out_wire_2_0(horizontal_tile_10_24_to_tile_10_23_0),
		.out_wire_2_1(horizontal_tile_10_24_to_tile_10_23_1),
		.out_wire_2_2(horizontal_tile_10_24_to_tile_10_23_2),
		.out_wire_2_3(horizontal_tile_10_24_to_tile_10_23_3),
		.in_wire_2_0(horizontal_tile_10_23_to_tile_10_24_0),
		.in_wire_2_1(horizontal_tile_10_23_to_tile_10_24_1),
		.in_wire_2_2(horizontal_tile_10_23_to_tile_10_24_2),
		.in_wire_2_3(horizontal_tile_10_23_to_tile_10_24_3),
		.out_wire_0_0(horizontal_tile_10_24_to_tile_10_25_0),
		.out_wire_0_1(horizontal_tile_10_24_to_tile_10_25_1),
		.out_wire_0_2(horizontal_tile_10_24_to_tile_10_25_2),
		.out_wire_0_3(horizontal_tile_10_24_to_tile_10_25_3),
		.in_wire_0_0(horizontal_tile_10_25_to_tile_10_24_0),
		.in_wire_0_1(horizontal_tile_10_25_to_tile_10_24_1),
		.in_wire_0_2(horizontal_tile_10_25_to_tile_10_24_2),
		.in_wire_0_3(horizontal_tile_10_25_to_tile_10_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(345)
	);

	pe_tile pe_tile_10_25(
		.out_wire_3_0(vertical_tile_10_25_to_tile_9_25_0),
		.out_wire_3_1(vertical_tile_10_25_to_tile_9_25_1),
		.out_wire_3_2(vertical_tile_10_25_to_tile_9_25_2),
		.out_wire_3_3(vertical_tile_10_25_to_tile_9_25_3),
		.in_wire_3_0(vertical_tile_9_25_to_tile_10_25_0),
		.in_wire_3_1(vertical_tile_9_25_to_tile_10_25_1),
		.in_wire_3_2(vertical_tile_9_25_to_tile_10_25_2),
		.in_wire_3_3(vertical_tile_9_25_to_tile_10_25_3),
		.out_wire_1_0(vertical_tile_10_25_to_tile_11_25_0),
		.out_wire_1_1(vertical_tile_10_25_to_tile_11_25_1),
		.out_wire_1_2(vertical_tile_10_25_to_tile_11_25_2),
		.out_wire_1_3(vertical_tile_10_25_to_tile_11_25_3),
		.in_wire_1_0(vertical_tile_11_25_to_tile_10_25_0),
		.in_wire_1_1(vertical_tile_11_25_to_tile_10_25_1),
		.in_wire_1_2(vertical_tile_11_25_to_tile_10_25_2),
		.in_wire_1_3(vertical_tile_11_25_to_tile_10_25_3),
		.out_wire_2_0(horizontal_tile_10_25_to_tile_10_24_0),
		.out_wire_2_1(horizontal_tile_10_25_to_tile_10_24_1),
		.out_wire_2_2(horizontal_tile_10_25_to_tile_10_24_2),
		.out_wire_2_3(horizontal_tile_10_25_to_tile_10_24_3),
		.in_wire_2_0(horizontal_tile_10_24_to_tile_10_25_0),
		.in_wire_2_1(horizontal_tile_10_24_to_tile_10_25_1),
		.in_wire_2_2(horizontal_tile_10_24_to_tile_10_25_2),
		.in_wire_2_3(horizontal_tile_10_24_to_tile_10_25_3),
		.out_wire_0_0(horizontal_tile_10_25_to_tile_10_26_0),
		.out_wire_0_1(horizontal_tile_10_25_to_tile_10_26_1),
		.out_wire_0_2(horizontal_tile_10_25_to_tile_10_26_2),
		.out_wire_0_3(horizontal_tile_10_25_to_tile_10_26_3),
		.in_wire_0_0(horizontal_tile_10_26_to_tile_10_25_0),
		.in_wire_0_1(horizontal_tile_10_26_to_tile_10_25_1),
		.in_wire_0_2(horizontal_tile_10_26_to_tile_10_25_2),
		.in_wire_0_3(horizontal_tile_10_26_to_tile_10_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(346)
	);

	pe_tile pe_tile_10_26(
		.out_wire_3_0(vertical_tile_10_26_to_tile_9_26_0),
		.out_wire_3_1(vertical_tile_10_26_to_tile_9_26_1),
		.out_wire_3_2(vertical_tile_10_26_to_tile_9_26_2),
		.out_wire_3_3(vertical_tile_10_26_to_tile_9_26_3),
		.in_wire_3_0(vertical_tile_9_26_to_tile_10_26_0),
		.in_wire_3_1(vertical_tile_9_26_to_tile_10_26_1),
		.in_wire_3_2(vertical_tile_9_26_to_tile_10_26_2),
		.in_wire_3_3(vertical_tile_9_26_to_tile_10_26_3),
		.out_wire_1_0(vertical_tile_10_26_to_tile_11_26_0),
		.out_wire_1_1(vertical_tile_10_26_to_tile_11_26_1),
		.out_wire_1_2(vertical_tile_10_26_to_tile_11_26_2),
		.out_wire_1_3(vertical_tile_10_26_to_tile_11_26_3),
		.in_wire_1_0(vertical_tile_11_26_to_tile_10_26_0),
		.in_wire_1_1(vertical_tile_11_26_to_tile_10_26_1),
		.in_wire_1_2(vertical_tile_11_26_to_tile_10_26_2),
		.in_wire_1_3(vertical_tile_11_26_to_tile_10_26_3),
		.out_wire_2_0(horizontal_tile_10_26_to_tile_10_25_0),
		.out_wire_2_1(horizontal_tile_10_26_to_tile_10_25_1),
		.out_wire_2_2(horizontal_tile_10_26_to_tile_10_25_2),
		.out_wire_2_3(horizontal_tile_10_26_to_tile_10_25_3),
		.in_wire_2_0(horizontal_tile_10_25_to_tile_10_26_0),
		.in_wire_2_1(horizontal_tile_10_25_to_tile_10_26_1),
		.in_wire_2_2(horizontal_tile_10_25_to_tile_10_26_2),
		.in_wire_2_3(horizontal_tile_10_25_to_tile_10_26_3),
		.out_wire_0_0(horizontal_tile_10_26_to_tile_10_27_0),
		.out_wire_0_1(horizontal_tile_10_26_to_tile_10_27_1),
		.out_wire_0_2(horizontal_tile_10_26_to_tile_10_27_2),
		.out_wire_0_3(horizontal_tile_10_26_to_tile_10_27_3),
		.in_wire_0_0(horizontal_tile_10_27_to_tile_10_26_0),
		.in_wire_0_1(horizontal_tile_10_27_to_tile_10_26_1),
		.in_wire_0_2(horizontal_tile_10_27_to_tile_10_26_2),
		.in_wire_0_3(horizontal_tile_10_27_to_tile_10_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(347)
	);

	pe_tile pe_tile_10_27(
		.out_wire_3_0(vertical_tile_10_27_to_tile_9_27_0),
		.out_wire_3_1(vertical_tile_10_27_to_tile_9_27_1),
		.out_wire_3_2(vertical_tile_10_27_to_tile_9_27_2),
		.out_wire_3_3(vertical_tile_10_27_to_tile_9_27_3),
		.in_wire_3_0(vertical_tile_9_27_to_tile_10_27_0),
		.in_wire_3_1(vertical_tile_9_27_to_tile_10_27_1),
		.in_wire_3_2(vertical_tile_9_27_to_tile_10_27_2),
		.in_wire_3_3(vertical_tile_9_27_to_tile_10_27_3),
		.out_wire_1_0(vertical_tile_10_27_to_tile_11_27_0),
		.out_wire_1_1(vertical_tile_10_27_to_tile_11_27_1),
		.out_wire_1_2(vertical_tile_10_27_to_tile_11_27_2),
		.out_wire_1_3(vertical_tile_10_27_to_tile_11_27_3),
		.in_wire_1_0(vertical_tile_11_27_to_tile_10_27_0),
		.in_wire_1_1(vertical_tile_11_27_to_tile_10_27_1),
		.in_wire_1_2(vertical_tile_11_27_to_tile_10_27_2),
		.in_wire_1_3(vertical_tile_11_27_to_tile_10_27_3),
		.out_wire_2_0(horizontal_tile_10_27_to_tile_10_26_0),
		.out_wire_2_1(horizontal_tile_10_27_to_tile_10_26_1),
		.out_wire_2_2(horizontal_tile_10_27_to_tile_10_26_2),
		.out_wire_2_3(horizontal_tile_10_27_to_tile_10_26_3),
		.in_wire_2_0(horizontal_tile_10_26_to_tile_10_27_0),
		.in_wire_2_1(horizontal_tile_10_26_to_tile_10_27_1),
		.in_wire_2_2(horizontal_tile_10_26_to_tile_10_27_2),
		.in_wire_2_3(horizontal_tile_10_26_to_tile_10_27_3),
		.out_wire_0_0(horizontal_tile_10_27_to_tile_10_28_0),
		.out_wire_0_1(horizontal_tile_10_27_to_tile_10_28_1),
		.out_wire_0_2(horizontal_tile_10_27_to_tile_10_28_2),
		.out_wire_0_3(horizontal_tile_10_27_to_tile_10_28_3),
		.in_wire_0_0(horizontal_tile_10_28_to_tile_10_27_0),
		.in_wire_0_1(horizontal_tile_10_28_to_tile_10_27_1),
		.in_wire_0_2(horizontal_tile_10_28_to_tile_10_27_2),
		.in_wire_0_3(horizontal_tile_10_28_to_tile_10_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(348)
	);

	pe_tile pe_tile_10_28(
		.out_wire_3_0(vertical_tile_10_28_to_tile_9_28_0),
		.out_wire_3_1(vertical_tile_10_28_to_tile_9_28_1),
		.out_wire_3_2(vertical_tile_10_28_to_tile_9_28_2),
		.out_wire_3_3(vertical_tile_10_28_to_tile_9_28_3),
		.in_wire_3_0(vertical_tile_9_28_to_tile_10_28_0),
		.in_wire_3_1(vertical_tile_9_28_to_tile_10_28_1),
		.in_wire_3_2(vertical_tile_9_28_to_tile_10_28_2),
		.in_wire_3_3(vertical_tile_9_28_to_tile_10_28_3),
		.out_wire_1_0(vertical_tile_10_28_to_tile_11_28_0),
		.out_wire_1_1(vertical_tile_10_28_to_tile_11_28_1),
		.out_wire_1_2(vertical_tile_10_28_to_tile_11_28_2),
		.out_wire_1_3(vertical_tile_10_28_to_tile_11_28_3),
		.in_wire_1_0(vertical_tile_11_28_to_tile_10_28_0),
		.in_wire_1_1(vertical_tile_11_28_to_tile_10_28_1),
		.in_wire_1_2(vertical_tile_11_28_to_tile_10_28_2),
		.in_wire_1_3(vertical_tile_11_28_to_tile_10_28_3),
		.out_wire_2_0(horizontal_tile_10_28_to_tile_10_27_0),
		.out_wire_2_1(horizontal_tile_10_28_to_tile_10_27_1),
		.out_wire_2_2(horizontal_tile_10_28_to_tile_10_27_2),
		.out_wire_2_3(horizontal_tile_10_28_to_tile_10_27_3),
		.in_wire_2_0(horizontal_tile_10_27_to_tile_10_28_0),
		.in_wire_2_1(horizontal_tile_10_27_to_tile_10_28_1),
		.in_wire_2_2(horizontal_tile_10_27_to_tile_10_28_2),
		.in_wire_2_3(horizontal_tile_10_27_to_tile_10_28_3),
		.out_wire_0_0(horizontal_tile_10_28_to_tile_10_29_0),
		.out_wire_0_1(horizontal_tile_10_28_to_tile_10_29_1),
		.out_wire_0_2(horizontal_tile_10_28_to_tile_10_29_2),
		.out_wire_0_3(horizontal_tile_10_28_to_tile_10_29_3),
		.in_wire_0_0(horizontal_tile_10_29_to_tile_10_28_0),
		.in_wire_0_1(horizontal_tile_10_29_to_tile_10_28_1),
		.in_wire_0_2(horizontal_tile_10_29_to_tile_10_28_2),
		.in_wire_0_3(horizontal_tile_10_29_to_tile_10_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(349)
	);

	pe_tile pe_tile_10_29(
		.out_wire_3_0(vertical_tile_10_29_to_tile_9_29_0),
		.out_wire_3_1(vertical_tile_10_29_to_tile_9_29_1),
		.out_wire_3_2(vertical_tile_10_29_to_tile_9_29_2),
		.out_wire_3_3(vertical_tile_10_29_to_tile_9_29_3),
		.in_wire_3_0(vertical_tile_9_29_to_tile_10_29_0),
		.in_wire_3_1(vertical_tile_9_29_to_tile_10_29_1),
		.in_wire_3_2(vertical_tile_9_29_to_tile_10_29_2),
		.in_wire_3_3(vertical_tile_9_29_to_tile_10_29_3),
		.out_wire_1_0(vertical_tile_10_29_to_tile_11_29_0),
		.out_wire_1_1(vertical_tile_10_29_to_tile_11_29_1),
		.out_wire_1_2(vertical_tile_10_29_to_tile_11_29_2),
		.out_wire_1_3(vertical_tile_10_29_to_tile_11_29_3),
		.in_wire_1_0(vertical_tile_11_29_to_tile_10_29_0),
		.in_wire_1_1(vertical_tile_11_29_to_tile_10_29_1),
		.in_wire_1_2(vertical_tile_11_29_to_tile_10_29_2),
		.in_wire_1_3(vertical_tile_11_29_to_tile_10_29_3),
		.out_wire_2_0(horizontal_tile_10_29_to_tile_10_28_0),
		.out_wire_2_1(horizontal_tile_10_29_to_tile_10_28_1),
		.out_wire_2_2(horizontal_tile_10_29_to_tile_10_28_2),
		.out_wire_2_3(horizontal_tile_10_29_to_tile_10_28_3),
		.in_wire_2_0(horizontal_tile_10_28_to_tile_10_29_0),
		.in_wire_2_1(horizontal_tile_10_28_to_tile_10_29_1),
		.in_wire_2_2(horizontal_tile_10_28_to_tile_10_29_2),
		.in_wire_2_3(horizontal_tile_10_28_to_tile_10_29_3),
		.out_wire_0_0(horizontal_tile_10_29_to_tile_10_30_0),
		.out_wire_0_1(horizontal_tile_10_29_to_tile_10_30_1),
		.out_wire_0_2(horizontal_tile_10_29_to_tile_10_30_2),
		.out_wire_0_3(horizontal_tile_10_29_to_tile_10_30_3),
		.in_wire_0_0(horizontal_tile_10_30_to_tile_10_29_0),
		.in_wire_0_1(horizontal_tile_10_30_to_tile_10_29_1),
		.in_wire_0_2(horizontal_tile_10_30_to_tile_10_29_2),
		.in_wire_0_3(horizontal_tile_10_30_to_tile_10_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(350)
	);

	pe_tile pe_tile_10_30(
		.out_wire_3_0(vertical_tile_10_30_to_tile_9_30_0),
		.out_wire_3_1(vertical_tile_10_30_to_tile_9_30_1),
		.out_wire_3_2(vertical_tile_10_30_to_tile_9_30_2),
		.out_wire_3_3(vertical_tile_10_30_to_tile_9_30_3),
		.in_wire_3_0(vertical_tile_9_30_to_tile_10_30_0),
		.in_wire_3_1(vertical_tile_9_30_to_tile_10_30_1),
		.in_wire_3_2(vertical_tile_9_30_to_tile_10_30_2),
		.in_wire_3_3(vertical_tile_9_30_to_tile_10_30_3),
		.out_wire_1_0(vertical_tile_10_30_to_tile_11_30_0),
		.out_wire_1_1(vertical_tile_10_30_to_tile_11_30_1),
		.out_wire_1_2(vertical_tile_10_30_to_tile_11_30_2),
		.out_wire_1_3(vertical_tile_10_30_to_tile_11_30_3),
		.in_wire_1_0(vertical_tile_11_30_to_tile_10_30_0),
		.in_wire_1_1(vertical_tile_11_30_to_tile_10_30_1),
		.in_wire_1_2(vertical_tile_11_30_to_tile_10_30_2),
		.in_wire_1_3(vertical_tile_11_30_to_tile_10_30_3),
		.out_wire_2_0(horizontal_tile_10_30_to_tile_10_29_0),
		.out_wire_2_1(horizontal_tile_10_30_to_tile_10_29_1),
		.out_wire_2_2(horizontal_tile_10_30_to_tile_10_29_2),
		.out_wire_2_3(horizontal_tile_10_30_to_tile_10_29_3),
		.in_wire_2_0(horizontal_tile_10_29_to_tile_10_30_0),
		.in_wire_2_1(horizontal_tile_10_29_to_tile_10_30_1),
		.in_wire_2_2(horizontal_tile_10_29_to_tile_10_30_2),
		.in_wire_2_3(horizontal_tile_10_29_to_tile_10_30_3),
		.out_wire_0_0(horizontal_tile_10_30_to_tile_10_31_0),
		.out_wire_0_1(horizontal_tile_10_30_to_tile_10_31_1),
		.out_wire_0_2(horizontal_tile_10_30_to_tile_10_31_2),
		.out_wire_0_3(horizontal_tile_10_30_to_tile_10_31_3),
		.in_wire_0_0(horizontal_tile_10_31_to_tile_10_30_0),
		.in_wire_0_1(horizontal_tile_10_31_to_tile_10_30_1),
		.in_wire_0_2(horizontal_tile_10_31_to_tile_10_30_2),
		.in_wire_0_3(horizontal_tile_10_31_to_tile_10_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(351)
	);

	pe_tile_right pe_tile_10_31(
		.out_wire_3_0(vertical_tile_10_31_to_tile_9_31_0),
		.out_wire_3_1(vertical_tile_10_31_to_tile_9_31_1),
		.out_wire_3_2(vertical_tile_10_31_to_tile_9_31_2),
		.out_wire_3_3(vertical_tile_10_31_to_tile_9_31_3),
		.in_wire_3_0(vertical_tile_9_31_to_tile_10_31_0),
		.in_wire_3_1(vertical_tile_9_31_to_tile_10_31_1),
		.in_wire_3_2(vertical_tile_9_31_to_tile_10_31_2),
		.in_wire_3_3(vertical_tile_9_31_to_tile_10_31_3),
		.out_wire_1_0(vertical_tile_10_31_to_tile_11_31_0),
		.out_wire_1_1(vertical_tile_10_31_to_tile_11_31_1),
		.out_wire_1_2(vertical_tile_10_31_to_tile_11_31_2),
		.out_wire_1_3(vertical_tile_10_31_to_tile_11_31_3),
		.in_wire_1_0(vertical_tile_11_31_to_tile_10_31_0),
		.in_wire_1_1(vertical_tile_11_31_to_tile_10_31_1),
		.in_wire_1_2(vertical_tile_11_31_to_tile_10_31_2),
		.in_wire_1_3(vertical_tile_11_31_to_tile_10_31_3),
		.out_wire_2_0(horizontal_tile_10_31_to_tile_10_30_0),
		.out_wire_2_1(horizontal_tile_10_31_to_tile_10_30_1),
		.out_wire_2_2(horizontal_tile_10_31_to_tile_10_30_2),
		.out_wire_2_3(horizontal_tile_10_31_to_tile_10_30_3),
		.in_wire_2_0(horizontal_tile_10_30_to_tile_10_31_0),
		.in_wire_2_1(horizontal_tile_10_30_to_tile_10_31_1),
		.in_wire_2_2(horizontal_tile_10_30_to_tile_10_31_2),
		.in_wire_2_3(horizontal_tile_10_30_to_tile_10_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(352)
	);

	pe_tile_left pe_tile_11_0(
		.out_wire_3_0(vertical_tile_11_0_to_tile_10_0_0),
		.out_wire_3_1(vertical_tile_11_0_to_tile_10_0_1),
		.out_wire_3_2(vertical_tile_11_0_to_tile_10_0_2),
		.out_wire_3_3(vertical_tile_11_0_to_tile_10_0_3),
		.in_wire_3_0(vertical_tile_10_0_to_tile_11_0_0),
		.in_wire_3_1(vertical_tile_10_0_to_tile_11_0_1),
		.in_wire_3_2(vertical_tile_10_0_to_tile_11_0_2),
		.in_wire_3_3(vertical_tile_10_0_to_tile_11_0_3),
		.out_wire_1_0(vertical_tile_11_0_to_tile_12_0_0),
		.out_wire_1_1(vertical_tile_11_0_to_tile_12_0_1),
		.out_wire_1_2(vertical_tile_11_0_to_tile_12_0_2),
		.out_wire_1_3(vertical_tile_11_0_to_tile_12_0_3),
		.in_wire_1_0(vertical_tile_12_0_to_tile_11_0_0),
		.in_wire_1_1(vertical_tile_12_0_to_tile_11_0_1),
		.in_wire_1_2(vertical_tile_12_0_to_tile_11_0_2),
		.in_wire_1_3(vertical_tile_12_0_to_tile_11_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_11_0_to_tile_11_1_0),
		.out_wire_0_1(horizontal_tile_11_0_to_tile_11_1_1),
		.out_wire_0_2(horizontal_tile_11_0_to_tile_11_1_2),
		.out_wire_0_3(horizontal_tile_11_0_to_tile_11_1_3),
		.in_wire_0_0(horizontal_tile_11_1_to_tile_11_0_0),
		.in_wire_0_1(horizontal_tile_11_1_to_tile_11_0_1),
		.in_wire_0_2(horizontal_tile_11_1_to_tile_11_0_2),
		.in_wire_0_3(horizontal_tile_11_1_to_tile_11_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(353)
	);

	pe_tile pe_tile_11_1(
		.out_wire_3_0(vertical_tile_11_1_to_tile_10_1_0),
		.out_wire_3_1(vertical_tile_11_1_to_tile_10_1_1),
		.out_wire_3_2(vertical_tile_11_1_to_tile_10_1_2),
		.out_wire_3_3(vertical_tile_11_1_to_tile_10_1_3),
		.in_wire_3_0(vertical_tile_10_1_to_tile_11_1_0),
		.in_wire_3_1(vertical_tile_10_1_to_tile_11_1_1),
		.in_wire_3_2(vertical_tile_10_1_to_tile_11_1_2),
		.in_wire_3_3(vertical_tile_10_1_to_tile_11_1_3),
		.out_wire_1_0(vertical_tile_11_1_to_tile_12_1_0),
		.out_wire_1_1(vertical_tile_11_1_to_tile_12_1_1),
		.out_wire_1_2(vertical_tile_11_1_to_tile_12_1_2),
		.out_wire_1_3(vertical_tile_11_1_to_tile_12_1_3),
		.in_wire_1_0(vertical_tile_12_1_to_tile_11_1_0),
		.in_wire_1_1(vertical_tile_12_1_to_tile_11_1_1),
		.in_wire_1_2(vertical_tile_12_1_to_tile_11_1_2),
		.in_wire_1_3(vertical_tile_12_1_to_tile_11_1_3),
		.out_wire_2_0(horizontal_tile_11_1_to_tile_11_0_0),
		.out_wire_2_1(horizontal_tile_11_1_to_tile_11_0_1),
		.out_wire_2_2(horizontal_tile_11_1_to_tile_11_0_2),
		.out_wire_2_3(horizontal_tile_11_1_to_tile_11_0_3),
		.in_wire_2_0(horizontal_tile_11_0_to_tile_11_1_0),
		.in_wire_2_1(horizontal_tile_11_0_to_tile_11_1_1),
		.in_wire_2_2(horizontal_tile_11_0_to_tile_11_1_2),
		.in_wire_2_3(horizontal_tile_11_0_to_tile_11_1_3),
		.out_wire_0_0(horizontal_tile_11_1_to_tile_11_2_0),
		.out_wire_0_1(horizontal_tile_11_1_to_tile_11_2_1),
		.out_wire_0_2(horizontal_tile_11_1_to_tile_11_2_2),
		.out_wire_0_3(horizontal_tile_11_1_to_tile_11_2_3),
		.in_wire_0_0(horizontal_tile_11_2_to_tile_11_1_0),
		.in_wire_0_1(horizontal_tile_11_2_to_tile_11_1_1),
		.in_wire_0_2(horizontal_tile_11_2_to_tile_11_1_2),
		.in_wire_0_3(horizontal_tile_11_2_to_tile_11_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(354)
	);

	pe_tile pe_tile_11_2(
		.out_wire_3_0(vertical_tile_11_2_to_tile_10_2_0),
		.out_wire_3_1(vertical_tile_11_2_to_tile_10_2_1),
		.out_wire_3_2(vertical_tile_11_2_to_tile_10_2_2),
		.out_wire_3_3(vertical_tile_11_2_to_tile_10_2_3),
		.in_wire_3_0(vertical_tile_10_2_to_tile_11_2_0),
		.in_wire_3_1(vertical_tile_10_2_to_tile_11_2_1),
		.in_wire_3_2(vertical_tile_10_2_to_tile_11_2_2),
		.in_wire_3_3(vertical_tile_10_2_to_tile_11_2_3),
		.out_wire_1_0(vertical_tile_11_2_to_tile_12_2_0),
		.out_wire_1_1(vertical_tile_11_2_to_tile_12_2_1),
		.out_wire_1_2(vertical_tile_11_2_to_tile_12_2_2),
		.out_wire_1_3(vertical_tile_11_2_to_tile_12_2_3),
		.in_wire_1_0(vertical_tile_12_2_to_tile_11_2_0),
		.in_wire_1_1(vertical_tile_12_2_to_tile_11_2_1),
		.in_wire_1_2(vertical_tile_12_2_to_tile_11_2_2),
		.in_wire_1_3(vertical_tile_12_2_to_tile_11_2_3),
		.out_wire_2_0(horizontal_tile_11_2_to_tile_11_1_0),
		.out_wire_2_1(horizontal_tile_11_2_to_tile_11_1_1),
		.out_wire_2_2(horizontal_tile_11_2_to_tile_11_1_2),
		.out_wire_2_3(horizontal_tile_11_2_to_tile_11_1_3),
		.in_wire_2_0(horizontal_tile_11_1_to_tile_11_2_0),
		.in_wire_2_1(horizontal_tile_11_1_to_tile_11_2_1),
		.in_wire_2_2(horizontal_tile_11_1_to_tile_11_2_2),
		.in_wire_2_3(horizontal_tile_11_1_to_tile_11_2_3),
		.out_wire_0_0(horizontal_tile_11_2_to_tile_11_3_0),
		.out_wire_0_1(horizontal_tile_11_2_to_tile_11_3_1),
		.out_wire_0_2(horizontal_tile_11_2_to_tile_11_3_2),
		.out_wire_0_3(horizontal_tile_11_2_to_tile_11_3_3),
		.in_wire_0_0(horizontal_tile_11_3_to_tile_11_2_0),
		.in_wire_0_1(horizontal_tile_11_3_to_tile_11_2_1),
		.in_wire_0_2(horizontal_tile_11_3_to_tile_11_2_2),
		.in_wire_0_3(horizontal_tile_11_3_to_tile_11_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(355)
	);

	pe_tile pe_tile_11_3(
		.out_wire_3_0(vertical_tile_11_3_to_tile_10_3_0),
		.out_wire_3_1(vertical_tile_11_3_to_tile_10_3_1),
		.out_wire_3_2(vertical_tile_11_3_to_tile_10_3_2),
		.out_wire_3_3(vertical_tile_11_3_to_tile_10_3_3),
		.in_wire_3_0(vertical_tile_10_3_to_tile_11_3_0),
		.in_wire_3_1(vertical_tile_10_3_to_tile_11_3_1),
		.in_wire_3_2(vertical_tile_10_3_to_tile_11_3_2),
		.in_wire_3_3(vertical_tile_10_3_to_tile_11_3_3),
		.out_wire_1_0(vertical_tile_11_3_to_tile_12_3_0),
		.out_wire_1_1(vertical_tile_11_3_to_tile_12_3_1),
		.out_wire_1_2(vertical_tile_11_3_to_tile_12_3_2),
		.out_wire_1_3(vertical_tile_11_3_to_tile_12_3_3),
		.in_wire_1_0(vertical_tile_12_3_to_tile_11_3_0),
		.in_wire_1_1(vertical_tile_12_3_to_tile_11_3_1),
		.in_wire_1_2(vertical_tile_12_3_to_tile_11_3_2),
		.in_wire_1_3(vertical_tile_12_3_to_tile_11_3_3),
		.out_wire_2_0(horizontal_tile_11_3_to_tile_11_2_0),
		.out_wire_2_1(horizontal_tile_11_3_to_tile_11_2_1),
		.out_wire_2_2(horizontal_tile_11_3_to_tile_11_2_2),
		.out_wire_2_3(horizontal_tile_11_3_to_tile_11_2_3),
		.in_wire_2_0(horizontal_tile_11_2_to_tile_11_3_0),
		.in_wire_2_1(horizontal_tile_11_2_to_tile_11_3_1),
		.in_wire_2_2(horizontal_tile_11_2_to_tile_11_3_2),
		.in_wire_2_3(horizontal_tile_11_2_to_tile_11_3_3),
		.out_wire_0_0(horizontal_tile_11_3_to_tile_11_4_0),
		.out_wire_0_1(horizontal_tile_11_3_to_tile_11_4_1),
		.out_wire_0_2(horizontal_tile_11_3_to_tile_11_4_2),
		.out_wire_0_3(horizontal_tile_11_3_to_tile_11_4_3),
		.in_wire_0_0(horizontal_tile_11_4_to_tile_11_3_0),
		.in_wire_0_1(horizontal_tile_11_4_to_tile_11_3_1),
		.in_wire_0_2(horizontal_tile_11_4_to_tile_11_3_2),
		.in_wire_0_3(horizontal_tile_11_4_to_tile_11_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(356)
	);

	pe_tile pe_tile_11_4(
		.out_wire_3_0(vertical_tile_11_4_to_tile_10_4_0),
		.out_wire_3_1(vertical_tile_11_4_to_tile_10_4_1),
		.out_wire_3_2(vertical_tile_11_4_to_tile_10_4_2),
		.out_wire_3_3(vertical_tile_11_4_to_tile_10_4_3),
		.in_wire_3_0(vertical_tile_10_4_to_tile_11_4_0),
		.in_wire_3_1(vertical_tile_10_4_to_tile_11_4_1),
		.in_wire_3_2(vertical_tile_10_4_to_tile_11_4_2),
		.in_wire_3_3(vertical_tile_10_4_to_tile_11_4_3),
		.out_wire_1_0(vertical_tile_11_4_to_tile_12_4_0),
		.out_wire_1_1(vertical_tile_11_4_to_tile_12_4_1),
		.out_wire_1_2(vertical_tile_11_4_to_tile_12_4_2),
		.out_wire_1_3(vertical_tile_11_4_to_tile_12_4_3),
		.in_wire_1_0(vertical_tile_12_4_to_tile_11_4_0),
		.in_wire_1_1(vertical_tile_12_4_to_tile_11_4_1),
		.in_wire_1_2(vertical_tile_12_4_to_tile_11_4_2),
		.in_wire_1_3(vertical_tile_12_4_to_tile_11_4_3),
		.out_wire_2_0(horizontal_tile_11_4_to_tile_11_3_0),
		.out_wire_2_1(horizontal_tile_11_4_to_tile_11_3_1),
		.out_wire_2_2(horizontal_tile_11_4_to_tile_11_3_2),
		.out_wire_2_3(horizontal_tile_11_4_to_tile_11_3_3),
		.in_wire_2_0(horizontal_tile_11_3_to_tile_11_4_0),
		.in_wire_2_1(horizontal_tile_11_3_to_tile_11_4_1),
		.in_wire_2_2(horizontal_tile_11_3_to_tile_11_4_2),
		.in_wire_2_3(horizontal_tile_11_3_to_tile_11_4_3),
		.out_wire_0_0(horizontal_tile_11_4_to_tile_11_5_0),
		.out_wire_0_1(horizontal_tile_11_4_to_tile_11_5_1),
		.out_wire_0_2(horizontal_tile_11_4_to_tile_11_5_2),
		.out_wire_0_3(horizontal_tile_11_4_to_tile_11_5_3),
		.in_wire_0_0(horizontal_tile_11_5_to_tile_11_4_0),
		.in_wire_0_1(horizontal_tile_11_5_to_tile_11_4_1),
		.in_wire_0_2(horizontal_tile_11_5_to_tile_11_4_2),
		.in_wire_0_3(horizontal_tile_11_5_to_tile_11_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(357)
	);

	pe_tile pe_tile_11_5(
		.out_wire_3_0(vertical_tile_11_5_to_tile_10_5_0),
		.out_wire_3_1(vertical_tile_11_5_to_tile_10_5_1),
		.out_wire_3_2(vertical_tile_11_5_to_tile_10_5_2),
		.out_wire_3_3(vertical_tile_11_5_to_tile_10_5_3),
		.in_wire_3_0(vertical_tile_10_5_to_tile_11_5_0),
		.in_wire_3_1(vertical_tile_10_5_to_tile_11_5_1),
		.in_wire_3_2(vertical_tile_10_5_to_tile_11_5_2),
		.in_wire_3_3(vertical_tile_10_5_to_tile_11_5_3),
		.out_wire_1_0(vertical_tile_11_5_to_tile_12_5_0),
		.out_wire_1_1(vertical_tile_11_5_to_tile_12_5_1),
		.out_wire_1_2(vertical_tile_11_5_to_tile_12_5_2),
		.out_wire_1_3(vertical_tile_11_5_to_tile_12_5_3),
		.in_wire_1_0(vertical_tile_12_5_to_tile_11_5_0),
		.in_wire_1_1(vertical_tile_12_5_to_tile_11_5_1),
		.in_wire_1_2(vertical_tile_12_5_to_tile_11_5_2),
		.in_wire_1_3(vertical_tile_12_5_to_tile_11_5_3),
		.out_wire_2_0(horizontal_tile_11_5_to_tile_11_4_0),
		.out_wire_2_1(horizontal_tile_11_5_to_tile_11_4_1),
		.out_wire_2_2(horizontal_tile_11_5_to_tile_11_4_2),
		.out_wire_2_3(horizontal_tile_11_5_to_tile_11_4_3),
		.in_wire_2_0(horizontal_tile_11_4_to_tile_11_5_0),
		.in_wire_2_1(horizontal_tile_11_4_to_tile_11_5_1),
		.in_wire_2_2(horizontal_tile_11_4_to_tile_11_5_2),
		.in_wire_2_3(horizontal_tile_11_4_to_tile_11_5_3),
		.out_wire_0_0(horizontal_tile_11_5_to_tile_11_6_0),
		.out_wire_0_1(horizontal_tile_11_5_to_tile_11_6_1),
		.out_wire_0_2(horizontal_tile_11_5_to_tile_11_6_2),
		.out_wire_0_3(horizontal_tile_11_5_to_tile_11_6_3),
		.in_wire_0_0(horizontal_tile_11_6_to_tile_11_5_0),
		.in_wire_0_1(horizontal_tile_11_6_to_tile_11_5_1),
		.in_wire_0_2(horizontal_tile_11_6_to_tile_11_5_2),
		.in_wire_0_3(horizontal_tile_11_6_to_tile_11_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(358)
	);

	pe_tile pe_tile_11_6(
		.out_wire_3_0(vertical_tile_11_6_to_tile_10_6_0),
		.out_wire_3_1(vertical_tile_11_6_to_tile_10_6_1),
		.out_wire_3_2(vertical_tile_11_6_to_tile_10_6_2),
		.out_wire_3_3(vertical_tile_11_6_to_tile_10_6_3),
		.in_wire_3_0(vertical_tile_10_6_to_tile_11_6_0),
		.in_wire_3_1(vertical_tile_10_6_to_tile_11_6_1),
		.in_wire_3_2(vertical_tile_10_6_to_tile_11_6_2),
		.in_wire_3_3(vertical_tile_10_6_to_tile_11_6_3),
		.out_wire_1_0(vertical_tile_11_6_to_tile_12_6_0),
		.out_wire_1_1(vertical_tile_11_6_to_tile_12_6_1),
		.out_wire_1_2(vertical_tile_11_6_to_tile_12_6_2),
		.out_wire_1_3(vertical_tile_11_6_to_tile_12_6_3),
		.in_wire_1_0(vertical_tile_12_6_to_tile_11_6_0),
		.in_wire_1_1(vertical_tile_12_6_to_tile_11_6_1),
		.in_wire_1_2(vertical_tile_12_6_to_tile_11_6_2),
		.in_wire_1_3(vertical_tile_12_6_to_tile_11_6_3),
		.out_wire_2_0(horizontal_tile_11_6_to_tile_11_5_0),
		.out_wire_2_1(horizontal_tile_11_6_to_tile_11_5_1),
		.out_wire_2_2(horizontal_tile_11_6_to_tile_11_5_2),
		.out_wire_2_3(horizontal_tile_11_6_to_tile_11_5_3),
		.in_wire_2_0(horizontal_tile_11_5_to_tile_11_6_0),
		.in_wire_2_1(horizontal_tile_11_5_to_tile_11_6_1),
		.in_wire_2_2(horizontal_tile_11_5_to_tile_11_6_2),
		.in_wire_2_3(horizontal_tile_11_5_to_tile_11_6_3),
		.out_wire_0_0(horizontal_tile_11_6_to_tile_11_7_0),
		.out_wire_0_1(horizontal_tile_11_6_to_tile_11_7_1),
		.out_wire_0_2(horizontal_tile_11_6_to_tile_11_7_2),
		.out_wire_0_3(horizontal_tile_11_6_to_tile_11_7_3),
		.in_wire_0_0(horizontal_tile_11_7_to_tile_11_6_0),
		.in_wire_0_1(horizontal_tile_11_7_to_tile_11_6_1),
		.in_wire_0_2(horizontal_tile_11_7_to_tile_11_6_2),
		.in_wire_0_3(horizontal_tile_11_7_to_tile_11_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(359)
	);

	pe_tile pe_tile_11_7(
		.out_wire_3_0(vertical_tile_11_7_to_tile_10_7_0),
		.out_wire_3_1(vertical_tile_11_7_to_tile_10_7_1),
		.out_wire_3_2(vertical_tile_11_7_to_tile_10_7_2),
		.out_wire_3_3(vertical_tile_11_7_to_tile_10_7_3),
		.in_wire_3_0(vertical_tile_10_7_to_tile_11_7_0),
		.in_wire_3_1(vertical_tile_10_7_to_tile_11_7_1),
		.in_wire_3_2(vertical_tile_10_7_to_tile_11_7_2),
		.in_wire_3_3(vertical_tile_10_7_to_tile_11_7_3),
		.out_wire_1_0(vertical_tile_11_7_to_tile_12_7_0),
		.out_wire_1_1(vertical_tile_11_7_to_tile_12_7_1),
		.out_wire_1_2(vertical_tile_11_7_to_tile_12_7_2),
		.out_wire_1_3(vertical_tile_11_7_to_tile_12_7_3),
		.in_wire_1_0(vertical_tile_12_7_to_tile_11_7_0),
		.in_wire_1_1(vertical_tile_12_7_to_tile_11_7_1),
		.in_wire_1_2(vertical_tile_12_7_to_tile_11_7_2),
		.in_wire_1_3(vertical_tile_12_7_to_tile_11_7_3),
		.out_wire_2_0(horizontal_tile_11_7_to_tile_11_6_0),
		.out_wire_2_1(horizontal_tile_11_7_to_tile_11_6_1),
		.out_wire_2_2(horizontal_tile_11_7_to_tile_11_6_2),
		.out_wire_2_3(horizontal_tile_11_7_to_tile_11_6_3),
		.in_wire_2_0(horizontal_tile_11_6_to_tile_11_7_0),
		.in_wire_2_1(horizontal_tile_11_6_to_tile_11_7_1),
		.in_wire_2_2(horizontal_tile_11_6_to_tile_11_7_2),
		.in_wire_2_3(horizontal_tile_11_6_to_tile_11_7_3),
		.out_wire_0_0(horizontal_tile_11_7_to_tile_11_8_0),
		.out_wire_0_1(horizontal_tile_11_7_to_tile_11_8_1),
		.out_wire_0_2(horizontal_tile_11_7_to_tile_11_8_2),
		.out_wire_0_3(horizontal_tile_11_7_to_tile_11_8_3),
		.in_wire_0_0(horizontal_tile_11_8_to_tile_11_7_0),
		.in_wire_0_1(horizontal_tile_11_8_to_tile_11_7_1),
		.in_wire_0_2(horizontal_tile_11_8_to_tile_11_7_2),
		.in_wire_0_3(horizontal_tile_11_8_to_tile_11_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(360)
	);

	pe_tile pe_tile_11_8(
		.out_wire_3_0(vertical_tile_11_8_to_tile_10_8_0),
		.out_wire_3_1(vertical_tile_11_8_to_tile_10_8_1),
		.out_wire_3_2(vertical_tile_11_8_to_tile_10_8_2),
		.out_wire_3_3(vertical_tile_11_8_to_tile_10_8_3),
		.in_wire_3_0(vertical_tile_10_8_to_tile_11_8_0),
		.in_wire_3_1(vertical_tile_10_8_to_tile_11_8_1),
		.in_wire_3_2(vertical_tile_10_8_to_tile_11_8_2),
		.in_wire_3_3(vertical_tile_10_8_to_tile_11_8_3),
		.out_wire_1_0(vertical_tile_11_8_to_tile_12_8_0),
		.out_wire_1_1(vertical_tile_11_8_to_tile_12_8_1),
		.out_wire_1_2(vertical_tile_11_8_to_tile_12_8_2),
		.out_wire_1_3(vertical_tile_11_8_to_tile_12_8_3),
		.in_wire_1_0(vertical_tile_12_8_to_tile_11_8_0),
		.in_wire_1_1(vertical_tile_12_8_to_tile_11_8_1),
		.in_wire_1_2(vertical_tile_12_8_to_tile_11_8_2),
		.in_wire_1_3(vertical_tile_12_8_to_tile_11_8_3),
		.out_wire_2_0(horizontal_tile_11_8_to_tile_11_7_0),
		.out_wire_2_1(horizontal_tile_11_8_to_tile_11_7_1),
		.out_wire_2_2(horizontal_tile_11_8_to_tile_11_7_2),
		.out_wire_2_3(horizontal_tile_11_8_to_tile_11_7_3),
		.in_wire_2_0(horizontal_tile_11_7_to_tile_11_8_0),
		.in_wire_2_1(horizontal_tile_11_7_to_tile_11_8_1),
		.in_wire_2_2(horizontal_tile_11_7_to_tile_11_8_2),
		.in_wire_2_3(horizontal_tile_11_7_to_tile_11_8_3),
		.out_wire_0_0(horizontal_tile_11_8_to_tile_11_9_0),
		.out_wire_0_1(horizontal_tile_11_8_to_tile_11_9_1),
		.out_wire_0_2(horizontal_tile_11_8_to_tile_11_9_2),
		.out_wire_0_3(horizontal_tile_11_8_to_tile_11_9_3),
		.in_wire_0_0(horizontal_tile_11_9_to_tile_11_8_0),
		.in_wire_0_1(horizontal_tile_11_9_to_tile_11_8_1),
		.in_wire_0_2(horizontal_tile_11_9_to_tile_11_8_2),
		.in_wire_0_3(horizontal_tile_11_9_to_tile_11_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(361)
	);

	pe_tile pe_tile_11_9(
		.out_wire_3_0(vertical_tile_11_9_to_tile_10_9_0),
		.out_wire_3_1(vertical_tile_11_9_to_tile_10_9_1),
		.out_wire_3_2(vertical_tile_11_9_to_tile_10_9_2),
		.out_wire_3_3(vertical_tile_11_9_to_tile_10_9_3),
		.in_wire_3_0(vertical_tile_10_9_to_tile_11_9_0),
		.in_wire_3_1(vertical_tile_10_9_to_tile_11_9_1),
		.in_wire_3_2(vertical_tile_10_9_to_tile_11_9_2),
		.in_wire_3_3(vertical_tile_10_9_to_tile_11_9_3),
		.out_wire_1_0(vertical_tile_11_9_to_tile_12_9_0),
		.out_wire_1_1(vertical_tile_11_9_to_tile_12_9_1),
		.out_wire_1_2(vertical_tile_11_9_to_tile_12_9_2),
		.out_wire_1_3(vertical_tile_11_9_to_tile_12_9_3),
		.in_wire_1_0(vertical_tile_12_9_to_tile_11_9_0),
		.in_wire_1_1(vertical_tile_12_9_to_tile_11_9_1),
		.in_wire_1_2(vertical_tile_12_9_to_tile_11_9_2),
		.in_wire_1_3(vertical_tile_12_9_to_tile_11_9_3),
		.out_wire_2_0(horizontal_tile_11_9_to_tile_11_8_0),
		.out_wire_2_1(horizontal_tile_11_9_to_tile_11_8_1),
		.out_wire_2_2(horizontal_tile_11_9_to_tile_11_8_2),
		.out_wire_2_3(horizontal_tile_11_9_to_tile_11_8_3),
		.in_wire_2_0(horizontal_tile_11_8_to_tile_11_9_0),
		.in_wire_2_1(horizontal_tile_11_8_to_tile_11_9_1),
		.in_wire_2_2(horizontal_tile_11_8_to_tile_11_9_2),
		.in_wire_2_3(horizontal_tile_11_8_to_tile_11_9_3),
		.out_wire_0_0(horizontal_tile_11_9_to_tile_11_10_0),
		.out_wire_0_1(horizontal_tile_11_9_to_tile_11_10_1),
		.out_wire_0_2(horizontal_tile_11_9_to_tile_11_10_2),
		.out_wire_0_3(horizontal_tile_11_9_to_tile_11_10_3),
		.in_wire_0_0(horizontal_tile_11_10_to_tile_11_9_0),
		.in_wire_0_1(horizontal_tile_11_10_to_tile_11_9_1),
		.in_wire_0_2(horizontal_tile_11_10_to_tile_11_9_2),
		.in_wire_0_3(horizontal_tile_11_10_to_tile_11_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(362)
	);

	pe_tile pe_tile_11_10(
		.out_wire_3_0(vertical_tile_11_10_to_tile_10_10_0),
		.out_wire_3_1(vertical_tile_11_10_to_tile_10_10_1),
		.out_wire_3_2(vertical_tile_11_10_to_tile_10_10_2),
		.out_wire_3_3(vertical_tile_11_10_to_tile_10_10_3),
		.in_wire_3_0(vertical_tile_10_10_to_tile_11_10_0),
		.in_wire_3_1(vertical_tile_10_10_to_tile_11_10_1),
		.in_wire_3_2(vertical_tile_10_10_to_tile_11_10_2),
		.in_wire_3_3(vertical_tile_10_10_to_tile_11_10_3),
		.out_wire_1_0(vertical_tile_11_10_to_tile_12_10_0),
		.out_wire_1_1(vertical_tile_11_10_to_tile_12_10_1),
		.out_wire_1_2(vertical_tile_11_10_to_tile_12_10_2),
		.out_wire_1_3(vertical_tile_11_10_to_tile_12_10_3),
		.in_wire_1_0(vertical_tile_12_10_to_tile_11_10_0),
		.in_wire_1_1(vertical_tile_12_10_to_tile_11_10_1),
		.in_wire_1_2(vertical_tile_12_10_to_tile_11_10_2),
		.in_wire_1_3(vertical_tile_12_10_to_tile_11_10_3),
		.out_wire_2_0(horizontal_tile_11_10_to_tile_11_9_0),
		.out_wire_2_1(horizontal_tile_11_10_to_tile_11_9_1),
		.out_wire_2_2(horizontal_tile_11_10_to_tile_11_9_2),
		.out_wire_2_3(horizontal_tile_11_10_to_tile_11_9_3),
		.in_wire_2_0(horizontal_tile_11_9_to_tile_11_10_0),
		.in_wire_2_1(horizontal_tile_11_9_to_tile_11_10_1),
		.in_wire_2_2(horizontal_tile_11_9_to_tile_11_10_2),
		.in_wire_2_3(horizontal_tile_11_9_to_tile_11_10_3),
		.out_wire_0_0(horizontal_tile_11_10_to_tile_11_11_0),
		.out_wire_0_1(horizontal_tile_11_10_to_tile_11_11_1),
		.out_wire_0_2(horizontal_tile_11_10_to_tile_11_11_2),
		.out_wire_0_3(horizontal_tile_11_10_to_tile_11_11_3),
		.in_wire_0_0(horizontal_tile_11_11_to_tile_11_10_0),
		.in_wire_0_1(horizontal_tile_11_11_to_tile_11_10_1),
		.in_wire_0_2(horizontal_tile_11_11_to_tile_11_10_2),
		.in_wire_0_3(horizontal_tile_11_11_to_tile_11_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(363)
	);

	pe_tile pe_tile_11_11(
		.out_wire_3_0(vertical_tile_11_11_to_tile_10_11_0),
		.out_wire_3_1(vertical_tile_11_11_to_tile_10_11_1),
		.out_wire_3_2(vertical_tile_11_11_to_tile_10_11_2),
		.out_wire_3_3(vertical_tile_11_11_to_tile_10_11_3),
		.in_wire_3_0(vertical_tile_10_11_to_tile_11_11_0),
		.in_wire_3_1(vertical_tile_10_11_to_tile_11_11_1),
		.in_wire_3_2(vertical_tile_10_11_to_tile_11_11_2),
		.in_wire_3_3(vertical_tile_10_11_to_tile_11_11_3),
		.out_wire_1_0(vertical_tile_11_11_to_tile_12_11_0),
		.out_wire_1_1(vertical_tile_11_11_to_tile_12_11_1),
		.out_wire_1_2(vertical_tile_11_11_to_tile_12_11_2),
		.out_wire_1_3(vertical_tile_11_11_to_tile_12_11_3),
		.in_wire_1_0(vertical_tile_12_11_to_tile_11_11_0),
		.in_wire_1_1(vertical_tile_12_11_to_tile_11_11_1),
		.in_wire_1_2(vertical_tile_12_11_to_tile_11_11_2),
		.in_wire_1_3(vertical_tile_12_11_to_tile_11_11_3),
		.out_wire_2_0(horizontal_tile_11_11_to_tile_11_10_0),
		.out_wire_2_1(horizontal_tile_11_11_to_tile_11_10_1),
		.out_wire_2_2(horizontal_tile_11_11_to_tile_11_10_2),
		.out_wire_2_3(horizontal_tile_11_11_to_tile_11_10_3),
		.in_wire_2_0(horizontal_tile_11_10_to_tile_11_11_0),
		.in_wire_2_1(horizontal_tile_11_10_to_tile_11_11_1),
		.in_wire_2_2(horizontal_tile_11_10_to_tile_11_11_2),
		.in_wire_2_3(horizontal_tile_11_10_to_tile_11_11_3),
		.out_wire_0_0(horizontal_tile_11_11_to_tile_11_12_0),
		.out_wire_0_1(horizontal_tile_11_11_to_tile_11_12_1),
		.out_wire_0_2(horizontal_tile_11_11_to_tile_11_12_2),
		.out_wire_0_3(horizontal_tile_11_11_to_tile_11_12_3),
		.in_wire_0_0(horizontal_tile_11_12_to_tile_11_11_0),
		.in_wire_0_1(horizontal_tile_11_12_to_tile_11_11_1),
		.in_wire_0_2(horizontal_tile_11_12_to_tile_11_11_2),
		.in_wire_0_3(horizontal_tile_11_12_to_tile_11_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(364)
	);

	pe_tile pe_tile_11_12(
		.out_wire_3_0(vertical_tile_11_12_to_tile_10_12_0),
		.out_wire_3_1(vertical_tile_11_12_to_tile_10_12_1),
		.out_wire_3_2(vertical_tile_11_12_to_tile_10_12_2),
		.out_wire_3_3(vertical_tile_11_12_to_tile_10_12_3),
		.in_wire_3_0(vertical_tile_10_12_to_tile_11_12_0),
		.in_wire_3_1(vertical_tile_10_12_to_tile_11_12_1),
		.in_wire_3_2(vertical_tile_10_12_to_tile_11_12_2),
		.in_wire_3_3(vertical_tile_10_12_to_tile_11_12_3),
		.out_wire_1_0(vertical_tile_11_12_to_tile_12_12_0),
		.out_wire_1_1(vertical_tile_11_12_to_tile_12_12_1),
		.out_wire_1_2(vertical_tile_11_12_to_tile_12_12_2),
		.out_wire_1_3(vertical_tile_11_12_to_tile_12_12_3),
		.in_wire_1_0(vertical_tile_12_12_to_tile_11_12_0),
		.in_wire_1_1(vertical_tile_12_12_to_tile_11_12_1),
		.in_wire_1_2(vertical_tile_12_12_to_tile_11_12_2),
		.in_wire_1_3(vertical_tile_12_12_to_tile_11_12_3),
		.out_wire_2_0(horizontal_tile_11_12_to_tile_11_11_0),
		.out_wire_2_1(horizontal_tile_11_12_to_tile_11_11_1),
		.out_wire_2_2(horizontal_tile_11_12_to_tile_11_11_2),
		.out_wire_2_3(horizontal_tile_11_12_to_tile_11_11_3),
		.in_wire_2_0(horizontal_tile_11_11_to_tile_11_12_0),
		.in_wire_2_1(horizontal_tile_11_11_to_tile_11_12_1),
		.in_wire_2_2(horizontal_tile_11_11_to_tile_11_12_2),
		.in_wire_2_3(horizontal_tile_11_11_to_tile_11_12_3),
		.out_wire_0_0(horizontal_tile_11_12_to_tile_11_13_0),
		.out_wire_0_1(horizontal_tile_11_12_to_tile_11_13_1),
		.out_wire_0_2(horizontal_tile_11_12_to_tile_11_13_2),
		.out_wire_0_3(horizontal_tile_11_12_to_tile_11_13_3),
		.in_wire_0_0(horizontal_tile_11_13_to_tile_11_12_0),
		.in_wire_0_1(horizontal_tile_11_13_to_tile_11_12_1),
		.in_wire_0_2(horizontal_tile_11_13_to_tile_11_12_2),
		.in_wire_0_3(horizontal_tile_11_13_to_tile_11_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(365)
	);

	pe_tile pe_tile_11_13(
		.out_wire_3_0(vertical_tile_11_13_to_tile_10_13_0),
		.out_wire_3_1(vertical_tile_11_13_to_tile_10_13_1),
		.out_wire_3_2(vertical_tile_11_13_to_tile_10_13_2),
		.out_wire_3_3(vertical_tile_11_13_to_tile_10_13_3),
		.in_wire_3_0(vertical_tile_10_13_to_tile_11_13_0),
		.in_wire_3_1(vertical_tile_10_13_to_tile_11_13_1),
		.in_wire_3_2(vertical_tile_10_13_to_tile_11_13_2),
		.in_wire_3_3(vertical_tile_10_13_to_tile_11_13_3),
		.out_wire_1_0(vertical_tile_11_13_to_tile_12_13_0),
		.out_wire_1_1(vertical_tile_11_13_to_tile_12_13_1),
		.out_wire_1_2(vertical_tile_11_13_to_tile_12_13_2),
		.out_wire_1_3(vertical_tile_11_13_to_tile_12_13_3),
		.in_wire_1_0(vertical_tile_12_13_to_tile_11_13_0),
		.in_wire_1_1(vertical_tile_12_13_to_tile_11_13_1),
		.in_wire_1_2(vertical_tile_12_13_to_tile_11_13_2),
		.in_wire_1_3(vertical_tile_12_13_to_tile_11_13_3),
		.out_wire_2_0(horizontal_tile_11_13_to_tile_11_12_0),
		.out_wire_2_1(horizontal_tile_11_13_to_tile_11_12_1),
		.out_wire_2_2(horizontal_tile_11_13_to_tile_11_12_2),
		.out_wire_2_3(horizontal_tile_11_13_to_tile_11_12_3),
		.in_wire_2_0(horizontal_tile_11_12_to_tile_11_13_0),
		.in_wire_2_1(horizontal_tile_11_12_to_tile_11_13_1),
		.in_wire_2_2(horizontal_tile_11_12_to_tile_11_13_2),
		.in_wire_2_3(horizontal_tile_11_12_to_tile_11_13_3),
		.out_wire_0_0(horizontal_tile_11_13_to_tile_11_14_0),
		.out_wire_0_1(horizontal_tile_11_13_to_tile_11_14_1),
		.out_wire_0_2(horizontal_tile_11_13_to_tile_11_14_2),
		.out_wire_0_3(horizontal_tile_11_13_to_tile_11_14_3),
		.in_wire_0_0(horizontal_tile_11_14_to_tile_11_13_0),
		.in_wire_0_1(horizontal_tile_11_14_to_tile_11_13_1),
		.in_wire_0_2(horizontal_tile_11_14_to_tile_11_13_2),
		.in_wire_0_3(horizontal_tile_11_14_to_tile_11_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(366)
	);

	pe_tile pe_tile_11_14(
		.out_wire_3_0(vertical_tile_11_14_to_tile_10_14_0),
		.out_wire_3_1(vertical_tile_11_14_to_tile_10_14_1),
		.out_wire_3_2(vertical_tile_11_14_to_tile_10_14_2),
		.out_wire_3_3(vertical_tile_11_14_to_tile_10_14_3),
		.in_wire_3_0(vertical_tile_10_14_to_tile_11_14_0),
		.in_wire_3_1(vertical_tile_10_14_to_tile_11_14_1),
		.in_wire_3_2(vertical_tile_10_14_to_tile_11_14_2),
		.in_wire_3_3(vertical_tile_10_14_to_tile_11_14_3),
		.out_wire_1_0(vertical_tile_11_14_to_tile_12_14_0),
		.out_wire_1_1(vertical_tile_11_14_to_tile_12_14_1),
		.out_wire_1_2(vertical_tile_11_14_to_tile_12_14_2),
		.out_wire_1_3(vertical_tile_11_14_to_tile_12_14_3),
		.in_wire_1_0(vertical_tile_12_14_to_tile_11_14_0),
		.in_wire_1_1(vertical_tile_12_14_to_tile_11_14_1),
		.in_wire_1_2(vertical_tile_12_14_to_tile_11_14_2),
		.in_wire_1_3(vertical_tile_12_14_to_tile_11_14_3),
		.out_wire_2_0(horizontal_tile_11_14_to_tile_11_13_0),
		.out_wire_2_1(horizontal_tile_11_14_to_tile_11_13_1),
		.out_wire_2_2(horizontal_tile_11_14_to_tile_11_13_2),
		.out_wire_2_3(horizontal_tile_11_14_to_tile_11_13_3),
		.in_wire_2_0(horizontal_tile_11_13_to_tile_11_14_0),
		.in_wire_2_1(horizontal_tile_11_13_to_tile_11_14_1),
		.in_wire_2_2(horizontal_tile_11_13_to_tile_11_14_2),
		.in_wire_2_3(horizontal_tile_11_13_to_tile_11_14_3),
		.out_wire_0_0(horizontal_tile_11_14_to_tile_11_15_0),
		.out_wire_0_1(horizontal_tile_11_14_to_tile_11_15_1),
		.out_wire_0_2(horizontal_tile_11_14_to_tile_11_15_2),
		.out_wire_0_3(horizontal_tile_11_14_to_tile_11_15_3),
		.in_wire_0_0(horizontal_tile_11_15_to_tile_11_14_0),
		.in_wire_0_1(horizontal_tile_11_15_to_tile_11_14_1),
		.in_wire_0_2(horizontal_tile_11_15_to_tile_11_14_2),
		.in_wire_0_3(horizontal_tile_11_15_to_tile_11_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(367)
	);

	pe_tile pe_tile_11_15(
		.out_wire_3_0(vertical_tile_11_15_to_tile_10_15_0),
		.out_wire_3_1(vertical_tile_11_15_to_tile_10_15_1),
		.out_wire_3_2(vertical_tile_11_15_to_tile_10_15_2),
		.out_wire_3_3(vertical_tile_11_15_to_tile_10_15_3),
		.in_wire_3_0(vertical_tile_10_15_to_tile_11_15_0),
		.in_wire_3_1(vertical_tile_10_15_to_tile_11_15_1),
		.in_wire_3_2(vertical_tile_10_15_to_tile_11_15_2),
		.in_wire_3_3(vertical_tile_10_15_to_tile_11_15_3),
		.out_wire_1_0(vertical_tile_11_15_to_tile_12_15_0),
		.out_wire_1_1(vertical_tile_11_15_to_tile_12_15_1),
		.out_wire_1_2(vertical_tile_11_15_to_tile_12_15_2),
		.out_wire_1_3(vertical_tile_11_15_to_tile_12_15_3),
		.in_wire_1_0(vertical_tile_12_15_to_tile_11_15_0),
		.in_wire_1_1(vertical_tile_12_15_to_tile_11_15_1),
		.in_wire_1_2(vertical_tile_12_15_to_tile_11_15_2),
		.in_wire_1_3(vertical_tile_12_15_to_tile_11_15_3),
		.out_wire_2_0(horizontal_tile_11_15_to_tile_11_14_0),
		.out_wire_2_1(horizontal_tile_11_15_to_tile_11_14_1),
		.out_wire_2_2(horizontal_tile_11_15_to_tile_11_14_2),
		.out_wire_2_3(horizontal_tile_11_15_to_tile_11_14_3),
		.in_wire_2_0(horizontal_tile_11_14_to_tile_11_15_0),
		.in_wire_2_1(horizontal_tile_11_14_to_tile_11_15_1),
		.in_wire_2_2(horizontal_tile_11_14_to_tile_11_15_2),
		.in_wire_2_3(horizontal_tile_11_14_to_tile_11_15_3),
		.out_wire_0_0(horizontal_tile_11_15_to_tile_11_16_0),
		.out_wire_0_1(horizontal_tile_11_15_to_tile_11_16_1),
		.out_wire_0_2(horizontal_tile_11_15_to_tile_11_16_2),
		.out_wire_0_3(horizontal_tile_11_15_to_tile_11_16_3),
		.in_wire_0_0(horizontal_tile_11_16_to_tile_11_15_0),
		.in_wire_0_1(horizontal_tile_11_16_to_tile_11_15_1),
		.in_wire_0_2(horizontal_tile_11_16_to_tile_11_15_2),
		.in_wire_0_3(horizontal_tile_11_16_to_tile_11_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(368)
	);

	pe_tile pe_tile_11_16(
		.out_wire_3_0(vertical_tile_11_16_to_tile_10_16_0),
		.out_wire_3_1(vertical_tile_11_16_to_tile_10_16_1),
		.out_wire_3_2(vertical_tile_11_16_to_tile_10_16_2),
		.out_wire_3_3(vertical_tile_11_16_to_tile_10_16_3),
		.in_wire_3_0(vertical_tile_10_16_to_tile_11_16_0),
		.in_wire_3_1(vertical_tile_10_16_to_tile_11_16_1),
		.in_wire_3_2(vertical_tile_10_16_to_tile_11_16_2),
		.in_wire_3_3(vertical_tile_10_16_to_tile_11_16_3),
		.out_wire_1_0(vertical_tile_11_16_to_tile_12_16_0),
		.out_wire_1_1(vertical_tile_11_16_to_tile_12_16_1),
		.out_wire_1_2(vertical_tile_11_16_to_tile_12_16_2),
		.out_wire_1_3(vertical_tile_11_16_to_tile_12_16_3),
		.in_wire_1_0(vertical_tile_12_16_to_tile_11_16_0),
		.in_wire_1_1(vertical_tile_12_16_to_tile_11_16_1),
		.in_wire_1_2(vertical_tile_12_16_to_tile_11_16_2),
		.in_wire_1_3(vertical_tile_12_16_to_tile_11_16_3),
		.out_wire_2_0(horizontal_tile_11_16_to_tile_11_15_0),
		.out_wire_2_1(horizontal_tile_11_16_to_tile_11_15_1),
		.out_wire_2_2(horizontal_tile_11_16_to_tile_11_15_2),
		.out_wire_2_3(horizontal_tile_11_16_to_tile_11_15_3),
		.in_wire_2_0(horizontal_tile_11_15_to_tile_11_16_0),
		.in_wire_2_1(horizontal_tile_11_15_to_tile_11_16_1),
		.in_wire_2_2(horizontal_tile_11_15_to_tile_11_16_2),
		.in_wire_2_3(horizontal_tile_11_15_to_tile_11_16_3),
		.out_wire_0_0(horizontal_tile_11_16_to_tile_11_17_0),
		.out_wire_0_1(horizontal_tile_11_16_to_tile_11_17_1),
		.out_wire_0_2(horizontal_tile_11_16_to_tile_11_17_2),
		.out_wire_0_3(horizontal_tile_11_16_to_tile_11_17_3),
		.in_wire_0_0(horizontal_tile_11_17_to_tile_11_16_0),
		.in_wire_0_1(horizontal_tile_11_17_to_tile_11_16_1),
		.in_wire_0_2(horizontal_tile_11_17_to_tile_11_16_2),
		.in_wire_0_3(horizontal_tile_11_17_to_tile_11_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(369)
	);

	pe_tile pe_tile_11_17(
		.out_wire_3_0(vertical_tile_11_17_to_tile_10_17_0),
		.out_wire_3_1(vertical_tile_11_17_to_tile_10_17_1),
		.out_wire_3_2(vertical_tile_11_17_to_tile_10_17_2),
		.out_wire_3_3(vertical_tile_11_17_to_tile_10_17_3),
		.in_wire_3_0(vertical_tile_10_17_to_tile_11_17_0),
		.in_wire_3_1(vertical_tile_10_17_to_tile_11_17_1),
		.in_wire_3_2(vertical_tile_10_17_to_tile_11_17_2),
		.in_wire_3_3(vertical_tile_10_17_to_tile_11_17_3),
		.out_wire_1_0(vertical_tile_11_17_to_tile_12_17_0),
		.out_wire_1_1(vertical_tile_11_17_to_tile_12_17_1),
		.out_wire_1_2(vertical_tile_11_17_to_tile_12_17_2),
		.out_wire_1_3(vertical_tile_11_17_to_tile_12_17_3),
		.in_wire_1_0(vertical_tile_12_17_to_tile_11_17_0),
		.in_wire_1_1(vertical_tile_12_17_to_tile_11_17_1),
		.in_wire_1_2(vertical_tile_12_17_to_tile_11_17_2),
		.in_wire_1_3(vertical_tile_12_17_to_tile_11_17_3),
		.out_wire_2_0(horizontal_tile_11_17_to_tile_11_16_0),
		.out_wire_2_1(horizontal_tile_11_17_to_tile_11_16_1),
		.out_wire_2_2(horizontal_tile_11_17_to_tile_11_16_2),
		.out_wire_2_3(horizontal_tile_11_17_to_tile_11_16_3),
		.in_wire_2_0(horizontal_tile_11_16_to_tile_11_17_0),
		.in_wire_2_1(horizontal_tile_11_16_to_tile_11_17_1),
		.in_wire_2_2(horizontal_tile_11_16_to_tile_11_17_2),
		.in_wire_2_3(horizontal_tile_11_16_to_tile_11_17_3),
		.out_wire_0_0(horizontal_tile_11_17_to_tile_11_18_0),
		.out_wire_0_1(horizontal_tile_11_17_to_tile_11_18_1),
		.out_wire_0_2(horizontal_tile_11_17_to_tile_11_18_2),
		.out_wire_0_3(horizontal_tile_11_17_to_tile_11_18_3),
		.in_wire_0_0(horizontal_tile_11_18_to_tile_11_17_0),
		.in_wire_0_1(horizontal_tile_11_18_to_tile_11_17_1),
		.in_wire_0_2(horizontal_tile_11_18_to_tile_11_17_2),
		.in_wire_0_3(horizontal_tile_11_18_to_tile_11_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(370)
	);

	pe_tile pe_tile_11_18(
		.out_wire_3_0(vertical_tile_11_18_to_tile_10_18_0),
		.out_wire_3_1(vertical_tile_11_18_to_tile_10_18_1),
		.out_wire_3_2(vertical_tile_11_18_to_tile_10_18_2),
		.out_wire_3_3(vertical_tile_11_18_to_tile_10_18_3),
		.in_wire_3_0(vertical_tile_10_18_to_tile_11_18_0),
		.in_wire_3_1(vertical_tile_10_18_to_tile_11_18_1),
		.in_wire_3_2(vertical_tile_10_18_to_tile_11_18_2),
		.in_wire_3_3(vertical_tile_10_18_to_tile_11_18_3),
		.out_wire_1_0(vertical_tile_11_18_to_tile_12_18_0),
		.out_wire_1_1(vertical_tile_11_18_to_tile_12_18_1),
		.out_wire_1_2(vertical_tile_11_18_to_tile_12_18_2),
		.out_wire_1_3(vertical_tile_11_18_to_tile_12_18_3),
		.in_wire_1_0(vertical_tile_12_18_to_tile_11_18_0),
		.in_wire_1_1(vertical_tile_12_18_to_tile_11_18_1),
		.in_wire_1_2(vertical_tile_12_18_to_tile_11_18_2),
		.in_wire_1_3(vertical_tile_12_18_to_tile_11_18_3),
		.out_wire_2_0(horizontal_tile_11_18_to_tile_11_17_0),
		.out_wire_2_1(horizontal_tile_11_18_to_tile_11_17_1),
		.out_wire_2_2(horizontal_tile_11_18_to_tile_11_17_2),
		.out_wire_2_3(horizontal_tile_11_18_to_tile_11_17_3),
		.in_wire_2_0(horizontal_tile_11_17_to_tile_11_18_0),
		.in_wire_2_1(horizontal_tile_11_17_to_tile_11_18_1),
		.in_wire_2_2(horizontal_tile_11_17_to_tile_11_18_2),
		.in_wire_2_3(horizontal_tile_11_17_to_tile_11_18_3),
		.out_wire_0_0(horizontal_tile_11_18_to_tile_11_19_0),
		.out_wire_0_1(horizontal_tile_11_18_to_tile_11_19_1),
		.out_wire_0_2(horizontal_tile_11_18_to_tile_11_19_2),
		.out_wire_0_3(horizontal_tile_11_18_to_tile_11_19_3),
		.in_wire_0_0(horizontal_tile_11_19_to_tile_11_18_0),
		.in_wire_0_1(horizontal_tile_11_19_to_tile_11_18_1),
		.in_wire_0_2(horizontal_tile_11_19_to_tile_11_18_2),
		.in_wire_0_3(horizontal_tile_11_19_to_tile_11_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(371)
	);

	pe_tile pe_tile_11_19(
		.out_wire_3_0(vertical_tile_11_19_to_tile_10_19_0),
		.out_wire_3_1(vertical_tile_11_19_to_tile_10_19_1),
		.out_wire_3_2(vertical_tile_11_19_to_tile_10_19_2),
		.out_wire_3_3(vertical_tile_11_19_to_tile_10_19_3),
		.in_wire_3_0(vertical_tile_10_19_to_tile_11_19_0),
		.in_wire_3_1(vertical_tile_10_19_to_tile_11_19_1),
		.in_wire_3_2(vertical_tile_10_19_to_tile_11_19_2),
		.in_wire_3_3(vertical_tile_10_19_to_tile_11_19_3),
		.out_wire_1_0(vertical_tile_11_19_to_tile_12_19_0),
		.out_wire_1_1(vertical_tile_11_19_to_tile_12_19_1),
		.out_wire_1_2(vertical_tile_11_19_to_tile_12_19_2),
		.out_wire_1_3(vertical_tile_11_19_to_tile_12_19_3),
		.in_wire_1_0(vertical_tile_12_19_to_tile_11_19_0),
		.in_wire_1_1(vertical_tile_12_19_to_tile_11_19_1),
		.in_wire_1_2(vertical_tile_12_19_to_tile_11_19_2),
		.in_wire_1_3(vertical_tile_12_19_to_tile_11_19_3),
		.out_wire_2_0(horizontal_tile_11_19_to_tile_11_18_0),
		.out_wire_2_1(horizontal_tile_11_19_to_tile_11_18_1),
		.out_wire_2_2(horizontal_tile_11_19_to_tile_11_18_2),
		.out_wire_2_3(horizontal_tile_11_19_to_tile_11_18_3),
		.in_wire_2_0(horizontal_tile_11_18_to_tile_11_19_0),
		.in_wire_2_1(horizontal_tile_11_18_to_tile_11_19_1),
		.in_wire_2_2(horizontal_tile_11_18_to_tile_11_19_2),
		.in_wire_2_3(horizontal_tile_11_18_to_tile_11_19_3),
		.out_wire_0_0(horizontal_tile_11_19_to_tile_11_20_0),
		.out_wire_0_1(horizontal_tile_11_19_to_tile_11_20_1),
		.out_wire_0_2(horizontal_tile_11_19_to_tile_11_20_2),
		.out_wire_0_3(horizontal_tile_11_19_to_tile_11_20_3),
		.in_wire_0_0(horizontal_tile_11_20_to_tile_11_19_0),
		.in_wire_0_1(horizontal_tile_11_20_to_tile_11_19_1),
		.in_wire_0_2(horizontal_tile_11_20_to_tile_11_19_2),
		.in_wire_0_3(horizontal_tile_11_20_to_tile_11_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(372)
	);

	pe_tile pe_tile_11_20(
		.out_wire_3_0(vertical_tile_11_20_to_tile_10_20_0),
		.out_wire_3_1(vertical_tile_11_20_to_tile_10_20_1),
		.out_wire_3_2(vertical_tile_11_20_to_tile_10_20_2),
		.out_wire_3_3(vertical_tile_11_20_to_tile_10_20_3),
		.in_wire_3_0(vertical_tile_10_20_to_tile_11_20_0),
		.in_wire_3_1(vertical_tile_10_20_to_tile_11_20_1),
		.in_wire_3_2(vertical_tile_10_20_to_tile_11_20_2),
		.in_wire_3_3(vertical_tile_10_20_to_tile_11_20_3),
		.out_wire_1_0(vertical_tile_11_20_to_tile_12_20_0),
		.out_wire_1_1(vertical_tile_11_20_to_tile_12_20_1),
		.out_wire_1_2(vertical_tile_11_20_to_tile_12_20_2),
		.out_wire_1_3(vertical_tile_11_20_to_tile_12_20_3),
		.in_wire_1_0(vertical_tile_12_20_to_tile_11_20_0),
		.in_wire_1_1(vertical_tile_12_20_to_tile_11_20_1),
		.in_wire_1_2(vertical_tile_12_20_to_tile_11_20_2),
		.in_wire_1_3(vertical_tile_12_20_to_tile_11_20_3),
		.out_wire_2_0(horizontal_tile_11_20_to_tile_11_19_0),
		.out_wire_2_1(horizontal_tile_11_20_to_tile_11_19_1),
		.out_wire_2_2(horizontal_tile_11_20_to_tile_11_19_2),
		.out_wire_2_3(horizontal_tile_11_20_to_tile_11_19_3),
		.in_wire_2_0(horizontal_tile_11_19_to_tile_11_20_0),
		.in_wire_2_1(horizontal_tile_11_19_to_tile_11_20_1),
		.in_wire_2_2(horizontal_tile_11_19_to_tile_11_20_2),
		.in_wire_2_3(horizontal_tile_11_19_to_tile_11_20_3),
		.out_wire_0_0(horizontal_tile_11_20_to_tile_11_21_0),
		.out_wire_0_1(horizontal_tile_11_20_to_tile_11_21_1),
		.out_wire_0_2(horizontal_tile_11_20_to_tile_11_21_2),
		.out_wire_0_3(horizontal_tile_11_20_to_tile_11_21_3),
		.in_wire_0_0(horizontal_tile_11_21_to_tile_11_20_0),
		.in_wire_0_1(horizontal_tile_11_21_to_tile_11_20_1),
		.in_wire_0_2(horizontal_tile_11_21_to_tile_11_20_2),
		.in_wire_0_3(horizontal_tile_11_21_to_tile_11_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(373)
	);

	pe_tile pe_tile_11_21(
		.out_wire_3_0(vertical_tile_11_21_to_tile_10_21_0),
		.out_wire_3_1(vertical_tile_11_21_to_tile_10_21_1),
		.out_wire_3_2(vertical_tile_11_21_to_tile_10_21_2),
		.out_wire_3_3(vertical_tile_11_21_to_tile_10_21_3),
		.in_wire_3_0(vertical_tile_10_21_to_tile_11_21_0),
		.in_wire_3_1(vertical_tile_10_21_to_tile_11_21_1),
		.in_wire_3_2(vertical_tile_10_21_to_tile_11_21_2),
		.in_wire_3_3(vertical_tile_10_21_to_tile_11_21_3),
		.out_wire_1_0(vertical_tile_11_21_to_tile_12_21_0),
		.out_wire_1_1(vertical_tile_11_21_to_tile_12_21_1),
		.out_wire_1_2(vertical_tile_11_21_to_tile_12_21_2),
		.out_wire_1_3(vertical_tile_11_21_to_tile_12_21_3),
		.in_wire_1_0(vertical_tile_12_21_to_tile_11_21_0),
		.in_wire_1_1(vertical_tile_12_21_to_tile_11_21_1),
		.in_wire_1_2(vertical_tile_12_21_to_tile_11_21_2),
		.in_wire_1_3(vertical_tile_12_21_to_tile_11_21_3),
		.out_wire_2_0(horizontal_tile_11_21_to_tile_11_20_0),
		.out_wire_2_1(horizontal_tile_11_21_to_tile_11_20_1),
		.out_wire_2_2(horizontal_tile_11_21_to_tile_11_20_2),
		.out_wire_2_3(horizontal_tile_11_21_to_tile_11_20_3),
		.in_wire_2_0(horizontal_tile_11_20_to_tile_11_21_0),
		.in_wire_2_1(horizontal_tile_11_20_to_tile_11_21_1),
		.in_wire_2_2(horizontal_tile_11_20_to_tile_11_21_2),
		.in_wire_2_3(horizontal_tile_11_20_to_tile_11_21_3),
		.out_wire_0_0(horizontal_tile_11_21_to_tile_11_22_0),
		.out_wire_0_1(horizontal_tile_11_21_to_tile_11_22_1),
		.out_wire_0_2(horizontal_tile_11_21_to_tile_11_22_2),
		.out_wire_0_3(horizontal_tile_11_21_to_tile_11_22_3),
		.in_wire_0_0(horizontal_tile_11_22_to_tile_11_21_0),
		.in_wire_0_1(horizontal_tile_11_22_to_tile_11_21_1),
		.in_wire_0_2(horizontal_tile_11_22_to_tile_11_21_2),
		.in_wire_0_3(horizontal_tile_11_22_to_tile_11_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(374)
	);

	pe_tile pe_tile_11_22(
		.out_wire_3_0(vertical_tile_11_22_to_tile_10_22_0),
		.out_wire_3_1(vertical_tile_11_22_to_tile_10_22_1),
		.out_wire_3_2(vertical_tile_11_22_to_tile_10_22_2),
		.out_wire_3_3(vertical_tile_11_22_to_tile_10_22_3),
		.in_wire_3_0(vertical_tile_10_22_to_tile_11_22_0),
		.in_wire_3_1(vertical_tile_10_22_to_tile_11_22_1),
		.in_wire_3_2(vertical_tile_10_22_to_tile_11_22_2),
		.in_wire_3_3(vertical_tile_10_22_to_tile_11_22_3),
		.out_wire_1_0(vertical_tile_11_22_to_tile_12_22_0),
		.out_wire_1_1(vertical_tile_11_22_to_tile_12_22_1),
		.out_wire_1_2(vertical_tile_11_22_to_tile_12_22_2),
		.out_wire_1_3(vertical_tile_11_22_to_tile_12_22_3),
		.in_wire_1_0(vertical_tile_12_22_to_tile_11_22_0),
		.in_wire_1_1(vertical_tile_12_22_to_tile_11_22_1),
		.in_wire_1_2(vertical_tile_12_22_to_tile_11_22_2),
		.in_wire_1_3(vertical_tile_12_22_to_tile_11_22_3),
		.out_wire_2_0(horizontal_tile_11_22_to_tile_11_21_0),
		.out_wire_2_1(horizontal_tile_11_22_to_tile_11_21_1),
		.out_wire_2_2(horizontal_tile_11_22_to_tile_11_21_2),
		.out_wire_2_3(horizontal_tile_11_22_to_tile_11_21_3),
		.in_wire_2_0(horizontal_tile_11_21_to_tile_11_22_0),
		.in_wire_2_1(horizontal_tile_11_21_to_tile_11_22_1),
		.in_wire_2_2(horizontal_tile_11_21_to_tile_11_22_2),
		.in_wire_2_3(horizontal_tile_11_21_to_tile_11_22_3),
		.out_wire_0_0(horizontal_tile_11_22_to_tile_11_23_0),
		.out_wire_0_1(horizontal_tile_11_22_to_tile_11_23_1),
		.out_wire_0_2(horizontal_tile_11_22_to_tile_11_23_2),
		.out_wire_0_3(horizontal_tile_11_22_to_tile_11_23_3),
		.in_wire_0_0(horizontal_tile_11_23_to_tile_11_22_0),
		.in_wire_0_1(horizontal_tile_11_23_to_tile_11_22_1),
		.in_wire_0_2(horizontal_tile_11_23_to_tile_11_22_2),
		.in_wire_0_3(horizontal_tile_11_23_to_tile_11_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(375)
	);

	pe_tile pe_tile_11_23(
		.out_wire_3_0(vertical_tile_11_23_to_tile_10_23_0),
		.out_wire_3_1(vertical_tile_11_23_to_tile_10_23_1),
		.out_wire_3_2(vertical_tile_11_23_to_tile_10_23_2),
		.out_wire_3_3(vertical_tile_11_23_to_tile_10_23_3),
		.in_wire_3_0(vertical_tile_10_23_to_tile_11_23_0),
		.in_wire_3_1(vertical_tile_10_23_to_tile_11_23_1),
		.in_wire_3_2(vertical_tile_10_23_to_tile_11_23_2),
		.in_wire_3_3(vertical_tile_10_23_to_tile_11_23_3),
		.out_wire_1_0(vertical_tile_11_23_to_tile_12_23_0),
		.out_wire_1_1(vertical_tile_11_23_to_tile_12_23_1),
		.out_wire_1_2(vertical_tile_11_23_to_tile_12_23_2),
		.out_wire_1_3(vertical_tile_11_23_to_tile_12_23_3),
		.in_wire_1_0(vertical_tile_12_23_to_tile_11_23_0),
		.in_wire_1_1(vertical_tile_12_23_to_tile_11_23_1),
		.in_wire_1_2(vertical_tile_12_23_to_tile_11_23_2),
		.in_wire_1_3(vertical_tile_12_23_to_tile_11_23_3),
		.out_wire_2_0(horizontal_tile_11_23_to_tile_11_22_0),
		.out_wire_2_1(horizontal_tile_11_23_to_tile_11_22_1),
		.out_wire_2_2(horizontal_tile_11_23_to_tile_11_22_2),
		.out_wire_2_3(horizontal_tile_11_23_to_tile_11_22_3),
		.in_wire_2_0(horizontal_tile_11_22_to_tile_11_23_0),
		.in_wire_2_1(horizontal_tile_11_22_to_tile_11_23_1),
		.in_wire_2_2(horizontal_tile_11_22_to_tile_11_23_2),
		.in_wire_2_3(horizontal_tile_11_22_to_tile_11_23_3),
		.out_wire_0_0(horizontal_tile_11_23_to_tile_11_24_0),
		.out_wire_0_1(horizontal_tile_11_23_to_tile_11_24_1),
		.out_wire_0_2(horizontal_tile_11_23_to_tile_11_24_2),
		.out_wire_0_3(horizontal_tile_11_23_to_tile_11_24_3),
		.in_wire_0_0(horizontal_tile_11_24_to_tile_11_23_0),
		.in_wire_0_1(horizontal_tile_11_24_to_tile_11_23_1),
		.in_wire_0_2(horizontal_tile_11_24_to_tile_11_23_2),
		.in_wire_0_3(horizontal_tile_11_24_to_tile_11_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(376)
	);

	pe_tile pe_tile_11_24(
		.out_wire_3_0(vertical_tile_11_24_to_tile_10_24_0),
		.out_wire_3_1(vertical_tile_11_24_to_tile_10_24_1),
		.out_wire_3_2(vertical_tile_11_24_to_tile_10_24_2),
		.out_wire_3_3(vertical_tile_11_24_to_tile_10_24_3),
		.in_wire_3_0(vertical_tile_10_24_to_tile_11_24_0),
		.in_wire_3_1(vertical_tile_10_24_to_tile_11_24_1),
		.in_wire_3_2(vertical_tile_10_24_to_tile_11_24_2),
		.in_wire_3_3(vertical_tile_10_24_to_tile_11_24_3),
		.out_wire_1_0(vertical_tile_11_24_to_tile_12_24_0),
		.out_wire_1_1(vertical_tile_11_24_to_tile_12_24_1),
		.out_wire_1_2(vertical_tile_11_24_to_tile_12_24_2),
		.out_wire_1_3(vertical_tile_11_24_to_tile_12_24_3),
		.in_wire_1_0(vertical_tile_12_24_to_tile_11_24_0),
		.in_wire_1_1(vertical_tile_12_24_to_tile_11_24_1),
		.in_wire_1_2(vertical_tile_12_24_to_tile_11_24_2),
		.in_wire_1_3(vertical_tile_12_24_to_tile_11_24_3),
		.out_wire_2_0(horizontal_tile_11_24_to_tile_11_23_0),
		.out_wire_2_1(horizontal_tile_11_24_to_tile_11_23_1),
		.out_wire_2_2(horizontal_tile_11_24_to_tile_11_23_2),
		.out_wire_2_3(horizontal_tile_11_24_to_tile_11_23_3),
		.in_wire_2_0(horizontal_tile_11_23_to_tile_11_24_0),
		.in_wire_2_1(horizontal_tile_11_23_to_tile_11_24_1),
		.in_wire_2_2(horizontal_tile_11_23_to_tile_11_24_2),
		.in_wire_2_3(horizontal_tile_11_23_to_tile_11_24_3),
		.out_wire_0_0(horizontal_tile_11_24_to_tile_11_25_0),
		.out_wire_0_1(horizontal_tile_11_24_to_tile_11_25_1),
		.out_wire_0_2(horizontal_tile_11_24_to_tile_11_25_2),
		.out_wire_0_3(horizontal_tile_11_24_to_tile_11_25_3),
		.in_wire_0_0(horizontal_tile_11_25_to_tile_11_24_0),
		.in_wire_0_1(horizontal_tile_11_25_to_tile_11_24_1),
		.in_wire_0_2(horizontal_tile_11_25_to_tile_11_24_2),
		.in_wire_0_3(horizontal_tile_11_25_to_tile_11_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(377)
	);

	pe_tile pe_tile_11_25(
		.out_wire_3_0(vertical_tile_11_25_to_tile_10_25_0),
		.out_wire_3_1(vertical_tile_11_25_to_tile_10_25_1),
		.out_wire_3_2(vertical_tile_11_25_to_tile_10_25_2),
		.out_wire_3_3(vertical_tile_11_25_to_tile_10_25_3),
		.in_wire_3_0(vertical_tile_10_25_to_tile_11_25_0),
		.in_wire_3_1(vertical_tile_10_25_to_tile_11_25_1),
		.in_wire_3_2(vertical_tile_10_25_to_tile_11_25_2),
		.in_wire_3_3(vertical_tile_10_25_to_tile_11_25_3),
		.out_wire_1_0(vertical_tile_11_25_to_tile_12_25_0),
		.out_wire_1_1(vertical_tile_11_25_to_tile_12_25_1),
		.out_wire_1_2(vertical_tile_11_25_to_tile_12_25_2),
		.out_wire_1_3(vertical_tile_11_25_to_tile_12_25_3),
		.in_wire_1_0(vertical_tile_12_25_to_tile_11_25_0),
		.in_wire_1_1(vertical_tile_12_25_to_tile_11_25_1),
		.in_wire_1_2(vertical_tile_12_25_to_tile_11_25_2),
		.in_wire_1_3(vertical_tile_12_25_to_tile_11_25_3),
		.out_wire_2_0(horizontal_tile_11_25_to_tile_11_24_0),
		.out_wire_2_1(horizontal_tile_11_25_to_tile_11_24_1),
		.out_wire_2_2(horizontal_tile_11_25_to_tile_11_24_2),
		.out_wire_2_3(horizontal_tile_11_25_to_tile_11_24_3),
		.in_wire_2_0(horizontal_tile_11_24_to_tile_11_25_0),
		.in_wire_2_1(horizontal_tile_11_24_to_tile_11_25_1),
		.in_wire_2_2(horizontal_tile_11_24_to_tile_11_25_2),
		.in_wire_2_3(horizontal_tile_11_24_to_tile_11_25_3),
		.out_wire_0_0(horizontal_tile_11_25_to_tile_11_26_0),
		.out_wire_0_1(horizontal_tile_11_25_to_tile_11_26_1),
		.out_wire_0_2(horizontal_tile_11_25_to_tile_11_26_2),
		.out_wire_0_3(horizontal_tile_11_25_to_tile_11_26_3),
		.in_wire_0_0(horizontal_tile_11_26_to_tile_11_25_0),
		.in_wire_0_1(horizontal_tile_11_26_to_tile_11_25_1),
		.in_wire_0_2(horizontal_tile_11_26_to_tile_11_25_2),
		.in_wire_0_3(horizontal_tile_11_26_to_tile_11_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(378)
	);

	pe_tile pe_tile_11_26(
		.out_wire_3_0(vertical_tile_11_26_to_tile_10_26_0),
		.out_wire_3_1(vertical_tile_11_26_to_tile_10_26_1),
		.out_wire_3_2(vertical_tile_11_26_to_tile_10_26_2),
		.out_wire_3_3(vertical_tile_11_26_to_tile_10_26_3),
		.in_wire_3_0(vertical_tile_10_26_to_tile_11_26_0),
		.in_wire_3_1(vertical_tile_10_26_to_tile_11_26_1),
		.in_wire_3_2(vertical_tile_10_26_to_tile_11_26_2),
		.in_wire_3_3(vertical_tile_10_26_to_tile_11_26_3),
		.out_wire_1_0(vertical_tile_11_26_to_tile_12_26_0),
		.out_wire_1_1(vertical_tile_11_26_to_tile_12_26_1),
		.out_wire_1_2(vertical_tile_11_26_to_tile_12_26_2),
		.out_wire_1_3(vertical_tile_11_26_to_tile_12_26_3),
		.in_wire_1_0(vertical_tile_12_26_to_tile_11_26_0),
		.in_wire_1_1(vertical_tile_12_26_to_tile_11_26_1),
		.in_wire_1_2(vertical_tile_12_26_to_tile_11_26_2),
		.in_wire_1_3(vertical_tile_12_26_to_tile_11_26_3),
		.out_wire_2_0(horizontal_tile_11_26_to_tile_11_25_0),
		.out_wire_2_1(horizontal_tile_11_26_to_tile_11_25_1),
		.out_wire_2_2(horizontal_tile_11_26_to_tile_11_25_2),
		.out_wire_2_3(horizontal_tile_11_26_to_tile_11_25_3),
		.in_wire_2_0(horizontal_tile_11_25_to_tile_11_26_0),
		.in_wire_2_1(horizontal_tile_11_25_to_tile_11_26_1),
		.in_wire_2_2(horizontal_tile_11_25_to_tile_11_26_2),
		.in_wire_2_3(horizontal_tile_11_25_to_tile_11_26_3),
		.out_wire_0_0(horizontal_tile_11_26_to_tile_11_27_0),
		.out_wire_0_1(horizontal_tile_11_26_to_tile_11_27_1),
		.out_wire_0_2(horizontal_tile_11_26_to_tile_11_27_2),
		.out_wire_0_3(horizontal_tile_11_26_to_tile_11_27_3),
		.in_wire_0_0(horizontal_tile_11_27_to_tile_11_26_0),
		.in_wire_0_1(horizontal_tile_11_27_to_tile_11_26_1),
		.in_wire_0_2(horizontal_tile_11_27_to_tile_11_26_2),
		.in_wire_0_3(horizontal_tile_11_27_to_tile_11_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(379)
	);

	pe_tile pe_tile_11_27(
		.out_wire_3_0(vertical_tile_11_27_to_tile_10_27_0),
		.out_wire_3_1(vertical_tile_11_27_to_tile_10_27_1),
		.out_wire_3_2(vertical_tile_11_27_to_tile_10_27_2),
		.out_wire_3_3(vertical_tile_11_27_to_tile_10_27_3),
		.in_wire_3_0(vertical_tile_10_27_to_tile_11_27_0),
		.in_wire_3_1(vertical_tile_10_27_to_tile_11_27_1),
		.in_wire_3_2(vertical_tile_10_27_to_tile_11_27_2),
		.in_wire_3_3(vertical_tile_10_27_to_tile_11_27_3),
		.out_wire_1_0(vertical_tile_11_27_to_tile_12_27_0),
		.out_wire_1_1(vertical_tile_11_27_to_tile_12_27_1),
		.out_wire_1_2(vertical_tile_11_27_to_tile_12_27_2),
		.out_wire_1_3(vertical_tile_11_27_to_tile_12_27_3),
		.in_wire_1_0(vertical_tile_12_27_to_tile_11_27_0),
		.in_wire_1_1(vertical_tile_12_27_to_tile_11_27_1),
		.in_wire_1_2(vertical_tile_12_27_to_tile_11_27_2),
		.in_wire_1_3(vertical_tile_12_27_to_tile_11_27_3),
		.out_wire_2_0(horizontal_tile_11_27_to_tile_11_26_0),
		.out_wire_2_1(horizontal_tile_11_27_to_tile_11_26_1),
		.out_wire_2_2(horizontal_tile_11_27_to_tile_11_26_2),
		.out_wire_2_3(horizontal_tile_11_27_to_tile_11_26_3),
		.in_wire_2_0(horizontal_tile_11_26_to_tile_11_27_0),
		.in_wire_2_1(horizontal_tile_11_26_to_tile_11_27_1),
		.in_wire_2_2(horizontal_tile_11_26_to_tile_11_27_2),
		.in_wire_2_3(horizontal_tile_11_26_to_tile_11_27_3),
		.out_wire_0_0(horizontal_tile_11_27_to_tile_11_28_0),
		.out_wire_0_1(horizontal_tile_11_27_to_tile_11_28_1),
		.out_wire_0_2(horizontal_tile_11_27_to_tile_11_28_2),
		.out_wire_0_3(horizontal_tile_11_27_to_tile_11_28_3),
		.in_wire_0_0(horizontal_tile_11_28_to_tile_11_27_0),
		.in_wire_0_1(horizontal_tile_11_28_to_tile_11_27_1),
		.in_wire_0_2(horizontal_tile_11_28_to_tile_11_27_2),
		.in_wire_0_3(horizontal_tile_11_28_to_tile_11_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(380)
	);

	pe_tile pe_tile_11_28(
		.out_wire_3_0(vertical_tile_11_28_to_tile_10_28_0),
		.out_wire_3_1(vertical_tile_11_28_to_tile_10_28_1),
		.out_wire_3_2(vertical_tile_11_28_to_tile_10_28_2),
		.out_wire_3_3(vertical_tile_11_28_to_tile_10_28_3),
		.in_wire_3_0(vertical_tile_10_28_to_tile_11_28_0),
		.in_wire_3_1(vertical_tile_10_28_to_tile_11_28_1),
		.in_wire_3_2(vertical_tile_10_28_to_tile_11_28_2),
		.in_wire_3_3(vertical_tile_10_28_to_tile_11_28_3),
		.out_wire_1_0(vertical_tile_11_28_to_tile_12_28_0),
		.out_wire_1_1(vertical_tile_11_28_to_tile_12_28_1),
		.out_wire_1_2(vertical_tile_11_28_to_tile_12_28_2),
		.out_wire_1_3(vertical_tile_11_28_to_tile_12_28_3),
		.in_wire_1_0(vertical_tile_12_28_to_tile_11_28_0),
		.in_wire_1_1(vertical_tile_12_28_to_tile_11_28_1),
		.in_wire_1_2(vertical_tile_12_28_to_tile_11_28_2),
		.in_wire_1_3(vertical_tile_12_28_to_tile_11_28_3),
		.out_wire_2_0(horizontal_tile_11_28_to_tile_11_27_0),
		.out_wire_2_1(horizontal_tile_11_28_to_tile_11_27_1),
		.out_wire_2_2(horizontal_tile_11_28_to_tile_11_27_2),
		.out_wire_2_3(horizontal_tile_11_28_to_tile_11_27_3),
		.in_wire_2_0(horizontal_tile_11_27_to_tile_11_28_0),
		.in_wire_2_1(horizontal_tile_11_27_to_tile_11_28_1),
		.in_wire_2_2(horizontal_tile_11_27_to_tile_11_28_2),
		.in_wire_2_3(horizontal_tile_11_27_to_tile_11_28_3),
		.out_wire_0_0(horizontal_tile_11_28_to_tile_11_29_0),
		.out_wire_0_1(horizontal_tile_11_28_to_tile_11_29_1),
		.out_wire_0_2(horizontal_tile_11_28_to_tile_11_29_2),
		.out_wire_0_3(horizontal_tile_11_28_to_tile_11_29_3),
		.in_wire_0_0(horizontal_tile_11_29_to_tile_11_28_0),
		.in_wire_0_1(horizontal_tile_11_29_to_tile_11_28_1),
		.in_wire_0_2(horizontal_tile_11_29_to_tile_11_28_2),
		.in_wire_0_3(horizontal_tile_11_29_to_tile_11_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(381)
	);

	pe_tile pe_tile_11_29(
		.out_wire_3_0(vertical_tile_11_29_to_tile_10_29_0),
		.out_wire_3_1(vertical_tile_11_29_to_tile_10_29_1),
		.out_wire_3_2(vertical_tile_11_29_to_tile_10_29_2),
		.out_wire_3_3(vertical_tile_11_29_to_tile_10_29_3),
		.in_wire_3_0(vertical_tile_10_29_to_tile_11_29_0),
		.in_wire_3_1(vertical_tile_10_29_to_tile_11_29_1),
		.in_wire_3_2(vertical_tile_10_29_to_tile_11_29_2),
		.in_wire_3_3(vertical_tile_10_29_to_tile_11_29_3),
		.out_wire_1_0(vertical_tile_11_29_to_tile_12_29_0),
		.out_wire_1_1(vertical_tile_11_29_to_tile_12_29_1),
		.out_wire_1_2(vertical_tile_11_29_to_tile_12_29_2),
		.out_wire_1_3(vertical_tile_11_29_to_tile_12_29_3),
		.in_wire_1_0(vertical_tile_12_29_to_tile_11_29_0),
		.in_wire_1_1(vertical_tile_12_29_to_tile_11_29_1),
		.in_wire_1_2(vertical_tile_12_29_to_tile_11_29_2),
		.in_wire_1_3(vertical_tile_12_29_to_tile_11_29_3),
		.out_wire_2_0(horizontal_tile_11_29_to_tile_11_28_0),
		.out_wire_2_1(horizontal_tile_11_29_to_tile_11_28_1),
		.out_wire_2_2(horizontal_tile_11_29_to_tile_11_28_2),
		.out_wire_2_3(horizontal_tile_11_29_to_tile_11_28_3),
		.in_wire_2_0(horizontal_tile_11_28_to_tile_11_29_0),
		.in_wire_2_1(horizontal_tile_11_28_to_tile_11_29_1),
		.in_wire_2_2(horizontal_tile_11_28_to_tile_11_29_2),
		.in_wire_2_3(horizontal_tile_11_28_to_tile_11_29_3),
		.out_wire_0_0(horizontal_tile_11_29_to_tile_11_30_0),
		.out_wire_0_1(horizontal_tile_11_29_to_tile_11_30_1),
		.out_wire_0_2(horizontal_tile_11_29_to_tile_11_30_2),
		.out_wire_0_3(horizontal_tile_11_29_to_tile_11_30_3),
		.in_wire_0_0(horizontal_tile_11_30_to_tile_11_29_0),
		.in_wire_0_1(horizontal_tile_11_30_to_tile_11_29_1),
		.in_wire_0_2(horizontal_tile_11_30_to_tile_11_29_2),
		.in_wire_0_3(horizontal_tile_11_30_to_tile_11_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(382)
	);

	pe_tile pe_tile_11_30(
		.out_wire_3_0(vertical_tile_11_30_to_tile_10_30_0),
		.out_wire_3_1(vertical_tile_11_30_to_tile_10_30_1),
		.out_wire_3_2(vertical_tile_11_30_to_tile_10_30_2),
		.out_wire_3_3(vertical_tile_11_30_to_tile_10_30_3),
		.in_wire_3_0(vertical_tile_10_30_to_tile_11_30_0),
		.in_wire_3_1(vertical_tile_10_30_to_tile_11_30_1),
		.in_wire_3_2(vertical_tile_10_30_to_tile_11_30_2),
		.in_wire_3_3(vertical_tile_10_30_to_tile_11_30_3),
		.out_wire_1_0(vertical_tile_11_30_to_tile_12_30_0),
		.out_wire_1_1(vertical_tile_11_30_to_tile_12_30_1),
		.out_wire_1_2(vertical_tile_11_30_to_tile_12_30_2),
		.out_wire_1_3(vertical_tile_11_30_to_tile_12_30_3),
		.in_wire_1_0(vertical_tile_12_30_to_tile_11_30_0),
		.in_wire_1_1(vertical_tile_12_30_to_tile_11_30_1),
		.in_wire_1_2(vertical_tile_12_30_to_tile_11_30_2),
		.in_wire_1_3(vertical_tile_12_30_to_tile_11_30_3),
		.out_wire_2_0(horizontal_tile_11_30_to_tile_11_29_0),
		.out_wire_2_1(horizontal_tile_11_30_to_tile_11_29_1),
		.out_wire_2_2(horizontal_tile_11_30_to_tile_11_29_2),
		.out_wire_2_3(horizontal_tile_11_30_to_tile_11_29_3),
		.in_wire_2_0(horizontal_tile_11_29_to_tile_11_30_0),
		.in_wire_2_1(horizontal_tile_11_29_to_tile_11_30_1),
		.in_wire_2_2(horizontal_tile_11_29_to_tile_11_30_2),
		.in_wire_2_3(horizontal_tile_11_29_to_tile_11_30_3),
		.out_wire_0_0(horizontal_tile_11_30_to_tile_11_31_0),
		.out_wire_0_1(horizontal_tile_11_30_to_tile_11_31_1),
		.out_wire_0_2(horizontal_tile_11_30_to_tile_11_31_2),
		.out_wire_0_3(horizontal_tile_11_30_to_tile_11_31_3),
		.in_wire_0_0(horizontal_tile_11_31_to_tile_11_30_0),
		.in_wire_0_1(horizontal_tile_11_31_to_tile_11_30_1),
		.in_wire_0_2(horizontal_tile_11_31_to_tile_11_30_2),
		.in_wire_0_3(horizontal_tile_11_31_to_tile_11_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(383)
	);

	pe_tile_right pe_tile_11_31(
		.out_wire_3_0(vertical_tile_11_31_to_tile_10_31_0),
		.out_wire_3_1(vertical_tile_11_31_to_tile_10_31_1),
		.out_wire_3_2(vertical_tile_11_31_to_tile_10_31_2),
		.out_wire_3_3(vertical_tile_11_31_to_tile_10_31_3),
		.in_wire_3_0(vertical_tile_10_31_to_tile_11_31_0),
		.in_wire_3_1(vertical_tile_10_31_to_tile_11_31_1),
		.in_wire_3_2(vertical_tile_10_31_to_tile_11_31_2),
		.in_wire_3_3(vertical_tile_10_31_to_tile_11_31_3),
		.out_wire_1_0(vertical_tile_11_31_to_tile_12_31_0),
		.out_wire_1_1(vertical_tile_11_31_to_tile_12_31_1),
		.out_wire_1_2(vertical_tile_11_31_to_tile_12_31_2),
		.out_wire_1_3(vertical_tile_11_31_to_tile_12_31_3),
		.in_wire_1_0(vertical_tile_12_31_to_tile_11_31_0),
		.in_wire_1_1(vertical_tile_12_31_to_tile_11_31_1),
		.in_wire_1_2(vertical_tile_12_31_to_tile_11_31_2),
		.in_wire_1_3(vertical_tile_12_31_to_tile_11_31_3),
		.out_wire_2_0(horizontal_tile_11_31_to_tile_11_30_0),
		.out_wire_2_1(horizontal_tile_11_31_to_tile_11_30_1),
		.out_wire_2_2(horizontal_tile_11_31_to_tile_11_30_2),
		.out_wire_2_3(horizontal_tile_11_31_to_tile_11_30_3),
		.in_wire_2_0(horizontal_tile_11_30_to_tile_11_31_0),
		.in_wire_2_1(horizontal_tile_11_30_to_tile_11_31_1),
		.in_wire_2_2(horizontal_tile_11_30_to_tile_11_31_2),
		.in_wire_2_3(horizontal_tile_11_30_to_tile_11_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(384)
	);

	pe_tile_left pe_tile_12_0(
		.out_wire_3_0(vertical_tile_12_0_to_tile_11_0_0),
		.out_wire_3_1(vertical_tile_12_0_to_tile_11_0_1),
		.out_wire_3_2(vertical_tile_12_0_to_tile_11_0_2),
		.out_wire_3_3(vertical_tile_12_0_to_tile_11_0_3),
		.in_wire_3_0(vertical_tile_11_0_to_tile_12_0_0),
		.in_wire_3_1(vertical_tile_11_0_to_tile_12_0_1),
		.in_wire_3_2(vertical_tile_11_0_to_tile_12_0_2),
		.in_wire_3_3(vertical_tile_11_0_to_tile_12_0_3),
		.out_wire_1_0(vertical_tile_12_0_to_tile_13_0_0),
		.out_wire_1_1(vertical_tile_12_0_to_tile_13_0_1),
		.out_wire_1_2(vertical_tile_12_0_to_tile_13_0_2),
		.out_wire_1_3(vertical_tile_12_0_to_tile_13_0_3),
		.in_wire_1_0(vertical_tile_13_0_to_tile_12_0_0),
		.in_wire_1_1(vertical_tile_13_0_to_tile_12_0_1),
		.in_wire_1_2(vertical_tile_13_0_to_tile_12_0_2),
		.in_wire_1_3(vertical_tile_13_0_to_tile_12_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_12_0_to_tile_12_1_0),
		.out_wire_0_1(horizontal_tile_12_0_to_tile_12_1_1),
		.out_wire_0_2(horizontal_tile_12_0_to_tile_12_1_2),
		.out_wire_0_3(horizontal_tile_12_0_to_tile_12_1_3),
		.in_wire_0_0(horizontal_tile_12_1_to_tile_12_0_0),
		.in_wire_0_1(horizontal_tile_12_1_to_tile_12_0_1),
		.in_wire_0_2(horizontal_tile_12_1_to_tile_12_0_2),
		.in_wire_0_3(horizontal_tile_12_1_to_tile_12_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(385)
	);

	pe_tile pe_tile_12_1(
		.out_wire_3_0(vertical_tile_12_1_to_tile_11_1_0),
		.out_wire_3_1(vertical_tile_12_1_to_tile_11_1_1),
		.out_wire_3_2(vertical_tile_12_1_to_tile_11_1_2),
		.out_wire_3_3(vertical_tile_12_1_to_tile_11_1_3),
		.in_wire_3_0(vertical_tile_11_1_to_tile_12_1_0),
		.in_wire_3_1(vertical_tile_11_1_to_tile_12_1_1),
		.in_wire_3_2(vertical_tile_11_1_to_tile_12_1_2),
		.in_wire_3_3(vertical_tile_11_1_to_tile_12_1_3),
		.out_wire_1_0(vertical_tile_12_1_to_tile_13_1_0),
		.out_wire_1_1(vertical_tile_12_1_to_tile_13_1_1),
		.out_wire_1_2(vertical_tile_12_1_to_tile_13_1_2),
		.out_wire_1_3(vertical_tile_12_1_to_tile_13_1_3),
		.in_wire_1_0(vertical_tile_13_1_to_tile_12_1_0),
		.in_wire_1_1(vertical_tile_13_1_to_tile_12_1_1),
		.in_wire_1_2(vertical_tile_13_1_to_tile_12_1_2),
		.in_wire_1_3(vertical_tile_13_1_to_tile_12_1_3),
		.out_wire_2_0(horizontal_tile_12_1_to_tile_12_0_0),
		.out_wire_2_1(horizontal_tile_12_1_to_tile_12_0_1),
		.out_wire_2_2(horizontal_tile_12_1_to_tile_12_0_2),
		.out_wire_2_3(horizontal_tile_12_1_to_tile_12_0_3),
		.in_wire_2_0(horizontal_tile_12_0_to_tile_12_1_0),
		.in_wire_2_1(horizontal_tile_12_0_to_tile_12_1_1),
		.in_wire_2_2(horizontal_tile_12_0_to_tile_12_1_2),
		.in_wire_2_3(horizontal_tile_12_0_to_tile_12_1_3),
		.out_wire_0_0(horizontal_tile_12_1_to_tile_12_2_0),
		.out_wire_0_1(horizontal_tile_12_1_to_tile_12_2_1),
		.out_wire_0_2(horizontal_tile_12_1_to_tile_12_2_2),
		.out_wire_0_3(horizontal_tile_12_1_to_tile_12_2_3),
		.in_wire_0_0(horizontal_tile_12_2_to_tile_12_1_0),
		.in_wire_0_1(horizontal_tile_12_2_to_tile_12_1_1),
		.in_wire_0_2(horizontal_tile_12_2_to_tile_12_1_2),
		.in_wire_0_3(horizontal_tile_12_2_to_tile_12_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(386)
	);

	pe_tile pe_tile_12_2(
		.out_wire_3_0(vertical_tile_12_2_to_tile_11_2_0),
		.out_wire_3_1(vertical_tile_12_2_to_tile_11_2_1),
		.out_wire_3_2(vertical_tile_12_2_to_tile_11_2_2),
		.out_wire_3_3(vertical_tile_12_2_to_tile_11_2_3),
		.in_wire_3_0(vertical_tile_11_2_to_tile_12_2_0),
		.in_wire_3_1(vertical_tile_11_2_to_tile_12_2_1),
		.in_wire_3_2(vertical_tile_11_2_to_tile_12_2_2),
		.in_wire_3_3(vertical_tile_11_2_to_tile_12_2_3),
		.out_wire_1_0(vertical_tile_12_2_to_tile_13_2_0),
		.out_wire_1_1(vertical_tile_12_2_to_tile_13_2_1),
		.out_wire_1_2(vertical_tile_12_2_to_tile_13_2_2),
		.out_wire_1_3(vertical_tile_12_2_to_tile_13_2_3),
		.in_wire_1_0(vertical_tile_13_2_to_tile_12_2_0),
		.in_wire_1_1(vertical_tile_13_2_to_tile_12_2_1),
		.in_wire_1_2(vertical_tile_13_2_to_tile_12_2_2),
		.in_wire_1_3(vertical_tile_13_2_to_tile_12_2_3),
		.out_wire_2_0(horizontal_tile_12_2_to_tile_12_1_0),
		.out_wire_2_1(horizontal_tile_12_2_to_tile_12_1_1),
		.out_wire_2_2(horizontal_tile_12_2_to_tile_12_1_2),
		.out_wire_2_3(horizontal_tile_12_2_to_tile_12_1_3),
		.in_wire_2_0(horizontal_tile_12_1_to_tile_12_2_0),
		.in_wire_2_1(horizontal_tile_12_1_to_tile_12_2_1),
		.in_wire_2_2(horizontal_tile_12_1_to_tile_12_2_2),
		.in_wire_2_3(horizontal_tile_12_1_to_tile_12_2_3),
		.out_wire_0_0(horizontal_tile_12_2_to_tile_12_3_0),
		.out_wire_0_1(horizontal_tile_12_2_to_tile_12_3_1),
		.out_wire_0_2(horizontal_tile_12_2_to_tile_12_3_2),
		.out_wire_0_3(horizontal_tile_12_2_to_tile_12_3_3),
		.in_wire_0_0(horizontal_tile_12_3_to_tile_12_2_0),
		.in_wire_0_1(horizontal_tile_12_3_to_tile_12_2_1),
		.in_wire_0_2(horizontal_tile_12_3_to_tile_12_2_2),
		.in_wire_0_3(horizontal_tile_12_3_to_tile_12_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(387)
	);

	pe_tile pe_tile_12_3(
		.out_wire_3_0(vertical_tile_12_3_to_tile_11_3_0),
		.out_wire_3_1(vertical_tile_12_3_to_tile_11_3_1),
		.out_wire_3_2(vertical_tile_12_3_to_tile_11_3_2),
		.out_wire_3_3(vertical_tile_12_3_to_tile_11_3_3),
		.in_wire_3_0(vertical_tile_11_3_to_tile_12_3_0),
		.in_wire_3_1(vertical_tile_11_3_to_tile_12_3_1),
		.in_wire_3_2(vertical_tile_11_3_to_tile_12_3_2),
		.in_wire_3_3(vertical_tile_11_3_to_tile_12_3_3),
		.out_wire_1_0(vertical_tile_12_3_to_tile_13_3_0),
		.out_wire_1_1(vertical_tile_12_3_to_tile_13_3_1),
		.out_wire_1_2(vertical_tile_12_3_to_tile_13_3_2),
		.out_wire_1_3(vertical_tile_12_3_to_tile_13_3_3),
		.in_wire_1_0(vertical_tile_13_3_to_tile_12_3_0),
		.in_wire_1_1(vertical_tile_13_3_to_tile_12_3_1),
		.in_wire_1_2(vertical_tile_13_3_to_tile_12_3_2),
		.in_wire_1_3(vertical_tile_13_3_to_tile_12_3_3),
		.out_wire_2_0(horizontal_tile_12_3_to_tile_12_2_0),
		.out_wire_2_1(horizontal_tile_12_3_to_tile_12_2_1),
		.out_wire_2_2(horizontal_tile_12_3_to_tile_12_2_2),
		.out_wire_2_3(horizontal_tile_12_3_to_tile_12_2_3),
		.in_wire_2_0(horizontal_tile_12_2_to_tile_12_3_0),
		.in_wire_2_1(horizontal_tile_12_2_to_tile_12_3_1),
		.in_wire_2_2(horizontal_tile_12_2_to_tile_12_3_2),
		.in_wire_2_3(horizontal_tile_12_2_to_tile_12_3_3),
		.out_wire_0_0(horizontal_tile_12_3_to_tile_12_4_0),
		.out_wire_0_1(horizontal_tile_12_3_to_tile_12_4_1),
		.out_wire_0_2(horizontal_tile_12_3_to_tile_12_4_2),
		.out_wire_0_3(horizontal_tile_12_3_to_tile_12_4_3),
		.in_wire_0_0(horizontal_tile_12_4_to_tile_12_3_0),
		.in_wire_0_1(horizontal_tile_12_4_to_tile_12_3_1),
		.in_wire_0_2(horizontal_tile_12_4_to_tile_12_3_2),
		.in_wire_0_3(horizontal_tile_12_4_to_tile_12_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(388)
	);

	pe_tile pe_tile_12_4(
		.out_wire_3_0(vertical_tile_12_4_to_tile_11_4_0),
		.out_wire_3_1(vertical_tile_12_4_to_tile_11_4_1),
		.out_wire_3_2(vertical_tile_12_4_to_tile_11_4_2),
		.out_wire_3_3(vertical_tile_12_4_to_tile_11_4_3),
		.in_wire_3_0(vertical_tile_11_4_to_tile_12_4_0),
		.in_wire_3_1(vertical_tile_11_4_to_tile_12_4_1),
		.in_wire_3_2(vertical_tile_11_4_to_tile_12_4_2),
		.in_wire_3_3(vertical_tile_11_4_to_tile_12_4_3),
		.out_wire_1_0(vertical_tile_12_4_to_tile_13_4_0),
		.out_wire_1_1(vertical_tile_12_4_to_tile_13_4_1),
		.out_wire_1_2(vertical_tile_12_4_to_tile_13_4_2),
		.out_wire_1_3(vertical_tile_12_4_to_tile_13_4_3),
		.in_wire_1_0(vertical_tile_13_4_to_tile_12_4_0),
		.in_wire_1_1(vertical_tile_13_4_to_tile_12_4_1),
		.in_wire_1_2(vertical_tile_13_4_to_tile_12_4_2),
		.in_wire_1_3(vertical_tile_13_4_to_tile_12_4_3),
		.out_wire_2_0(horizontal_tile_12_4_to_tile_12_3_0),
		.out_wire_2_1(horizontal_tile_12_4_to_tile_12_3_1),
		.out_wire_2_2(horizontal_tile_12_4_to_tile_12_3_2),
		.out_wire_2_3(horizontal_tile_12_4_to_tile_12_3_3),
		.in_wire_2_0(horizontal_tile_12_3_to_tile_12_4_0),
		.in_wire_2_1(horizontal_tile_12_3_to_tile_12_4_1),
		.in_wire_2_2(horizontal_tile_12_3_to_tile_12_4_2),
		.in_wire_2_3(horizontal_tile_12_3_to_tile_12_4_3),
		.out_wire_0_0(horizontal_tile_12_4_to_tile_12_5_0),
		.out_wire_0_1(horizontal_tile_12_4_to_tile_12_5_1),
		.out_wire_0_2(horizontal_tile_12_4_to_tile_12_5_2),
		.out_wire_0_3(horizontal_tile_12_4_to_tile_12_5_3),
		.in_wire_0_0(horizontal_tile_12_5_to_tile_12_4_0),
		.in_wire_0_1(horizontal_tile_12_5_to_tile_12_4_1),
		.in_wire_0_2(horizontal_tile_12_5_to_tile_12_4_2),
		.in_wire_0_3(horizontal_tile_12_5_to_tile_12_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(389)
	);

	pe_tile pe_tile_12_5(
		.out_wire_3_0(vertical_tile_12_5_to_tile_11_5_0),
		.out_wire_3_1(vertical_tile_12_5_to_tile_11_5_1),
		.out_wire_3_2(vertical_tile_12_5_to_tile_11_5_2),
		.out_wire_3_3(vertical_tile_12_5_to_tile_11_5_3),
		.in_wire_3_0(vertical_tile_11_5_to_tile_12_5_0),
		.in_wire_3_1(vertical_tile_11_5_to_tile_12_5_1),
		.in_wire_3_2(vertical_tile_11_5_to_tile_12_5_2),
		.in_wire_3_3(vertical_tile_11_5_to_tile_12_5_3),
		.out_wire_1_0(vertical_tile_12_5_to_tile_13_5_0),
		.out_wire_1_1(vertical_tile_12_5_to_tile_13_5_1),
		.out_wire_1_2(vertical_tile_12_5_to_tile_13_5_2),
		.out_wire_1_3(vertical_tile_12_5_to_tile_13_5_3),
		.in_wire_1_0(vertical_tile_13_5_to_tile_12_5_0),
		.in_wire_1_1(vertical_tile_13_5_to_tile_12_5_1),
		.in_wire_1_2(vertical_tile_13_5_to_tile_12_5_2),
		.in_wire_1_3(vertical_tile_13_5_to_tile_12_5_3),
		.out_wire_2_0(horizontal_tile_12_5_to_tile_12_4_0),
		.out_wire_2_1(horizontal_tile_12_5_to_tile_12_4_1),
		.out_wire_2_2(horizontal_tile_12_5_to_tile_12_4_2),
		.out_wire_2_3(horizontal_tile_12_5_to_tile_12_4_3),
		.in_wire_2_0(horizontal_tile_12_4_to_tile_12_5_0),
		.in_wire_2_1(horizontal_tile_12_4_to_tile_12_5_1),
		.in_wire_2_2(horizontal_tile_12_4_to_tile_12_5_2),
		.in_wire_2_3(horizontal_tile_12_4_to_tile_12_5_3),
		.out_wire_0_0(horizontal_tile_12_5_to_tile_12_6_0),
		.out_wire_0_1(horizontal_tile_12_5_to_tile_12_6_1),
		.out_wire_0_2(horizontal_tile_12_5_to_tile_12_6_2),
		.out_wire_0_3(horizontal_tile_12_5_to_tile_12_6_3),
		.in_wire_0_0(horizontal_tile_12_6_to_tile_12_5_0),
		.in_wire_0_1(horizontal_tile_12_6_to_tile_12_5_1),
		.in_wire_0_2(horizontal_tile_12_6_to_tile_12_5_2),
		.in_wire_0_3(horizontal_tile_12_6_to_tile_12_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(390)
	);

	pe_tile pe_tile_12_6(
		.out_wire_3_0(vertical_tile_12_6_to_tile_11_6_0),
		.out_wire_3_1(vertical_tile_12_6_to_tile_11_6_1),
		.out_wire_3_2(vertical_tile_12_6_to_tile_11_6_2),
		.out_wire_3_3(vertical_tile_12_6_to_tile_11_6_3),
		.in_wire_3_0(vertical_tile_11_6_to_tile_12_6_0),
		.in_wire_3_1(vertical_tile_11_6_to_tile_12_6_1),
		.in_wire_3_2(vertical_tile_11_6_to_tile_12_6_2),
		.in_wire_3_3(vertical_tile_11_6_to_tile_12_6_3),
		.out_wire_1_0(vertical_tile_12_6_to_tile_13_6_0),
		.out_wire_1_1(vertical_tile_12_6_to_tile_13_6_1),
		.out_wire_1_2(vertical_tile_12_6_to_tile_13_6_2),
		.out_wire_1_3(vertical_tile_12_6_to_tile_13_6_3),
		.in_wire_1_0(vertical_tile_13_6_to_tile_12_6_0),
		.in_wire_1_1(vertical_tile_13_6_to_tile_12_6_1),
		.in_wire_1_2(vertical_tile_13_6_to_tile_12_6_2),
		.in_wire_1_3(vertical_tile_13_6_to_tile_12_6_3),
		.out_wire_2_0(horizontal_tile_12_6_to_tile_12_5_0),
		.out_wire_2_1(horizontal_tile_12_6_to_tile_12_5_1),
		.out_wire_2_2(horizontal_tile_12_6_to_tile_12_5_2),
		.out_wire_2_3(horizontal_tile_12_6_to_tile_12_5_3),
		.in_wire_2_0(horizontal_tile_12_5_to_tile_12_6_0),
		.in_wire_2_1(horizontal_tile_12_5_to_tile_12_6_1),
		.in_wire_2_2(horizontal_tile_12_5_to_tile_12_6_2),
		.in_wire_2_3(horizontal_tile_12_5_to_tile_12_6_3),
		.out_wire_0_0(horizontal_tile_12_6_to_tile_12_7_0),
		.out_wire_0_1(horizontal_tile_12_6_to_tile_12_7_1),
		.out_wire_0_2(horizontal_tile_12_6_to_tile_12_7_2),
		.out_wire_0_3(horizontal_tile_12_6_to_tile_12_7_3),
		.in_wire_0_0(horizontal_tile_12_7_to_tile_12_6_0),
		.in_wire_0_1(horizontal_tile_12_7_to_tile_12_6_1),
		.in_wire_0_2(horizontal_tile_12_7_to_tile_12_6_2),
		.in_wire_0_3(horizontal_tile_12_7_to_tile_12_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(391)
	);

	pe_tile pe_tile_12_7(
		.out_wire_3_0(vertical_tile_12_7_to_tile_11_7_0),
		.out_wire_3_1(vertical_tile_12_7_to_tile_11_7_1),
		.out_wire_3_2(vertical_tile_12_7_to_tile_11_7_2),
		.out_wire_3_3(vertical_tile_12_7_to_tile_11_7_3),
		.in_wire_3_0(vertical_tile_11_7_to_tile_12_7_0),
		.in_wire_3_1(vertical_tile_11_7_to_tile_12_7_1),
		.in_wire_3_2(vertical_tile_11_7_to_tile_12_7_2),
		.in_wire_3_3(vertical_tile_11_7_to_tile_12_7_3),
		.out_wire_1_0(vertical_tile_12_7_to_tile_13_7_0),
		.out_wire_1_1(vertical_tile_12_7_to_tile_13_7_1),
		.out_wire_1_2(vertical_tile_12_7_to_tile_13_7_2),
		.out_wire_1_3(vertical_tile_12_7_to_tile_13_7_3),
		.in_wire_1_0(vertical_tile_13_7_to_tile_12_7_0),
		.in_wire_1_1(vertical_tile_13_7_to_tile_12_7_1),
		.in_wire_1_2(vertical_tile_13_7_to_tile_12_7_2),
		.in_wire_1_3(vertical_tile_13_7_to_tile_12_7_3),
		.out_wire_2_0(horizontal_tile_12_7_to_tile_12_6_0),
		.out_wire_2_1(horizontal_tile_12_7_to_tile_12_6_1),
		.out_wire_2_2(horizontal_tile_12_7_to_tile_12_6_2),
		.out_wire_2_3(horizontal_tile_12_7_to_tile_12_6_3),
		.in_wire_2_0(horizontal_tile_12_6_to_tile_12_7_0),
		.in_wire_2_1(horizontal_tile_12_6_to_tile_12_7_1),
		.in_wire_2_2(horizontal_tile_12_6_to_tile_12_7_2),
		.in_wire_2_3(horizontal_tile_12_6_to_tile_12_7_3),
		.out_wire_0_0(horizontal_tile_12_7_to_tile_12_8_0),
		.out_wire_0_1(horizontal_tile_12_7_to_tile_12_8_1),
		.out_wire_0_2(horizontal_tile_12_7_to_tile_12_8_2),
		.out_wire_0_3(horizontal_tile_12_7_to_tile_12_8_3),
		.in_wire_0_0(horizontal_tile_12_8_to_tile_12_7_0),
		.in_wire_0_1(horizontal_tile_12_8_to_tile_12_7_1),
		.in_wire_0_2(horizontal_tile_12_8_to_tile_12_7_2),
		.in_wire_0_3(horizontal_tile_12_8_to_tile_12_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(392)
	);

	pe_tile pe_tile_12_8(
		.out_wire_3_0(vertical_tile_12_8_to_tile_11_8_0),
		.out_wire_3_1(vertical_tile_12_8_to_tile_11_8_1),
		.out_wire_3_2(vertical_tile_12_8_to_tile_11_8_2),
		.out_wire_3_3(vertical_tile_12_8_to_tile_11_8_3),
		.in_wire_3_0(vertical_tile_11_8_to_tile_12_8_0),
		.in_wire_3_1(vertical_tile_11_8_to_tile_12_8_1),
		.in_wire_3_2(vertical_tile_11_8_to_tile_12_8_2),
		.in_wire_3_3(vertical_tile_11_8_to_tile_12_8_3),
		.out_wire_1_0(vertical_tile_12_8_to_tile_13_8_0),
		.out_wire_1_1(vertical_tile_12_8_to_tile_13_8_1),
		.out_wire_1_2(vertical_tile_12_8_to_tile_13_8_2),
		.out_wire_1_3(vertical_tile_12_8_to_tile_13_8_3),
		.in_wire_1_0(vertical_tile_13_8_to_tile_12_8_0),
		.in_wire_1_1(vertical_tile_13_8_to_tile_12_8_1),
		.in_wire_1_2(vertical_tile_13_8_to_tile_12_8_2),
		.in_wire_1_3(vertical_tile_13_8_to_tile_12_8_3),
		.out_wire_2_0(horizontal_tile_12_8_to_tile_12_7_0),
		.out_wire_2_1(horizontal_tile_12_8_to_tile_12_7_1),
		.out_wire_2_2(horizontal_tile_12_8_to_tile_12_7_2),
		.out_wire_2_3(horizontal_tile_12_8_to_tile_12_7_3),
		.in_wire_2_0(horizontal_tile_12_7_to_tile_12_8_0),
		.in_wire_2_1(horizontal_tile_12_7_to_tile_12_8_1),
		.in_wire_2_2(horizontal_tile_12_7_to_tile_12_8_2),
		.in_wire_2_3(horizontal_tile_12_7_to_tile_12_8_3),
		.out_wire_0_0(horizontal_tile_12_8_to_tile_12_9_0),
		.out_wire_0_1(horizontal_tile_12_8_to_tile_12_9_1),
		.out_wire_0_2(horizontal_tile_12_8_to_tile_12_9_2),
		.out_wire_0_3(horizontal_tile_12_8_to_tile_12_9_3),
		.in_wire_0_0(horizontal_tile_12_9_to_tile_12_8_0),
		.in_wire_0_1(horizontal_tile_12_9_to_tile_12_8_1),
		.in_wire_0_2(horizontal_tile_12_9_to_tile_12_8_2),
		.in_wire_0_3(horizontal_tile_12_9_to_tile_12_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(393)
	);

	pe_tile pe_tile_12_9(
		.out_wire_3_0(vertical_tile_12_9_to_tile_11_9_0),
		.out_wire_3_1(vertical_tile_12_9_to_tile_11_9_1),
		.out_wire_3_2(vertical_tile_12_9_to_tile_11_9_2),
		.out_wire_3_3(vertical_tile_12_9_to_tile_11_9_3),
		.in_wire_3_0(vertical_tile_11_9_to_tile_12_9_0),
		.in_wire_3_1(vertical_tile_11_9_to_tile_12_9_1),
		.in_wire_3_2(vertical_tile_11_9_to_tile_12_9_2),
		.in_wire_3_3(vertical_tile_11_9_to_tile_12_9_3),
		.out_wire_1_0(vertical_tile_12_9_to_tile_13_9_0),
		.out_wire_1_1(vertical_tile_12_9_to_tile_13_9_1),
		.out_wire_1_2(vertical_tile_12_9_to_tile_13_9_2),
		.out_wire_1_3(vertical_tile_12_9_to_tile_13_9_3),
		.in_wire_1_0(vertical_tile_13_9_to_tile_12_9_0),
		.in_wire_1_1(vertical_tile_13_9_to_tile_12_9_1),
		.in_wire_1_2(vertical_tile_13_9_to_tile_12_9_2),
		.in_wire_1_3(vertical_tile_13_9_to_tile_12_9_3),
		.out_wire_2_0(horizontal_tile_12_9_to_tile_12_8_0),
		.out_wire_2_1(horizontal_tile_12_9_to_tile_12_8_1),
		.out_wire_2_2(horizontal_tile_12_9_to_tile_12_8_2),
		.out_wire_2_3(horizontal_tile_12_9_to_tile_12_8_3),
		.in_wire_2_0(horizontal_tile_12_8_to_tile_12_9_0),
		.in_wire_2_1(horizontal_tile_12_8_to_tile_12_9_1),
		.in_wire_2_2(horizontal_tile_12_8_to_tile_12_9_2),
		.in_wire_2_3(horizontal_tile_12_8_to_tile_12_9_3),
		.out_wire_0_0(horizontal_tile_12_9_to_tile_12_10_0),
		.out_wire_0_1(horizontal_tile_12_9_to_tile_12_10_1),
		.out_wire_0_2(horizontal_tile_12_9_to_tile_12_10_2),
		.out_wire_0_3(horizontal_tile_12_9_to_tile_12_10_3),
		.in_wire_0_0(horizontal_tile_12_10_to_tile_12_9_0),
		.in_wire_0_1(horizontal_tile_12_10_to_tile_12_9_1),
		.in_wire_0_2(horizontal_tile_12_10_to_tile_12_9_2),
		.in_wire_0_3(horizontal_tile_12_10_to_tile_12_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(394)
	);

	pe_tile pe_tile_12_10(
		.out_wire_3_0(vertical_tile_12_10_to_tile_11_10_0),
		.out_wire_3_1(vertical_tile_12_10_to_tile_11_10_1),
		.out_wire_3_2(vertical_tile_12_10_to_tile_11_10_2),
		.out_wire_3_3(vertical_tile_12_10_to_tile_11_10_3),
		.in_wire_3_0(vertical_tile_11_10_to_tile_12_10_0),
		.in_wire_3_1(vertical_tile_11_10_to_tile_12_10_1),
		.in_wire_3_2(vertical_tile_11_10_to_tile_12_10_2),
		.in_wire_3_3(vertical_tile_11_10_to_tile_12_10_3),
		.out_wire_1_0(vertical_tile_12_10_to_tile_13_10_0),
		.out_wire_1_1(vertical_tile_12_10_to_tile_13_10_1),
		.out_wire_1_2(vertical_tile_12_10_to_tile_13_10_2),
		.out_wire_1_3(vertical_tile_12_10_to_tile_13_10_3),
		.in_wire_1_0(vertical_tile_13_10_to_tile_12_10_0),
		.in_wire_1_1(vertical_tile_13_10_to_tile_12_10_1),
		.in_wire_1_2(vertical_tile_13_10_to_tile_12_10_2),
		.in_wire_1_3(vertical_tile_13_10_to_tile_12_10_3),
		.out_wire_2_0(horizontal_tile_12_10_to_tile_12_9_0),
		.out_wire_2_1(horizontal_tile_12_10_to_tile_12_9_1),
		.out_wire_2_2(horizontal_tile_12_10_to_tile_12_9_2),
		.out_wire_2_3(horizontal_tile_12_10_to_tile_12_9_3),
		.in_wire_2_0(horizontal_tile_12_9_to_tile_12_10_0),
		.in_wire_2_1(horizontal_tile_12_9_to_tile_12_10_1),
		.in_wire_2_2(horizontal_tile_12_9_to_tile_12_10_2),
		.in_wire_2_3(horizontal_tile_12_9_to_tile_12_10_3),
		.out_wire_0_0(horizontal_tile_12_10_to_tile_12_11_0),
		.out_wire_0_1(horizontal_tile_12_10_to_tile_12_11_1),
		.out_wire_0_2(horizontal_tile_12_10_to_tile_12_11_2),
		.out_wire_0_3(horizontal_tile_12_10_to_tile_12_11_3),
		.in_wire_0_0(horizontal_tile_12_11_to_tile_12_10_0),
		.in_wire_0_1(horizontal_tile_12_11_to_tile_12_10_1),
		.in_wire_0_2(horizontal_tile_12_11_to_tile_12_10_2),
		.in_wire_0_3(horizontal_tile_12_11_to_tile_12_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(395)
	);

	pe_tile pe_tile_12_11(
		.out_wire_3_0(vertical_tile_12_11_to_tile_11_11_0),
		.out_wire_3_1(vertical_tile_12_11_to_tile_11_11_1),
		.out_wire_3_2(vertical_tile_12_11_to_tile_11_11_2),
		.out_wire_3_3(vertical_tile_12_11_to_tile_11_11_3),
		.in_wire_3_0(vertical_tile_11_11_to_tile_12_11_0),
		.in_wire_3_1(vertical_tile_11_11_to_tile_12_11_1),
		.in_wire_3_2(vertical_tile_11_11_to_tile_12_11_2),
		.in_wire_3_3(vertical_tile_11_11_to_tile_12_11_3),
		.out_wire_1_0(vertical_tile_12_11_to_tile_13_11_0),
		.out_wire_1_1(vertical_tile_12_11_to_tile_13_11_1),
		.out_wire_1_2(vertical_tile_12_11_to_tile_13_11_2),
		.out_wire_1_3(vertical_tile_12_11_to_tile_13_11_3),
		.in_wire_1_0(vertical_tile_13_11_to_tile_12_11_0),
		.in_wire_1_1(vertical_tile_13_11_to_tile_12_11_1),
		.in_wire_1_2(vertical_tile_13_11_to_tile_12_11_2),
		.in_wire_1_3(vertical_tile_13_11_to_tile_12_11_3),
		.out_wire_2_0(horizontal_tile_12_11_to_tile_12_10_0),
		.out_wire_2_1(horizontal_tile_12_11_to_tile_12_10_1),
		.out_wire_2_2(horizontal_tile_12_11_to_tile_12_10_2),
		.out_wire_2_3(horizontal_tile_12_11_to_tile_12_10_3),
		.in_wire_2_0(horizontal_tile_12_10_to_tile_12_11_0),
		.in_wire_2_1(horizontal_tile_12_10_to_tile_12_11_1),
		.in_wire_2_2(horizontal_tile_12_10_to_tile_12_11_2),
		.in_wire_2_3(horizontal_tile_12_10_to_tile_12_11_3),
		.out_wire_0_0(horizontal_tile_12_11_to_tile_12_12_0),
		.out_wire_0_1(horizontal_tile_12_11_to_tile_12_12_1),
		.out_wire_0_2(horizontal_tile_12_11_to_tile_12_12_2),
		.out_wire_0_3(horizontal_tile_12_11_to_tile_12_12_3),
		.in_wire_0_0(horizontal_tile_12_12_to_tile_12_11_0),
		.in_wire_0_1(horizontal_tile_12_12_to_tile_12_11_1),
		.in_wire_0_2(horizontal_tile_12_12_to_tile_12_11_2),
		.in_wire_0_3(horizontal_tile_12_12_to_tile_12_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(396)
	);

	pe_tile pe_tile_12_12(
		.out_wire_3_0(vertical_tile_12_12_to_tile_11_12_0),
		.out_wire_3_1(vertical_tile_12_12_to_tile_11_12_1),
		.out_wire_3_2(vertical_tile_12_12_to_tile_11_12_2),
		.out_wire_3_3(vertical_tile_12_12_to_tile_11_12_3),
		.in_wire_3_0(vertical_tile_11_12_to_tile_12_12_0),
		.in_wire_3_1(vertical_tile_11_12_to_tile_12_12_1),
		.in_wire_3_2(vertical_tile_11_12_to_tile_12_12_2),
		.in_wire_3_3(vertical_tile_11_12_to_tile_12_12_3),
		.out_wire_1_0(vertical_tile_12_12_to_tile_13_12_0),
		.out_wire_1_1(vertical_tile_12_12_to_tile_13_12_1),
		.out_wire_1_2(vertical_tile_12_12_to_tile_13_12_2),
		.out_wire_1_3(vertical_tile_12_12_to_tile_13_12_3),
		.in_wire_1_0(vertical_tile_13_12_to_tile_12_12_0),
		.in_wire_1_1(vertical_tile_13_12_to_tile_12_12_1),
		.in_wire_1_2(vertical_tile_13_12_to_tile_12_12_2),
		.in_wire_1_3(vertical_tile_13_12_to_tile_12_12_3),
		.out_wire_2_0(horizontal_tile_12_12_to_tile_12_11_0),
		.out_wire_2_1(horizontal_tile_12_12_to_tile_12_11_1),
		.out_wire_2_2(horizontal_tile_12_12_to_tile_12_11_2),
		.out_wire_2_3(horizontal_tile_12_12_to_tile_12_11_3),
		.in_wire_2_0(horizontal_tile_12_11_to_tile_12_12_0),
		.in_wire_2_1(horizontal_tile_12_11_to_tile_12_12_1),
		.in_wire_2_2(horizontal_tile_12_11_to_tile_12_12_2),
		.in_wire_2_3(horizontal_tile_12_11_to_tile_12_12_3),
		.out_wire_0_0(horizontal_tile_12_12_to_tile_12_13_0),
		.out_wire_0_1(horizontal_tile_12_12_to_tile_12_13_1),
		.out_wire_0_2(horizontal_tile_12_12_to_tile_12_13_2),
		.out_wire_0_3(horizontal_tile_12_12_to_tile_12_13_3),
		.in_wire_0_0(horizontal_tile_12_13_to_tile_12_12_0),
		.in_wire_0_1(horizontal_tile_12_13_to_tile_12_12_1),
		.in_wire_0_2(horizontal_tile_12_13_to_tile_12_12_2),
		.in_wire_0_3(horizontal_tile_12_13_to_tile_12_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(397)
	);

	pe_tile pe_tile_12_13(
		.out_wire_3_0(vertical_tile_12_13_to_tile_11_13_0),
		.out_wire_3_1(vertical_tile_12_13_to_tile_11_13_1),
		.out_wire_3_2(vertical_tile_12_13_to_tile_11_13_2),
		.out_wire_3_3(vertical_tile_12_13_to_tile_11_13_3),
		.in_wire_3_0(vertical_tile_11_13_to_tile_12_13_0),
		.in_wire_3_1(vertical_tile_11_13_to_tile_12_13_1),
		.in_wire_3_2(vertical_tile_11_13_to_tile_12_13_2),
		.in_wire_3_3(vertical_tile_11_13_to_tile_12_13_3),
		.out_wire_1_0(vertical_tile_12_13_to_tile_13_13_0),
		.out_wire_1_1(vertical_tile_12_13_to_tile_13_13_1),
		.out_wire_1_2(vertical_tile_12_13_to_tile_13_13_2),
		.out_wire_1_3(vertical_tile_12_13_to_tile_13_13_3),
		.in_wire_1_0(vertical_tile_13_13_to_tile_12_13_0),
		.in_wire_1_1(vertical_tile_13_13_to_tile_12_13_1),
		.in_wire_1_2(vertical_tile_13_13_to_tile_12_13_2),
		.in_wire_1_3(vertical_tile_13_13_to_tile_12_13_3),
		.out_wire_2_0(horizontal_tile_12_13_to_tile_12_12_0),
		.out_wire_2_1(horizontal_tile_12_13_to_tile_12_12_1),
		.out_wire_2_2(horizontal_tile_12_13_to_tile_12_12_2),
		.out_wire_2_3(horizontal_tile_12_13_to_tile_12_12_3),
		.in_wire_2_0(horizontal_tile_12_12_to_tile_12_13_0),
		.in_wire_2_1(horizontal_tile_12_12_to_tile_12_13_1),
		.in_wire_2_2(horizontal_tile_12_12_to_tile_12_13_2),
		.in_wire_2_3(horizontal_tile_12_12_to_tile_12_13_3),
		.out_wire_0_0(horizontal_tile_12_13_to_tile_12_14_0),
		.out_wire_0_1(horizontal_tile_12_13_to_tile_12_14_1),
		.out_wire_0_2(horizontal_tile_12_13_to_tile_12_14_2),
		.out_wire_0_3(horizontal_tile_12_13_to_tile_12_14_3),
		.in_wire_0_0(horizontal_tile_12_14_to_tile_12_13_0),
		.in_wire_0_1(horizontal_tile_12_14_to_tile_12_13_1),
		.in_wire_0_2(horizontal_tile_12_14_to_tile_12_13_2),
		.in_wire_0_3(horizontal_tile_12_14_to_tile_12_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(398)
	);

	pe_tile pe_tile_12_14(
		.out_wire_3_0(vertical_tile_12_14_to_tile_11_14_0),
		.out_wire_3_1(vertical_tile_12_14_to_tile_11_14_1),
		.out_wire_3_2(vertical_tile_12_14_to_tile_11_14_2),
		.out_wire_3_3(vertical_tile_12_14_to_tile_11_14_3),
		.in_wire_3_0(vertical_tile_11_14_to_tile_12_14_0),
		.in_wire_3_1(vertical_tile_11_14_to_tile_12_14_1),
		.in_wire_3_2(vertical_tile_11_14_to_tile_12_14_2),
		.in_wire_3_3(vertical_tile_11_14_to_tile_12_14_3),
		.out_wire_1_0(vertical_tile_12_14_to_tile_13_14_0),
		.out_wire_1_1(vertical_tile_12_14_to_tile_13_14_1),
		.out_wire_1_2(vertical_tile_12_14_to_tile_13_14_2),
		.out_wire_1_3(vertical_tile_12_14_to_tile_13_14_3),
		.in_wire_1_0(vertical_tile_13_14_to_tile_12_14_0),
		.in_wire_1_1(vertical_tile_13_14_to_tile_12_14_1),
		.in_wire_1_2(vertical_tile_13_14_to_tile_12_14_2),
		.in_wire_1_3(vertical_tile_13_14_to_tile_12_14_3),
		.out_wire_2_0(horizontal_tile_12_14_to_tile_12_13_0),
		.out_wire_2_1(horizontal_tile_12_14_to_tile_12_13_1),
		.out_wire_2_2(horizontal_tile_12_14_to_tile_12_13_2),
		.out_wire_2_3(horizontal_tile_12_14_to_tile_12_13_3),
		.in_wire_2_0(horizontal_tile_12_13_to_tile_12_14_0),
		.in_wire_2_1(horizontal_tile_12_13_to_tile_12_14_1),
		.in_wire_2_2(horizontal_tile_12_13_to_tile_12_14_2),
		.in_wire_2_3(horizontal_tile_12_13_to_tile_12_14_3),
		.out_wire_0_0(horizontal_tile_12_14_to_tile_12_15_0),
		.out_wire_0_1(horizontal_tile_12_14_to_tile_12_15_1),
		.out_wire_0_2(horizontal_tile_12_14_to_tile_12_15_2),
		.out_wire_0_3(horizontal_tile_12_14_to_tile_12_15_3),
		.in_wire_0_0(horizontal_tile_12_15_to_tile_12_14_0),
		.in_wire_0_1(horizontal_tile_12_15_to_tile_12_14_1),
		.in_wire_0_2(horizontal_tile_12_15_to_tile_12_14_2),
		.in_wire_0_3(horizontal_tile_12_15_to_tile_12_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(399)
	);

	pe_tile pe_tile_12_15(
		.out_wire_3_0(vertical_tile_12_15_to_tile_11_15_0),
		.out_wire_3_1(vertical_tile_12_15_to_tile_11_15_1),
		.out_wire_3_2(vertical_tile_12_15_to_tile_11_15_2),
		.out_wire_3_3(vertical_tile_12_15_to_tile_11_15_3),
		.in_wire_3_0(vertical_tile_11_15_to_tile_12_15_0),
		.in_wire_3_1(vertical_tile_11_15_to_tile_12_15_1),
		.in_wire_3_2(vertical_tile_11_15_to_tile_12_15_2),
		.in_wire_3_3(vertical_tile_11_15_to_tile_12_15_3),
		.out_wire_1_0(vertical_tile_12_15_to_tile_13_15_0),
		.out_wire_1_1(vertical_tile_12_15_to_tile_13_15_1),
		.out_wire_1_2(vertical_tile_12_15_to_tile_13_15_2),
		.out_wire_1_3(vertical_tile_12_15_to_tile_13_15_3),
		.in_wire_1_0(vertical_tile_13_15_to_tile_12_15_0),
		.in_wire_1_1(vertical_tile_13_15_to_tile_12_15_1),
		.in_wire_1_2(vertical_tile_13_15_to_tile_12_15_2),
		.in_wire_1_3(vertical_tile_13_15_to_tile_12_15_3),
		.out_wire_2_0(horizontal_tile_12_15_to_tile_12_14_0),
		.out_wire_2_1(horizontal_tile_12_15_to_tile_12_14_1),
		.out_wire_2_2(horizontal_tile_12_15_to_tile_12_14_2),
		.out_wire_2_3(horizontal_tile_12_15_to_tile_12_14_3),
		.in_wire_2_0(horizontal_tile_12_14_to_tile_12_15_0),
		.in_wire_2_1(horizontal_tile_12_14_to_tile_12_15_1),
		.in_wire_2_2(horizontal_tile_12_14_to_tile_12_15_2),
		.in_wire_2_3(horizontal_tile_12_14_to_tile_12_15_3),
		.out_wire_0_0(horizontal_tile_12_15_to_tile_12_16_0),
		.out_wire_0_1(horizontal_tile_12_15_to_tile_12_16_1),
		.out_wire_0_2(horizontal_tile_12_15_to_tile_12_16_2),
		.out_wire_0_3(horizontal_tile_12_15_to_tile_12_16_3),
		.in_wire_0_0(horizontal_tile_12_16_to_tile_12_15_0),
		.in_wire_0_1(horizontal_tile_12_16_to_tile_12_15_1),
		.in_wire_0_2(horizontal_tile_12_16_to_tile_12_15_2),
		.in_wire_0_3(horizontal_tile_12_16_to_tile_12_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(400)
	);

	pe_tile pe_tile_12_16(
		.out_wire_3_0(vertical_tile_12_16_to_tile_11_16_0),
		.out_wire_3_1(vertical_tile_12_16_to_tile_11_16_1),
		.out_wire_3_2(vertical_tile_12_16_to_tile_11_16_2),
		.out_wire_3_3(vertical_tile_12_16_to_tile_11_16_3),
		.in_wire_3_0(vertical_tile_11_16_to_tile_12_16_0),
		.in_wire_3_1(vertical_tile_11_16_to_tile_12_16_1),
		.in_wire_3_2(vertical_tile_11_16_to_tile_12_16_2),
		.in_wire_3_3(vertical_tile_11_16_to_tile_12_16_3),
		.out_wire_1_0(vertical_tile_12_16_to_tile_13_16_0),
		.out_wire_1_1(vertical_tile_12_16_to_tile_13_16_1),
		.out_wire_1_2(vertical_tile_12_16_to_tile_13_16_2),
		.out_wire_1_3(vertical_tile_12_16_to_tile_13_16_3),
		.in_wire_1_0(vertical_tile_13_16_to_tile_12_16_0),
		.in_wire_1_1(vertical_tile_13_16_to_tile_12_16_1),
		.in_wire_1_2(vertical_tile_13_16_to_tile_12_16_2),
		.in_wire_1_3(vertical_tile_13_16_to_tile_12_16_3),
		.out_wire_2_0(horizontal_tile_12_16_to_tile_12_15_0),
		.out_wire_2_1(horizontal_tile_12_16_to_tile_12_15_1),
		.out_wire_2_2(horizontal_tile_12_16_to_tile_12_15_2),
		.out_wire_2_3(horizontal_tile_12_16_to_tile_12_15_3),
		.in_wire_2_0(horizontal_tile_12_15_to_tile_12_16_0),
		.in_wire_2_1(horizontal_tile_12_15_to_tile_12_16_1),
		.in_wire_2_2(horizontal_tile_12_15_to_tile_12_16_2),
		.in_wire_2_3(horizontal_tile_12_15_to_tile_12_16_3),
		.out_wire_0_0(horizontal_tile_12_16_to_tile_12_17_0),
		.out_wire_0_1(horizontal_tile_12_16_to_tile_12_17_1),
		.out_wire_0_2(horizontal_tile_12_16_to_tile_12_17_2),
		.out_wire_0_3(horizontal_tile_12_16_to_tile_12_17_3),
		.in_wire_0_0(horizontal_tile_12_17_to_tile_12_16_0),
		.in_wire_0_1(horizontal_tile_12_17_to_tile_12_16_1),
		.in_wire_0_2(horizontal_tile_12_17_to_tile_12_16_2),
		.in_wire_0_3(horizontal_tile_12_17_to_tile_12_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(401)
	);

	pe_tile pe_tile_12_17(
		.out_wire_3_0(vertical_tile_12_17_to_tile_11_17_0),
		.out_wire_3_1(vertical_tile_12_17_to_tile_11_17_1),
		.out_wire_3_2(vertical_tile_12_17_to_tile_11_17_2),
		.out_wire_3_3(vertical_tile_12_17_to_tile_11_17_3),
		.in_wire_3_0(vertical_tile_11_17_to_tile_12_17_0),
		.in_wire_3_1(vertical_tile_11_17_to_tile_12_17_1),
		.in_wire_3_2(vertical_tile_11_17_to_tile_12_17_2),
		.in_wire_3_3(vertical_tile_11_17_to_tile_12_17_3),
		.out_wire_1_0(vertical_tile_12_17_to_tile_13_17_0),
		.out_wire_1_1(vertical_tile_12_17_to_tile_13_17_1),
		.out_wire_1_2(vertical_tile_12_17_to_tile_13_17_2),
		.out_wire_1_3(vertical_tile_12_17_to_tile_13_17_3),
		.in_wire_1_0(vertical_tile_13_17_to_tile_12_17_0),
		.in_wire_1_1(vertical_tile_13_17_to_tile_12_17_1),
		.in_wire_1_2(vertical_tile_13_17_to_tile_12_17_2),
		.in_wire_1_3(vertical_tile_13_17_to_tile_12_17_3),
		.out_wire_2_0(horizontal_tile_12_17_to_tile_12_16_0),
		.out_wire_2_1(horizontal_tile_12_17_to_tile_12_16_1),
		.out_wire_2_2(horizontal_tile_12_17_to_tile_12_16_2),
		.out_wire_2_3(horizontal_tile_12_17_to_tile_12_16_3),
		.in_wire_2_0(horizontal_tile_12_16_to_tile_12_17_0),
		.in_wire_2_1(horizontal_tile_12_16_to_tile_12_17_1),
		.in_wire_2_2(horizontal_tile_12_16_to_tile_12_17_2),
		.in_wire_2_3(horizontal_tile_12_16_to_tile_12_17_3),
		.out_wire_0_0(horizontal_tile_12_17_to_tile_12_18_0),
		.out_wire_0_1(horizontal_tile_12_17_to_tile_12_18_1),
		.out_wire_0_2(horizontal_tile_12_17_to_tile_12_18_2),
		.out_wire_0_3(horizontal_tile_12_17_to_tile_12_18_3),
		.in_wire_0_0(horizontal_tile_12_18_to_tile_12_17_0),
		.in_wire_0_1(horizontal_tile_12_18_to_tile_12_17_1),
		.in_wire_0_2(horizontal_tile_12_18_to_tile_12_17_2),
		.in_wire_0_3(horizontal_tile_12_18_to_tile_12_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(402)
	);

	pe_tile pe_tile_12_18(
		.out_wire_3_0(vertical_tile_12_18_to_tile_11_18_0),
		.out_wire_3_1(vertical_tile_12_18_to_tile_11_18_1),
		.out_wire_3_2(vertical_tile_12_18_to_tile_11_18_2),
		.out_wire_3_3(vertical_tile_12_18_to_tile_11_18_3),
		.in_wire_3_0(vertical_tile_11_18_to_tile_12_18_0),
		.in_wire_3_1(vertical_tile_11_18_to_tile_12_18_1),
		.in_wire_3_2(vertical_tile_11_18_to_tile_12_18_2),
		.in_wire_3_3(vertical_tile_11_18_to_tile_12_18_3),
		.out_wire_1_0(vertical_tile_12_18_to_tile_13_18_0),
		.out_wire_1_1(vertical_tile_12_18_to_tile_13_18_1),
		.out_wire_1_2(vertical_tile_12_18_to_tile_13_18_2),
		.out_wire_1_3(vertical_tile_12_18_to_tile_13_18_3),
		.in_wire_1_0(vertical_tile_13_18_to_tile_12_18_0),
		.in_wire_1_1(vertical_tile_13_18_to_tile_12_18_1),
		.in_wire_1_2(vertical_tile_13_18_to_tile_12_18_2),
		.in_wire_1_3(vertical_tile_13_18_to_tile_12_18_3),
		.out_wire_2_0(horizontal_tile_12_18_to_tile_12_17_0),
		.out_wire_2_1(horizontal_tile_12_18_to_tile_12_17_1),
		.out_wire_2_2(horizontal_tile_12_18_to_tile_12_17_2),
		.out_wire_2_3(horizontal_tile_12_18_to_tile_12_17_3),
		.in_wire_2_0(horizontal_tile_12_17_to_tile_12_18_0),
		.in_wire_2_1(horizontal_tile_12_17_to_tile_12_18_1),
		.in_wire_2_2(horizontal_tile_12_17_to_tile_12_18_2),
		.in_wire_2_3(horizontal_tile_12_17_to_tile_12_18_3),
		.out_wire_0_0(horizontal_tile_12_18_to_tile_12_19_0),
		.out_wire_0_1(horizontal_tile_12_18_to_tile_12_19_1),
		.out_wire_0_2(horizontal_tile_12_18_to_tile_12_19_2),
		.out_wire_0_3(horizontal_tile_12_18_to_tile_12_19_3),
		.in_wire_0_0(horizontal_tile_12_19_to_tile_12_18_0),
		.in_wire_0_1(horizontal_tile_12_19_to_tile_12_18_1),
		.in_wire_0_2(horizontal_tile_12_19_to_tile_12_18_2),
		.in_wire_0_3(horizontal_tile_12_19_to_tile_12_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(403)
	);

	pe_tile pe_tile_12_19(
		.out_wire_3_0(vertical_tile_12_19_to_tile_11_19_0),
		.out_wire_3_1(vertical_tile_12_19_to_tile_11_19_1),
		.out_wire_3_2(vertical_tile_12_19_to_tile_11_19_2),
		.out_wire_3_3(vertical_tile_12_19_to_tile_11_19_3),
		.in_wire_3_0(vertical_tile_11_19_to_tile_12_19_0),
		.in_wire_3_1(vertical_tile_11_19_to_tile_12_19_1),
		.in_wire_3_2(vertical_tile_11_19_to_tile_12_19_2),
		.in_wire_3_3(vertical_tile_11_19_to_tile_12_19_3),
		.out_wire_1_0(vertical_tile_12_19_to_tile_13_19_0),
		.out_wire_1_1(vertical_tile_12_19_to_tile_13_19_1),
		.out_wire_1_2(vertical_tile_12_19_to_tile_13_19_2),
		.out_wire_1_3(vertical_tile_12_19_to_tile_13_19_3),
		.in_wire_1_0(vertical_tile_13_19_to_tile_12_19_0),
		.in_wire_1_1(vertical_tile_13_19_to_tile_12_19_1),
		.in_wire_1_2(vertical_tile_13_19_to_tile_12_19_2),
		.in_wire_1_3(vertical_tile_13_19_to_tile_12_19_3),
		.out_wire_2_0(horizontal_tile_12_19_to_tile_12_18_0),
		.out_wire_2_1(horizontal_tile_12_19_to_tile_12_18_1),
		.out_wire_2_2(horizontal_tile_12_19_to_tile_12_18_2),
		.out_wire_2_3(horizontal_tile_12_19_to_tile_12_18_3),
		.in_wire_2_0(horizontal_tile_12_18_to_tile_12_19_0),
		.in_wire_2_1(horizontal_tile_12_18_to_tile_12_19_1),
		.in_wire_2_2(horizontal_tile_12_18_to_tile_12_19_2),
		.in_wire_2_3(horizontal_tile_12_18_to_tile_12_19_3),
		.out_wire_0_0(horizontal_tile_12_19_to_tile_12_20_0),
		.out_wire_0_1(horizontal_tile_12_19_to_tile_12_20_1),
		.out_wire_0_2(horizontal_tile_12_19_to_tile_12_20_2),
		.out_wire_0_3(horizontal_tile_12_19_to_tile_12_20_3),
		.in_wire_0_0(horizontal_tile_12_20_to_tile_12_19_0),
		.in_wire_0_1(horizontal_tile_12_20_to_tile_12_19_1),
		.in_wire_0_2(horizontal_tile_12_20_to_tile_12_19_2),
		.in_wire_0_3(horizontal_tile_12_20_to_tile_12_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(404)
	);

	pe_tile pe_tile_12_20(
		.out_wire_3_0(vertical_tile_12_20_to_tile_11_20_0),
		.out_wire_3_1(vertical_tile_12_20_to_tile_11_20_1),
		.out_wire_3_2(vertical_tile_12_20_to_tile_11_20_2),
		.out_wire_3_3(vertical_tile_12_20_to_tile_11_20_3),
		.in_wire_3_0(vertical_tile_11_20_to_tile_12_20_0),
		.in_wire_3_1(vertical_tile_11_20_to_tile_12_20_1),
		.in_wire_3_2(vertical_tile_11_20_to_tile_12_20_2),
		.in_wire_3_3(vertical_tile_11_20_to_tile_12_20_3),
		.out_wire_1_0(vertical_tile_12_20_to_tile_13_20_0),
		.out_wire_1_1(vertical_tile_12_20_to_tile_13_20_1),
		.out_wire_1_2(vertical_tile_12_20_to_tile_13_20_2),
		.out_wire_1_3(vertical_tile_12_20_to_tile_13_20_3),
		.in_wire_1_0(vertical_tile_13_20_to_tile_12_20_0),
		.in_wire_1_1(vertical_tile_13_20_to_tile_12_20_1),
		.in_wire_1_2(vertical_tile_13_20_to_tile_12_20_2),
		.in_wire_1_3(vertical_tile_13_20_to_tile_12_20_3),
		.out_wire_2_0(horizontal_tile_12_20_to_tile_12_19_0),
		.out_wire_2_1(horizontal_tile_12_20_to_tile_12_19_1),
		.out_wire_2_2(horizontal_tile_12_20_to_tile_12_19_2),
		.out_wire_2_3(horizontal_tile_12_20_to_tile_12_19_3),
		.in_wire_2_0(horizontal_tile_12_19_to_tile_12_20_0),
		.in_wire_2_1(horizontal_tile_12_19_to_tile_12_20_1),
		.in_wire_2_2(horizontal_tile_12_19_to_tile_12_20_2),
		.in_wire_2_3(horizontal_tile_12_19_to_tile_12_20_3),
		.out_wire_0_0(horizontal_tile_12_20_to_tile_12_21_0),
		.out_wire_0_1(horizontal_tile_12_20_to_tile_12_21_1),
		.out_wire_0_2(horizontal_tile_12_20_to_tile_12_21_2),
		.out_wire_0_3(horizontal_tile_12_20_to_tile_12_21_3),
		.in_wire_0_0(horizontal_tile_12_21_to_tile_12_20_0),
		.in_wire_0_1(horizontal_tile_12_21_to_tile_12_20_1),
		.in_wire_0_2(horizontal_tile_12_21_to_tile_12_20_2),
		.in_wire_0_3(horizontal_tile_12_21_to_tile_12_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(405)
	);

	pe_tile pe_tile_12_21(
		.out_wire_3_0(vertical_tile_12_21_to_tile_11_21_0),
		.out_wire_3_1(vertical_tile_12_21_to_tile_11_21_1),
		.out_wire_3_2(vertical_tile_12_21_to_tile_11_21_2),
		.out_wire_3_3(vertical_tile_12_21_to_tile_11_21_3),
		.in_wire_3_0(vertical_tile_11_21_to_tile_12_21_0),
		.in_wire_3_1(vertical_tile_11_21_to_tile_12_21_1),
		.in_wire_3_2(vertical_tile_11_21_to_tile_12_21_2),
		.in_wire_3_3(vertical_tile_11_21_to_tile_12_21_3),
		.out_wire_1_0(vertical_tile_12_21_to_tile_13_21_0),
		.out_wire_1_1(vertical_tile_12_21_to_tile_13_21_1),
		.out_wire_1_2(vertical_tile_12_21_to_tile_13_21_2),
		.out_wire_1_3(vertical_tile_12_21_to_tile_13_21_3),
		.in_wire_1_0(vertical_tile_13_21_to_tile_12_21_0),
		.in_wire_1_1(vertical_tile_13_21_to_tile_12_21_1),
		.in_wire_1_2(vertical_tile_13_21_to_tile_12_21_2),
		.in_wire_1_3(vertical_tile_13_21_to_tile_12_21_3),
		.out_wire_2_0(horizontal_tile_12_21_to_tile_12_20_0),
		.out_wire_2_1(horizontal_tile_12_21_to_tile_12_20_1),
		.out_wire_2_2(horizontal_tile_12_21_to_tile_12_20_2),
		.out_wire_2_3(horizontal_tile_12_21_to_tile_12_20_3),
		.in_wire_2_0(horizontal_tile_12_20_to_tile_12_21_0),
		.in_wire_2_1(horizontal_tile_12_20_to_tile_12_21_1),
		.in_wire_2_2(horizontal_tile_12_20_to_tile_12_21_2),
		.in_wire_2_3(horizontal_tile_12_20_to_tile_12_21_3),
		.out_wire_0_0(horizontal_tile_12_21_to_tile_12_22_0),
		.out_wire_0_1(horizontal_tile_12_21_to_tile_12_22_1),
		.out_wire_0_2(horizontal_tile_12_21_to_tile_12_22_2),
		.out_wire_0_3(horizontal_tile_12_21_to_tile_12_22_3),
		.in_wire_0_0(horizontal_tile_12_22_to_tile_12_21_0),
		.in_wire_0_1(horizontal_tile_12_22_to_tile_12_21_1),
		.in_wire_0_2(horizontal_tile_12_22_to_tile_12_21_2),
		.in_wire_0_3(horizontal_tile_12_22_to_tile_12_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(406)
	);

	pe_tile pe_tile_12_22(
		.out_wire_3_0(vertical_tile_12_22_to_tile_11_22_0),
		.out_wire_3_1(vertical_tile_12_22_to_tile_11_22_1),
		.out_wire_3_2(vertical_tile_12_22_to_tile_11_22_2),
		.out_wire_3_3(vertical_tile_12_22_to_tile_11_22_3),
		.in_wire_3_0(vertical_tile_11_22_to_tile_12_22_0),
		.in_wire_3_1(vertical_tile_11_22_to_tile_12_22_1),
		.in_wire_3_2(vertical_tile_11_22_to_tile_12_22_2),
		.in_wire_3_3(vertical_tile_11_22_to_tile_12_22_3),
		.out_wire_1_0(vertical_tile_12_22_to_tile_13_22_0),
		.out_wire_1_1(vertical_tile_12_22_to_tile_13_22_1),
		.out_wire_1_2(vertical_tile_12_22_to_tile_13_22_2),
		.out_wire_1_3(vertical_tile_12_22_to_tile_13_22_3),
		.in_wire_1_0(vertical_tile_13_22_to_tile_12_22_0),
		.in_wire_1_1(vertical_tile_13_22_to_tile_12_22_1),
		.in_wire_1_2(vertical_tile_13_22_to_tile_12_22_2),
		.in_wire_1_3(vertical_tile_13_22_to_tile_12_22_3),
		.out_wire_2_0(horizontal_tile_12_22_to_tile_12_21_0),
		.out_wire_2_1(horizontal_tile_12_22_to_tile_12_21_1),
		.out_wire_2_2(horizontal_tile_12_22_to_tile_12_21_2),
		.out_wire_2_3(horizontal_tile_12_22_to_tile_12_21_3),
		.in_wire_2_0(horizontal_tile_12_21_to_tile_12_22_0),
		.in_wire_2_1(horizontal_tile_12_21_to_tile_12_22_1),
		.in_wire_2_2(horizontal_tile_12_21_to_tile_12_22_2),
		.in_wire_2_3(horizontal_tile_12_21_to_tile_12_22_3),
		.out_wire_0_0(horizontal_tile_12_22_to_tile_12_23_0),
		.out_wire_0_1(horizontal_tile_12_22_to_tile_12_23_1),
		.out_wire_0_2(horizontal_tile_12_22_to_tile_12_23_2),
		.out_wire_0_3(horizontal_tile_12_22_to_tile_12_23_3),
		.in_wire_0_0(horizontal_tile_12_23_to_tile_12_22_0),
		.in_wire_0_1(horizontal_tile_12_23_to_tile_12_22_1),
		.in_wire_0_2(horizontal_tile_12_23_to_tile_12_22_2),
		.in_wire_0_3(horizontal_tile_12_23_to_tile_12_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(407)
	);

	pe_tile pe_tile_12_23(
		.out_wire_3_0(vertical_tile_12_23_to_tile_11_23_0),
		.out_wire_3_1(vertical_tile_12_23_to_tile_11_23_1),
		.out_wire_3_2(vertical_tile_12_23_to_tile_11_23_2),
		.out_wire_3_3(vertical_tile_12_23_to_tile_11_23_3),
		.in_wire_3_0(vertical_tile_11_23_to_tile_12_23_0),
		.in_wire_3_1(vertical_tile_11_23_to_tile_12_23_1),
		.in_wire_3_2(vertical_tile_11_23_to_tile_12_23_2),
		.in_wire_3_3(vertical_tile_11_23_to_tile_12_23_3),
		.out_wire_1_0(vertical_tile_12_23_to_tile_13_23_0),
		.out_wire_1_1(vertical_tile_12_23_to_tile_13_23_1),
		.out_wire_1_2(vertical_tile_12_23_to_tile_13_23_2),
		.out_wire_1_3(vertical_tile_12_23_to_tile_13_23_3),
		.in_wire_1_0(vertical_tile_13_23_to_tile_12_23_0),
		.in_wire_1_1(vertical_tile_13_23_to_tile_12_23_1),
		.in_wire_1_2(vertical_tile_13_23_to_tile_12_23_2),
		.in_wire_1_3(vertical_tile_13_23_to_tile_12_23_3),
		.out_wire_2_0(horizontal_tile_12_23_to_tile_12_22_0),
		.out_wire_2_1(horizontal_tile_12_23_to_tile_12_22_1),
		.out_wire_2_2(horizontal_tile_12_23_to_tile_12_22_2),
		.out_wire_2_3(horizontal_tile_12_23_to_tile_12_22_3),
		.in_wire_2_0(horizontal_tile_12_22_to_tile_12_23_0),
		.in_wire_2_1(horizontal_tile_12_22_to_tile_12_23_1),
		.in_wire_2_2(horizontal_tile_12_22_to_tile_12_23_2),
		.in_wire_2_3(horizontal_tile_12_22_to_tile_12_23_3),
		.out_wire_0_0(horizontal_tile_12_23_to_tile_12_24_0),
		.out_wire_0_1(horizontal_tile_12_23_to_tile_12_24_1),
		.out_wire_0_2(horizontal_tile_12_23_to_tile_12_24_2),
		.out_wire_0_3(horizontal_tile_12_23_to_tile_12_24_3),
		.in_wire_0_0(horizontal_tile_12_24_to_tile_12_23_0),
		.in_wire_0_1(horizontal_tile_12_24_to_tile_12_23_1),
		.in_wire_0_2(horizontal_tile_12_24_to_tile_12_23_2),
		.in_wire_0_3(horizontal_tile_12_24_to_tile_12_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(408)
	);

	pe_tile pe_tile_12_24(
		.out_wire_3_0(vertical_tile_12_24_to_tile_11_24_0),
		.out_wire_3_1(vertical_tile_12_24_to_tile_11_24_1),
		.out_wire_3_2(vertical_tile_12_24_to_tile_11_24_2),
		.out_wire_3_3(vertical_tile_12_24_to_tile_11_24_3),
		.in_wire_3_0(vertical_tile_11_24_to_tile_12_24_0),
		.in_wire_3_1(vertical_tile_11_24_to_tile_12_24_1),
		.in_wire_3_2(vertical_tile_11_24_to_tile_12_24_2),
		.in_wire_3_3(vertical_tile_11_24_to_tile_12_24_3),
		.out_wire_1_0(vertical_tile_12_24_to_tile_13_24_0),
		.out_wire_1_1(vertical_tile_12_24_to_tile_13_24_1),
		.out_wire_1_2(vertical_tile_12_24_to_tile_13_24_2),
		.out_wire_1_3(vertical_tile_12_24_to_tile_13_24_3),
		.in_wire_1_0(vertical_tile_13_24_to_tile_12_24_0),
		.in_wire_1_1(vertical_tile_13_24_to_tile_12_24_1),
		.in_wire_1_2(vertical_tile_13_24_to_tile_12_24_2),
		.in_wire_1_3(vertical_tile_13_24_to_tile_12_24_3),
		.out_wire_2_0(horizontal_tile_12_24_to_tile_12_23_0),
		.out_wire_2_1(horizontal_tile_12_24_to_tile_12_23_1),
		.out_wire_2_2(horizontal_tile_12_24_to_tile_12_23_2),
		.out_wire_2_3(horizontal_tile_12_24_to_tile_12_23_3),
		.in_wire_2_0(horizontal_tile_12_23_to_tile_12_24_0),
		.in_wire_2_1(horizontal_tile_12_23_to_tile_12_24_1),
		.in_wire_2_2(horizontal_tile_12_23_to_tile_12_24_2),
		.in_wire_2_3(horizontal_tile_12_23_to_tile_12_24_3),
		.out_wire_0_0(horizontal_tile_12_24_to_tile_12_25_0),
		.out_wire_0_1(horizontal_tile_12_24_to_tile_12_25_1),
		.out_wire_0_2(horizontal_tile_12_24_to_tile_12_25_2),
		.out_wire_0_3(horizontal_tile_12_24_to_tile_12_25_3),
		.in_wire_0_0(horizontal_tile_12_25_to_tile_12_24_0),
		.in_wire_0_1(horizontal_tile_12_25_to_tile_12_24_1),
		.in_wire_0_2(horizontal_tile_12_25_to_tile_12_24_2),
		.in_wire_0_3(horizontal_tile_12_25_to_tile_12_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(409)
	);

	pe_tile pe_tile_12_25(
		.out_wire_3_0(vertical_tile_12_25_to_tile_11_25_0),
		.out_wire_3_1(vertical_tile_12_25_to_tile_11_25_1),
		.out_wire_3_2(vertical_tile_12_25_to_tile_11_25_2),
		.out_wire_3_3(vertical_tile_12_25_to_tile_11_25_3),
		.in_wire_3_0(vertical_tile_11_25_to_tile_12_25_0),
		.in_wire_3_1(vertical_tile_11_25_to_tile_12_25_1),
		.in_wire_3_2(vertical_tile_11_25_to_tile_12_25_2),
		.in_wire_3_3(vertical_tile_11_25_to_tile_12_25_3),
		.out_wire_1_0(vertical_tile_12_25_to_tile_13_25_0),
		.out_wire_1_1(vertical_tile_12_25_to_tile_13_25_1),
		.out_wire_1_2(vertical_tile_12_25_to_tile_13_25_2),
		.out_wire_1_3(vertical_tile_12_25_to_tile_13_25_3),
		.in_wire_1_0(vertical_tile_13_25_to_tile_12_25_0),
		.in_wire_1_1(vertical_tile_13_25_to_tile_12_25_1),
		.in_wire_1_2(vertical_tile_13_25_to_tile_12_25_2),
		.in_wire_1_3(vertical_tile_13_25_to_tile_12_25_3),
		.out_wire_2_0(horizontal_tile_12_25_to_tile_12_24_0),
		.out_wire_2_1(horizontal_tile_12_25_to_tile_12_24_1),
		.out_wire_2_2(horizontal_tile_12_25_to_tile_12_24_2),
		.out_wire_2_3(horizontal_tile_12_25_to_tile_12_24_3),
		.in_wire_2_0(horizontal_tile_12_24_to_tile_12_25_0),
		.in_wire_2_1(horizontal_tile_12_24_to_tile_12_25_1),
		.in_wire_2_2(horizontal_tile_12_24_to_tile_12_25_2),
		.in_wire_2_3(horizontal_tile_12_24_to_tile_12_25_3),
		.out_wire_0_0(horizontal_tile_12_25_to_tile_12_26_0),
		.out_wire_0_1(horizontal_tile_12_25_to_tile_12_26_1),
		.out_wire_0_2(horizontal_tile_12_25_to_tile_12_26_2),
		.out_wire_0_3(horizontal_tile_12_25_to_tile_12_26_3),
		.in_wire_0_0(horizontal_tile_12_26_to_tile_12_25_0),
		.in_wire_0_1(horizontal_tile_12_26_to_tile_12_25_1),
		.in_wire_0_2(horizontal_tile_12_26_to_tile_12_25_2),
		.in_wire_0_3(horizontal_tile_12_26_to_tile_12_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(410)
	);

	pe_tile pe_tile_12_26(
		.out_wire_3_0(vertical_tile_12_26_to_tile_11_26_0),
		.out_wire_3_1(vertical_tile_12_26_to_tile_11_26_1),
		.out_wire_3_2(vertical_tile_12_26_to_tile_11_26_2),
		.out_wire_3_3(vertical_tile_12_26_to_tile_11_26_3),
		.in_wire_3_0(vertical_tile_11_26_to_tile_12_26_0),
		.in_wire_3_1(vertical_tile_11_26_to_tile_12_26_1),
		.in_wire_3_2(vertical_tile_11_26_to_tile_12_26_2),
		.in_wire_3_3(vertical_tile_11_26_to_tile_12_26_3),
		.out_wire_1_0(vertical_tile_12_26_to_tile_13_26_0),
		.out_wire_1_1(vertical_tile_12_26_to_tile_13_26_1),
		.out_wire_1_2(vertical_tile_12_26_to_tile_13_26_2),
		.out_wire_1_3(vertical_tile_12_26_to_tile_13_26_3),
		.in_wire_1_0(vertical_tile_13_26_to_tile_12_26_0),
		.in_wire_1_1(vertical_tile_13_26_to_tile_12_26_1),
		.in_wire_1_2(vertical_tile_13_26_to_tile_12_26_2),
		.in_wire_1_3(vertical_tile_13_26_to_tile_12_26_3),
		.out_wire_2_0(horizontal_tile_12_26_to_tile_12_25_0),
		.out_wire_2_1(horizontal_tile_12_26_to_tile_12_25_1),
		.out_wire_2_2(horizontal_tile_12_26_to_tile_12_25_2),
		.out_wire_2_3(horizontal_tile_12_26_to_tile_12_25_3),
		.in_wire_2_0(horizontal_tile_12_25_to_tile_12_26_0),
		.in_wire_2_1(horizontal_tile_12_25_to_tile_12_26_1),
		.in_wire_2_2(horizontal_tile_12_25_to_tile_12_26_2),
		.in_wire_2_3(horizontal_tile_12_25_to_tile_12_26_3),
		.out_wire_0_0(horizontal_tile_12_26_to_tile_12_27_0),
		.out_wire_0_1(horizontal_tile_12_26_to_tile_12_27_1),
		.out_wire_0_2(horizontal_tile_12_26_to_tile_12_27_2),
		.out_wire_0_3(horizontal_tile_12_26_to_tile_12_27_3),
		.in_wire_0_0(horizontal_tile_12_27_to_tile_12_26_0),
		.in_wire_0_1(horizontal_tile_12_27_to_tile_12_26_1),
		.in_wire_0_2(horizontal_tile_12_27_to_tile_12_26_2),
		.in_wire_0_3(horizontal_tile_12_27_to_tile_12_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(411)
	);

	pe_tile pe_tile_12_27(
		.out_wire_3_0(vertical_tile_12_27_to_tile_11_27_0),
		.out_wire_3_1(vertical_tile_12_27_to_tile_11_27_1),
		.out_wire_3_2(vertical_tile_12_27_to_tile_11_27_2),
		.out_wire_3_3(vertical_tile_12_27_to_tile_11_27_3),
		.in_wire_3_0(vertical_tile_11_27_to_tile_12_27_0),
		.in_wire_3_1(vertical_tile_11_27_to_tile_12_27_1),
		.in_wire_3_2(vertical_tile_11_27_to_tile_12_27_2),
		.in_wire_3_3(vertical_tile_11_27_to_tile_12_27_3),
		.out_wire_1_0(vertical_tile_12_27_to_tile_13_27_0),
		.out_wire_1_1(vertical_tile_12_27_to_tile_13_27_1),
		.out_wire_1_2(vertical_tile_12_27_to_tile_13_27_2),
		.out_wire_1_3(vertical_tile_12_27_to_tile_13_27_3),
		.in_wire_1_0(vertical_tile_13_27_to_tile_12_27_0),
		.in_wire_1_1(vertical_tile_13_27_to_tile_12_27_1),
		.in_wire_1_2(vertical_tile_13_27_to_tile_12_27_2),
		.in_wire_1_3(vertical_tile_13_27_to_tile_12_27_3),
		.out_wire_2_0(horizontal_tile_12_27_to_tile_12_26_0),
		.out_wire_2_1(horizontal_tile_12_27_to_tile_12_26_1),
		.out_wire_2_2(horizontal_tile_12_27_to_tile_12_26_2),
		.out_wire_2_3(horizontal_tile_12_27_to_tile_12_26_3),
		.in_wire_2_0(horizontal_tile_12_26_to_tile_12_27_0),
		.in_wire_2_1(horizontal_tile_12_26_to_tile_12_27_1),
		.in_wire_2_2(horizontal_tile_12_26_to_tile_12_27_2),
		.in_wire_2_3(horizontal_tile_12_26_to_tile_12_27_3),
		.out_wire_0_0(horizontal_tile_12_27_to_tile_12_28_0),
		.out_wire_0_1(horizontal_tile_12_27_to_tile_12_28_1),
		.out_wire_0_2(horizontal_tile_12_27_to_tile_12_28_2),
		.out_wire_0_3(horizontal_tile_12_27_to_tile_12_28_3),
		.in_wire_0_0(horizontal_tile_12_28_to_tile_12_27_0),
		.in_wire_0_1(horizontal_tile_12_28_to_tile_12_27_1),
		.in_wire_0_2(horizontal_tile_12_28_to_tile_12_27_2),
		.in_wire_0_3(horizontal_tile_12_28_to_tile_12_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(412)
	);

	pe_tile pe_tile_12_28(
		.out_wire_3_0(vertical_tile_12_28_to_tile_11_28_0),
		.out_wire_3_1(vertical_tile_12_28_to_tile_11_28_1),
		.out_wire_3_2(vertical_tile_12_28_to_tile_11_28_2),
		.out_wire_3_3(vertical_tile_12_28_to_tile_11_28_3),
		.in_wire_3_0(vertical_tile_11_28_to_tile_12_28_0),
		.in_wire_3_1(vertical_tile_11_28_to_tile_12_28_1),
		.in_wire_3_2(vertical_tile_11_28_to_tile_12_28_2),
		.in_wire_3_3(vertical_tile_11_28_to_tile_12_28_3),
		.out_wire_1_0(vertical_tile_12_28_to_tile_13_28_0),
		.out_wire_1_1(vertical_tile_12_28_to_tile_13_28_1),
		.out_wire_1_2(vertical_tile_12_28_to_tile_13_28_2),
		.out_wire_1_3(vertical_tile_12_28_to_tile_13_28_3),
		.in_wire_1_0(vertical_tile_13_28_to_tile_12_28_0),
		.in_wire_1_1(vertical_tile_13_28_to_tile_12_28_1),
		.in_wire_1_2(vertical_tile_13_28_to_tile_12_28_2),
		.in_wire_1_3(vertical_tile_13_28_to_tile_12_28_3),
		.out_wire_2_0(horizontal_tile_12_28_to_tile_12_27_0),
		.out_wire_2_1(horizontal_tile_12_28_to_tile_12_27_1),
		.out_wire_2_2(horizontal_tile_12_28_to_tile_12_27_2),
		.out_wire_2_3(horizontal_tile_12_28_to_tile_12_27_3),
		.in_wire_2_0(horizontal_tile_12_27_to_tile_12_28_0),
		.in_wire_2_1(horizontal_tile_12_27_to_tile_12_28_1),
		.in_wire_2_2(horizontal_tile_12_27_to_tile_12_28_2),
		.in_wire_2_3(horizontal_tile_12_27_to_tile_12_28_3),
		.out_wire_0_0(horizontal_tile_12_28_to_tile_12_29_0),
		.out_wire_0_1(horizontal_tile_12_28_to_tile_12_29_1),
		.out_wire_0_2(horizontal_tile_12_28_to_tile_12_29_2),
		.out_wire_0_3(horizontal_tile_12_28_to_tile_12_29_3),
		.in_wire_0_0(horizontal_tile_12_29_to_tile_12_28_0),
		.in_wire_0_1(horizontal_tile_12_29_to_tile_12_28_1),
		.in_wire_0_2(horizontal_tile_12_29_to_tile_12_28_2),
		.in_wire_0_3(horizontal_tile_12_29_to_tile_12_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(413)
	);

	pe_tile pe_tile_12_29(
		.out_wire_3_0(vertical_tile_12_29_to_tile_11_29_0),
		.out_wire_3_1(vertical_tile_12_29_to_tile_11_29_1),
		.out_wire_3_2(vertical_tile_12_29_to_tile_11_29_2),
		.out_wire_3_3(vertical_tile_12_29_to_tile_11_29_3),
		.in_wire_3_0(vertical_tile_11_29_to_tile_12_29_0),
		.in_wire_3_1(vertical_tile_11_29_to_tile_12_29_1),
		.in_wire_3_2(vertical_tile_11_29_to_tile_12_29_2),
		.in_wire_3_3(vertical_tile_11_29_to_tile_12_29_3),
		.out_wire_1_0(vertical_tile_12_29_to_tile_13_29_0),
		.out_wire_1_1(vertical_tile_12_29_to_tile_13_29_1),
		.out_wire_1_2(vertical_tile_12_29_to_tile_13_29_2),
		.out_wire_1_3(vertical_tile_12_29_to_tile_13_29_3),
		.in_wire_1_0(vertical_tile_13_29_to_tile_12_29_0),
		.in_wire_1_1(vertical_tile_13_29_to_tile_12_29_1),
		.in_wire_1_2(vertical_tile_13_29_to_tile_12_29_2),
		.in_wire_1_3(vertical_tile_13_29_to_tile_12_29_3),
		.out_wire_2_0(horizontal_tile_12_29_to_tile_12_28_0),
		.out_wire_2_1(horizontal_tile_12_29_to_tile_12_28_1),
		.out_wire_2_2(horizontal_tile_12_29_to_tile_12_28_2),
		.out_wire_2_3(horizontal_tile_12_29_to_tile_12_28_3),
		.in_wire_2_0(horizontal_tile_12_28_to_tile_12_29_0),
		.in_wire_2_1(horizontal_tile_12_28_to_tile_12_29_1),
		.in_wire_2_2(horizontal_tile_12_28_to_tile_12_29_2),
		.in_wire_2_3(horizontal_tile_12_28_to_tile_12_29_3),
		.out_wire_0_0(horizontal_tile_12_29_to_tile_12_30_0),
		.out_wire_0_1(horizontal_tile_12_29_to_tile_12_30_1),
		.out_wire_0_2(horizontal_tile_12_29_to_tile_12_30_2),
		.out_wire_0_3(horizontal_tile_12_29_to_tile_12_30_3),
		.in_wire_0_0(horizontal_tile_12_30_to_tile_12_29_0),
		.in_wire_0_1(horizontal_tile_12_30_to_tile_12_29_1),
		.in_wire_0_2(horizontal_tile_12_30_to_tile_12_29_2),
		.in_wire_0_3(horizontal_tile_12_30_to_tile_12_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(414)
	);

	pe_tile pe_tile_12_30(
		.out_wire_3_0(vertical_tile_12_30_to_tile_11_30_0),
		.out_wire_3_1(vertical_tile_12_30_to_tile_11_30_1),
		.out_wire_3_2(vertical_tile_12_30_to_tile_11_30_2),
		.out_wire_3_3(vertical_tile_12_30_to_tile_11_30_3),
		.in_wire_3_0(vertical_tile_11_30_to_tile_12_30_0),
		.in_wire_3_1(vertical_tile_11_30_to_tile_12_30_1),
		.in_wire_3_2(vertical_tile_11_30_to_tile_12_30_2),
		.in_wire_3_3(vertical_tile_11_30_to_tile_12_30_3),
		.out_wire_1_0(vertical_tile_12_30_to_tile_13_30_0),
		.out_wire_1_1(vertical_tile_12_30_to_tile_13_30_1),
		.out_wire_1_2(vertical_tile_12_30_to_tile_13_30_2),
		.out_wire_1_3(vertical_tile_12_30_to_tile_13_30_3),
		.in_wire_1_0(vertical_tile_13_30_to_tile_12_30_0),
		.in_wire_1_1(vertical_tile_13_30_to_tile_12_30_1),
		.in_wire_1_2(vertical_tile_13_30_to_tile_12_30_2),
		.in_wire_1_3(vertical_tile_13_30_to_tile_12_30_3),
		.out_wire_2_0(horizontal_tile_12_30_to_tile_12_29_0),
		.out_wire_2_1(horizontal_tile_12_30_to_tile_12_29_1),
		.out_wire_2_2(horizontal_tile_12_30_to_tile_12_29_2),
		.out_wire_2_3(horizontal_tile_12_30_to_tile_12_29_3),
		.in_wire_2_0(horizontal_tile_12_29_to_tile_12_30_0),
		.in_wire_2_1(horizontal_tile_12_29_to_tile_12_30_1),
		.in_wire_2_2(horizontal_tile_12_29_to_tile_12_30_2),
		.in_wire_2_3(horizontal_tile_12_29_to_tile_12_30_3),
		.out_wire_0_0(horizontal_tile_12_30_to_tile_12_31_0),
		.out_wire_0_1(horizontal_tile_12_30_to_tile_12_31_1),
		.out_wire_0_2(horizontal_tile_12_30_to_tile_12_31_2),
		.out_wire_0_3(horizontal_tile_12_30_to_tile_12_31_3),
		.in_wire_0_0(horizontal_tile_12_31_to_tile_12_30_0),
		.in_wire_0_1(horizontal_tile_12_31_to_tile_12_30_1),
		.in_wire_0_2(horizontal_tile_12_31_to_tile_12_30_2),
		.in_wire_0_3(horizontal_tile_12_31_to_tile_12_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(415)
	);

	pe_tile_right pe_tile_12_31(
		.out_wire_3_0(vertical_tile_12_31_to_tile_11_31_0),
		.out_wire_3_1(vertical_tile_12_31_to_tile_11_31_1),
		.out_wire_3_2(vertical_tile_12_31_to_tile_11_31_2),
		.out_wire_3_3(vertical_tile_12_31_to_tile_11_31_3),
		.in_wire_3_0(vertical_tile_11_31_to_tile_12_31_0),
		.in_wire_3_1(vertical_tile_11_31_to_tile_12_31_1),
		.in_wire_3_2(vertical_tile_11_31_to_tile_12_31_2),
		.in_wire_3_3(vertical_tile_11_31_to_tile_12_31_3),
		.out_wire_1_0(vertical_tile_12_31_to_tile_13_31_0),
		.out_wire_1_1(vertical_tile_12_31_to_tile_13_31_1),
		.out_wire_1_2(vertical_tile_12_31_to_tile_13_31_2),
		.out_wire_1_3(vertical_tile_12_31_to_tile_13_31_3),
		.in_wire_1_0(vertical_tile_13_31_to_tile_12_31_0),
		.in_wire_1_1(vertical_tile_13_31_to_tile_12_31_1),
		.in_wire_1_2(vertical_tile_13_31_to_tile_12_31_2),
		.in_wire_1_3(vertical_tile_13_31_to_tile_12_31_3),
		.out_wire_2_0(horizontal_tile_12_31_to_tile_12_30_0),
		.out_wire_2_1(horizontal_tile_12_31_to_tile_12_30_1),
		.out_wire_2_2(horizontal_tile_12_31_to_tile_12_30_2),
		.out_wire_2_3(horizontal_tile_12_31_to_tile_12_30_3),
		.in_wire_2_0(horizontal_tile_12_30_to_tile_12_31_0),
		.in_wire_2_1(horizontal_tile_12_30_to_tile_12_31_1),
		.in_wire_2_2(horizontal_tile_12_30_to_tile_12_31_2),
		.in_wire_2_3(horizontal_tile_12_30_to_tile_12_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(416)
	);

	pe_tile_left pe_tile_13_0(
		.out_wire_3_0(vertical_tile_13_0_to_tile_12_0_0),
		.out_wire_3_1(vertical_tile_13_0_to_tile_12_0_1),
		.out_wire_3_2(vertical_tile_13_0_to_tile_12_0_2),
		.out_wire_3_3(vertical_tile_13_0_to_tile_12_0_3),
		.in_wire_3_0(vertical_tile_12_0_to_tile_13_0_0),
		.in_wire_3_1(vertical_tile_12_0_to_tile_13_0_1),
		.in_wire_3_2(vertical_tile_12_0_to_tile_13_0_2),
		.in_wire_3_3(vertical_tile_12_0_to_tile_13_0_3),
		.out_wire_1_0(vertical_tile_13_0_to_tile_14_0_0),
		.out_wire_1_1(vertical_tile_13_0_to_tile_14_0_1),
		.out_wire_1_2(vertical_tile_13_0_to_tile_14_0_2),
		.out_wire_1_3(vertical_tile_13_0_to_tile_14_0_3),
		.in_wire_1_0(vertical_tile_14_0_to_tile_13_0_0),
		.in_wire_1_1(vertical_tile_14_0_to_tile_13_0_1),
		.in_wire_1_2(vertical_tile_14_0_to_tile_13_0_2),
		.in_wire_1_3(vertical_tile_14_0_to_tile_13_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_13_0_to_tile_13_1_0),
		.out_wire_0_1(horizontal_tile_13_0_to_tile_13_1_1),
		.out_wire_0_2(horizontal_tile_13_0_to_tile_13_1_2),
		.out_wire_0_3(horizontal_tile_13_0_to_tile_13_1_3),
		.in_wire_0_0(horizontal_tile_13_1_to_tile_13_0_0),
		.in_wire_0_1(horizontal_tile_13_1_to_tile_13_0_1),
		.in_wire_0_2(horizontal_tile_13_1_to_tile_13_0_2),
		.in_wire_0_3(horizontal_tile_13_1_to_tile_13_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(417)
	);

	pe_tile pe_tile_13_1(
		.out_wire_3_0(vertical_tile_13_1_to_tile_12_1_0),
		.out_wire_3_1(vertical_tile_13_1_to_tile_12_1_1),
		.out_wire_3_2(vertical_tile_13_1_to_tile_12_1_2),
		.out_wire_3_3(vertical_tile_13_1_to_tile_12_1_3),
		.in_wire_3_0(vertical_tile_12_1_to_tile_13_1_0),
		.in_wire_3_1(vertical_tile_12_1_to_tile_13_1_1),
		.in_wire_3_2(vertical_tile_12_1_to_tile_13_1_2),
		.in_wire_3_3(vertical_tile_12_1_to_tile_13_1_3),
		.out_wire_1_0(vertical_tile_13_1_to_tile_14_1_0),
		.out_wire_1_1(vertical_tile_13_1_to_tile_14_1_1),
		.out_wire_1_2(vertical_tile_13_1_to_tile_14_1_2),
		.out_wire_1_3(vertical_tile_13_1_to_tile_14_1_3),
		.in_wire_1_0(vertical_tile_14_1_to_tile_13_1_0),
		.in_wire_1_1(vertical_tile_14_1_to_tile_13_1_1),
		.in_wire_1_2(vertical_tile_14_1_to_tile_13_1_2),
		.in_wire_1_3(vertical_tile_14_1_to_tile_13_1_3),
		.out_wire_2_0(horizontal_tile_13_1_to_tile_13_0_0),
		.out_wire_2_1(horizontal_tile_13_1_to_tile_13_0_1),
		.out_wire_2_2(horizontal_tile_13_1_to_tile_13_0_2),
		.out_wire_2_3(horizontal_tile_13_1_to_tile_13_0_3),
		.in_wire_2_0(horizontal_tile_13_0_to_tile_13_1_0),
		.in_wire_2_1(horizontal_tile_13_0_to_tile_13_1_1),
		.in_wire_2_2(horizontal_tile_13_0_to_tile_13_1_2),
		.in_wire_2_3(horizontal_tile_13_0_to_tile_13_1_3),
		.out_wire_0_0(horizontal_tile_13_1_to_tile_13_2_0),
		.out_wire_0_1(horizontal_tile_13_1_to_tile_13_2_1),
		.out_wire_0_2(horizontal_tile_13_1_to_tile_13_2_2),
		.out_wire_0_3(horizontal_tile_13_1_to_tile_13_2_3),
		.in_wire_0_0(horizontal_tile_13_2_to_tile_13_1_0),
		.in_wire_0_1(horizontal_tile_13_2_to_tile_13_1_1),
		.in_wire_0_2(horizontal_tile_13_2_to_tile_13_1_2),
		.in_wire_0_3(horizontal_tile_13_2_to_tile_13_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(418)
	);

	pe_tile pe_tile_13_2(
		.out_wire_3_0(vertical_tile_13_2_to_tile_12_2_0),
		.out_wire_3_1(vertical_tile_13_2_to_tile_12_2_1),
		.out_wire_3_2(vertical_tile_13_2_to_tile_12_2_2),
		.out_wire_3_3(vertical_tile_13_2_to_tile_12_2_3),
		.in_wire_3_0(vertical_tile_12_2_to_tile_13_2_0),
		.in_wire_3_1(vertical_tile_12_2_to_tile_13_2_1),
		.in_wire_3_2(vertical_tile_12_2_to_tile_13_2_2),
		.in_wire_3_3(vertical_tile_12_2_to_tile_13_2_3),
		.out_wire_1_0(vertical_tile_13_2_to_tile_14_2_0),
		.out_wire_1_1(vertical_tile_13_2_to_tile_14_2_1),
		.out_wire_1_2(vertical_tile_13_2_to_tile_14_2_2),
		.out_wire_1_3(vertical_tile_13_2_to_tile_14_2_3),
		.in_wire_1_0(vertical_tile_14_2_to_tile_13_2_0),
		.in_wire_1_1(vertical_tile_14_2_to_tile_13_2_1),
		.in_wire_1_2(vertical_tile_14_2_to_tile_13_2_2),
		.in_wire_1_3(vertical_tile_14_2_to_tile_13_2_3),
		.out_wire_2_0(horizontal_tile_13_2_to_tile_13_1_0),
		.out_wire_2_1(horizontal_tile_13_2_to_tile_13_1_1),
		.out_wire_2_2(horizontal_tile_13_2_to_tile_13_1_2),
		.out_wire_2_3(horizontal_tile_13_2_to_tile_13_1_3),
		.in_wire_2_0(horizontal_tile_13_1_to_tile_13_2_0),
		.in_wire_2_1(horizontal_tile_13_1_to_tile_13_2_1),
		.in_wire_2_2(horizontal_tile_13_1_to_tile_13_2_2),
		.in_wire_2_3(horizontal_tile_13_1_to_tile_13_2_3),
		.out_wire_0_0(horizontal_tile_13_2_to_tile_13_3_0),
		.out_wire_0_1(horizontal_tile_13_2_to_tile_13_3_1),
		.out_wire_0_2(horizontal_tile_13_2_to_tile_13_3_2),
		.out_wire_0_3(horizontal_tile_13_2_to_tile_13_3_3),
		.in_wire_0_0(horizontal_tile_13_3_to_tile_13_2_0),
		.in_wire_0_1(horizontal_tile_13_3_to_tile_13_2_1),
		.in_wire_0_2(horizontal_tile_13_3_to_tile_13_2_2),
		.in_wire_0_3(horizontal_tile_13_3_to_tile_13_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(419)
	);

	pe_tile pe_tile_13_3(
		.out_wire_3_0(vertical_tile_13_3_to_tile_12_3_0),
		.out_wire_3_1(vertical_tile_13_3_to_tile_12_3_1),
		.out_wire_3_2(vertical_tile_13_3_to_tile_12_3_2),
		.out_wire_3_3(vertical_tile_13_3_to_tile_12_3_3),
		.in_wire_3_0(vertical_tile_12_3_to_tile_13_3_0),
		.in_wire_3_1(vertical_tile_12_3_to_tile_13_3_1),
		.in_wire_3_2(vertical_tile_12_3_to_tile_13_3_2),
		.in_wire_3_3(vertical_tile_12_3_to_tile_13_3_3),
		.out_wire_1_0(vertical_tile_13_3_to_tile_14_3_0),
		.out_wire_1_1(vertical_tile_13_3_to_tile_14_3_1),
		.out_wire_1_2(vertical_tile_13_3_to_tile_14_3_2),
		.out_wire_1_3(vertical_tile_13_3_to_tile_14_3_3),
		.in_wire_1_0(vertical_tile_14_3_to_tile_13_3_0),
		.in_wire_1_1(vertical_tile_14_3_to_tile_13_3_1),
		.in_wire_1_2(vertical_tile_14_3_to_tile_13_3_2),
		.in_wire_1_3(vertical_tile_14_3_to_tile_13_3_3),
		.out_wire_2_0(horizontal_tile_13_3_to_tile_13_2_0),
		.out_wire_2_1(horizontal_tile_13_3_to_tile_13_2_1),
		.out_wire_2_2(horizontal_tile_13_3_to_tile_13_2_2),
		.out_wire_2_3(horizontal_tile_13_3_to_tile_13_2_3),
		.in_wire_2_0(horizontal_tile_13_2_to_tile_13_3_0),
		.in_wire_2_1(horizontal_tile_13_2_to_tile_13_3_1),
		.in_wire_2_2(horizontal_tile_13_2_to_tile_13_3_2),
		.in_wire_2_3(horizontal_tile_13_2_to_tile_13_3_3),
		.out_wire_0_0(horizontal_tile_13_3_to_tile_13_4_0),
		.out_wire_0_1(horizontal_tile_13_3_to_tile_13_4_1),
		.out_wire_0_2(horizontal_tile_13_3_to_tile_13_4_2),
		.out_wire_0_3(horizontal_tile_13_3_to_tile_13_4_3),
		.in_wire_0_0(horizontal_tile_13_4_to_tile_13_3_0),
		.in_wire_0_1(horizontal_tile_13_4_to_tile_13_3_1),
		.in_wire_0_2(horizontal_tile_13_4_to_tile_13_3_2),
		.in_wire_0_3(horizontal_tile_13_4_to_tile_13_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(420)
	);

	pe_tile pe_tile_13_4(
		.out_wire_3_0(vertical_tile_13_4_to_tile_12_4_0),
		.out_wire_3_1(vertical_tile_13_4_to_tile_12_4_1),
		.out_wire_3_2(vertical_tile_13_4_to_tile_12_4_2),
		.out_wire_3_3(vertical_tile_13_4_to_tile_12_4_3),
		.in_wire_3_0(vertical_tile_12_4_to_tile_13_4_0),
		.in_wire_3_1(vertical_tile_12_4_to_tile_13_4_1),
		.in_wire_3_2(vertical_tile_12_4_to_tile_13_4_2),
		.in_wire_3_3(vertical_tile_12_4_to_tile_13_4_3),
		.out_wire_1_0(vertical_tile_13_4_to_tile_14_4_0),
		.out_wire_1_1(vertical_tile_13_4_to_tile_14_4_1),
		.out_wire_1_2(vertical_tile_13_4_to_tile_14_4_2),
		.out_wire_1_3(vertical_tile_13_4_to_tile_14_4_3),
		.in_wire_1_0(vertical_tile_14_4_to_tile_13_4_0),
		.in_wire_1_1(vertical_tile_14_4_to_tile_13_4_1),
		.in_wire_1_2(vertical_tile_14_4_to_tile_13_4_2),
		.in_wire_1_3(vertical_tile_14_4_to_tile_13_4_3),
		.out_wire_2_0(horizontal_tile_13_4_to_tile_13_3_0),
		.out_wire_2_1(horizontal_tile_13_4_to_tile_13_3_1),
		.out_wire_2_2(horizontal_tile_13_4_to_tile_13_3_2),
		.out_wire_2_3(horizontal_tile_13_4_to_tile_13_3_3),
		.in_wire_2_0(horizontal_tile_13_3_to_tile_13_4_0),
		.in_wire_2_1(horizontal_tile_13_3_to_tile_13_4_1),
		.in_wire_2_2(horizontal_tile_13_3_to_tile_13_4_2),
		.in_wire_2_3(horizontal_tile_13_3_to_tile_13_4_3),
		.out_wire_0_0(horizontal_tile_13_4_to_tile_13_5_0),
		.out_wire_0_1(horizontal_tile_13_4_to_tile_13_5_1),
		.out_wire_0_2(horizontal_tile_13_4_to_tile_13_5_2),
		.out_wire_0_3(horizontal_tile_13_4_to_tile_13_5_3),
		.in_wire_0_0(horizontal_tile_13_5_to_tile_13_4_0),
		.in_wire_0_1(horizontal_tile_13_5_to_tile_13_4_1),
		.in_wire_0_2(horizontal_tile_13_5_to_tile_13_4_2),
		.in_wire_0_3(horizontal_tile_13_5_to_tile_13_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(421)
	);

	pe_tile pe_tile_13_5(
		.out_wire_3_0(vertical_tile_13_5_to_tile_12_5_0),
		.out_wire_3_1(vertical_tile_13_5_to_tile_12_5_1),
		.out_wire_3_2(vertical_tile_13_5_to_tile_12_5_2),
		.out_wire_3_3(vertical_tile_13_5_to_tile_12_5_3),
		.in_wire_3_0(vertical_tile_12_5_to_tile_13_5_0),
		.in_wire_3_1(vertical_tile_12_5_to_tile_13_5_1),
		.in_wire_3_2(vertical_tile_12_5_to_tile_13_5_2),
		.in_wire_3_3(vertical_tile_12_5_to_tile_13_5_3),
		.out_wire_1_0(vertical_tile_13_5_to_tile_14_5_0),
		.out_wire_1_1(vertical_tile_13_5_to_tile_14_5_1),
		.out_wire_1_2(vertical_tile_13_5_to_tile_14_5_2),
		.out_wire_1_3(vertical_tile_13_5_to_tile_14_5_3),
		.in_wire_1_0(vertical_tile_14_5_to_tile_13_5_0),
		.in_wire_1_1(vertical_tile_14_5_to_tile_13_5_1),
		.in_wire_1_2(vertical_tile_14_5_to_tile_13_5_2),
		.in_wire_1_3(vertical_tile_14_5_to_tile_13_5_3),
		.out_wire_2_0(horizontal_tile_13_5_to_tile_13_4_0),
		.out_wire_2_1(horizontal_tile_13_5_to_tile_13_4_1),
		.out_wire_2_2(horizontal_tile_13_5_to_tile_13_4_2),
		.out_wire_2_3(horizontal_tile_13_5_to_tile_13_4_3),
		.in_wire_2_0(horizontal_tile_13_4_to_tile_13_5_0),
		.in_wire_2_1(horizontal_tile_13_4_to_tile_13_5_1),
		.in_wire_2_2(horizontal_tile_13_4_to_tile_13_5_2),
		.in_wire_2_3(horizontal_tile_13_4_to_tile_13_5_3),
		.out_wire_0_0(horizontal_tile_13_5_to_tile_13_6_0),
		.out_wire_0_1(horizontal_tile_13_5_to_tile_13_6_1),
		.out_wire_0_2(horizontal_tile_13_5_to_tile_13_6_2),
		.out_wire_0_3(horizontal_tile_13_5_to_tile_13_6_3),
		.in_wire_0_0(horizontal_tile_13_6_to_tile_13_5_0),
		.in_wire_0_1(horizontal_tile_13_6_to_tile_13_5_1),
		.in_wire_0_2(horizontal_tile_13_6_to_tile_13_5_2),
		.in_wire_0_3(horizontal_tile_13_6_to_tile_13_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(422)
	);

	pe_tile pe_tile_13_6(
		.out_wire_3_0(vertical_tile_13_6_to_tile_12_6_0),
		.out_wire_3_1(vertical_tile_13_6_to_tile_12_6_1),
		.out_wire_3_2(vertical_tile_13_6_to_tile_12_6_2),
		.out_wire_3_3(vertical_tile_13_6_to_tile_12_6_3),
		.in_wire_3_0(vertical_tile_12_6_to_tile_13_6_0),
		.in_wire_3_1(vertical_tile_12_6_to_tile_13_6_1),
		.in_wire_3_2(vertical_tile_12_6_to_tile_13_6_2),
		.in_wire_3_3(vertical_tile_12_6_to_tile_13_6_3),
		.out_wire_1_0(vertical_tile_13_6_to_tile_14_6_0),
		.out_wire_1_1(vertical_tile_13_6_to_tile_14_6_1),
		.out_wire_1_2(vertical_tile_13_6_to_tile_14_6_2),
		.out_wire_1_3(vertical_tile_13_6_to_tile_14_6_3),
		.in_wire_1_0(vertical_tile_14_6_to_tile_13_6_0),
		.in_wire_1_1(vertical_tile_14_6_to_tile_13_6_1),
		.in_wire_1_2(vertical_tile_14_6_to_tile_13_6_2),
		.in_wire_1_3(vertical_tile_14_6_to_tile_13_6_3),
		.out_wire_2_0(horizontal_tile_13_6_to_tile_13_5_0),
		.out_wire_2_1(horizontal_tile_13_6_to_tile_13_5_1),
		.out_wire_2_2(horizontal_tile_13_6_to_tile_13_5_2),
		.out_wire_2_3(horizontal_tile_13_6_to_tile_13_5_3),
		.in_wire_2_0(horizontal_tile_13_5_to_tile_13_6_0),
		.in_wire_2_1(horizontal_tile_13_5_to_tile_13_6_1),
		.in_wire_2_2(horizontal_tile_13_5_to_tile_13_6_2),
		.in_wire_2_3(horizontal_tile_13_5_to_tile_13_6_3),
		.out_wire_0_0(horizontal_tile_13_6_to_tile_13_7_0),
		.out_wire_0_1(horizontal_tile_13_6_to_tile_13_7_1),
		.out_wire_0_2(horizontal_tile_13_6_to_tile_13_7_2),
		.out_wire_0_3(horizontal_tile_13_6_to_tile_13_7_3),
		.in_wire_0_0(horizontal_tile_13_7_to_tile_13_6_0),
		.in_wire_0_1(horizontal_tile_13_7_to_tile_13_6_1),
		.in_wire_0_2(horizontal_tile_13_7_to_tile_13_6_2),
		.in_wire_0_3(horizontal_tile_13_7_to_tile_13_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(423)
	);

	pe_tile pe_tile_13_7(
		.out_wire_3_0(vertical_tile_13_7_to_tile_12_7_0),
		.out_wire_3_1(vertical_tile_13_7_to_tile_12_7_1),
		.out_wire_3_2(vertical_tile_13_7_to_tile_12_7_2),
		.out_wire_3_3(vertical_tile_13_7_to_tile_12_7_3),
		.in_wire_3_0(vertical_tile_12_7_to_tile_13_7_0),
		.in_wire_3_1(vertical_tile_12_7_to_tile_13_7_1),
		.in_wire_3_2(vertical_tile_12_7_to_tile_13_7_2),
		.in_wire_3_3(vertical_tile_12_7_to_tile_13_7_3),
		.out_wire_1_0(vertical_tile_13_7_to_tile_14_7_0),
		.out_wire_1_1(vertical_tile_13_7_to_tile_14_7_1),
		.out_wire_1_2(vertical_tile_13_7_to_tile_14_7_2),
		.out_wire_1_3(vertical_tile_13_7_to_tile_14_7_3),
		.in_wire_1_0(vertical_tile_14_7_to_tile_13_7_0),
		.in_wire_1_1(vertical_tile_14_7_to_tile_13_7_1),
		.in_wire_1_2(vertical_tile_14_7_to_tile_13_7_2),
		.in_wire_1_3(vertical_tile_14_7_to_tile_13_7_3),
		.out_wire_2_0(horizontal_tile_13_7_to_tile_13_6_0),
		.out_wire_2_1(horizontal_tile_13_7_to_tile_13_6_1),
		.out_wire_2_2(horizontal_tile_13_7_to_tile_13_6_2),
		.out_wire_2_3(horizontal_tile_13_7_to_tile_13_6_3),
		.in_wire_2_0(horizontal_tile_13_6_to_tile_13_7_0),
		.in_wire_2_1(horizontal_tile_13_6_to_tile_13_7_1),
		.in_wire_2_2(horizontal_tile_13_6_to_tile_13_7_2),
		.in_wire_2_3(horizontal_tile_13_6_to_tile_13_7_3),
		.out_wire_0_0(horizontal_tile_13_7_to_tile_13_8_0),
		.out_wire_0_1(horizontal_tile_13_7_to_tile_13_8_1),
		.out_wire_0_2(horizontal_tile_13_7_to_tile_13_8_2),
		.out_wire_0_3(horizontal_tile_13_7_to_tile_13_8_3),
		.in_wire_0_0(horizontal_tile_13_8_to_tile_13_7_0),
		.in_wire_0_1(horizontal_tile_13_8_to_tile_13_7_1),
		.in_wire_0_2(horizontal_tile_13_8_to_tile_13_7_2),
		.in_wire_0_3(horizontal_tile_13_8_to_tile_13_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(424)
	);

	pe_tile pe_tile_13_8(
		.out_wire_3_0(vertical_tile_13_8_to_tile_12_8_0),
		.out_wire_3_1(vertical_tile_13_8_to_tile_12_8_1),
		.out_wire_3_2(vertical_tile_13_8_to_tile_12_8_2),
		.out_wire_3_3(vertical_tile_13_8_to_tile_12_8_3),
		.in_wire_3_0(vertical_tile_12_8_to_tile_13_8_0),
		.in_wire_3_1(vertical_tile_12_8_to_tile_13_8_1),
		.in_wire_3_2(vertical_tile_12_8_to_tile_13_8_2),
		.in_wire_3_3(vertical_tile_12_8_to_tile_13_8_3),
		.out_wire_1_0(vertical_tile_13_8_to_tile_14_8_0),
		.out_wire_1_1(vertical_tile_13_8_to_tile_14_8_1),
		.out_wire_1_2(vertical_tile_13_8_to_tile_14_8_2),
		.out_wire_1_3(vertical_tile_13_8_to_tile_14_8_3),
		.in_wire_1_0(vertical_tile_14_8_to_tile_13_8_0),
		.in_wire_1_1(vertical_tile_14_8_to_tile_13_8_1),
		.in_wire_1_2(vertical_tile_14_8_to_tile_13_8_2),
		.in_wire_1_3(vertical_tile_14_8_to_tile_13_8_3),
		.out_wire_2_0(horizontal_tile_13_8_to_tile_13_7_0),
		.out_wire_2_1(horizontal_tile_13_8_to_tile_13_7_1),
		.out_wire_2_2(horizontal_tile_13_8_to_tile_13_7_2),
		.out_wire_2_3(horizontal_tile_13_8_to_tile_13_7_3),
		.in_wire_2_0(horizontal_tile_13_7_to_tile_13_8_0),
		.in_wire_2_1(horizontal_tile_13_7_to_tile_13_8_1),
		.in_wire_2_2(horizontal_tile_13_7_to_tile_13_8_2),
		.in_wire_2_3(horizontal_tile_13_7_to_tile_13_8_3),
		.out_wire_0_0(horizontal_tile_13_8_to_tile_13_9_0),
		.out_wire_0_1(horizontal_tile_13_8_to_tile_13_9_1),
		.out_wire_0_2(horizontal_tile_13_8_to_tile_13_9_2),
		.out_wire_0_3(horizontal_tile_13_8_to_tile_13_9_3),
		.in_wire_0_0(horizontal_tile_13_9_to_tile_13_8_0),
		.in_wire_0_1(horizontal_tile_13_9_to_tile_13_8_1),
		.in_wire_0_2(horizontal_tile_13_9_to_tile_13_8_2),
		.in_wire_0_3(horizontal_tile_13_9_to_tile_13_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(425)
	);

	pe_tile pe_tile_13_9(
		.out_wire_3_0(vertical_tile_13_9_to_tile_12_9_0),
		.out_wire_3_1(vertical_tile_13_9_to_tile_12_9_1),
		.out_wire_3_2(vertical_tile_13_9_to_tile_12_9_2),
		.out_wire_3_3(vertical_tile_13_9_to_tile_12_9_3),
		.in_wire_3_0(vertical_tile_12_9_to_tile_13_9_0),
		.in_wire_3_1(vertical_tile_12_9_to_tile_13_9_1),
		.in_wire_3_2(vertical_tile_12_9_to_tile_13_9_2),
		.in_wire_3_3(vertical_tile_12_9_to_tile_13_9_3),
		.out_wire_1_0(vertical_tile_13_9_to_tile_14_9_0),
		.out_wire_1_1(vertical_tile_13_9_to_tile_14_9_1),
		.out_wire_1_2(vertical_tile_13_9_to_tile_14_9_2),
		.out_wire_1_3(vertical_tile_13_9_to_tile_14_9_3),
		.in_wire_1_0(vertical_tile_14_9_to_tile_13_9_0),
		.in_wire_1_1(vertical_tile_14_9_to_tile_13_9_1),
		.in_wire_1_2(vertical_tile_14_9_to_tile_13_9_2),
		.in_wire_1_3(vertical_tile_14_9_to_tile_13_9_3),
		.out_wire_2_0(horizontal_tile_13_9_to_tile_13_8_0),
		.out_wire_2_1(horizontal_tile_13_9_to_tile_13_8_1),
		.out_wire_2_2(horizontal_tile_13_9_to_tile_13_8_2),
		.out_wire_2_3(horizontal_tile_13_9_to_tile_13_8_3),
		.in_wire_2_0(horizontal_tile_13_8_to_tile_13_9_0),
		.in_wire_2_1(horizontal_tile_13_8_to_tile_13_9_1),
		.in_wire_2_2(horizontal_tile_13_8_to_tile_13_9_2),
		.in_wire_2_3(horizontal_tile_13_8_to_tile_13_9_3),
		.out_wire_0_0(horizontal_tile_13_9_to_tile_13_10_0),
		.out_wire_0_1(horizontal_tile_13_9_to_tile_13_10_1),
		.out_wire_0_2(horizontal_tile_13_9_to_tile_13_10_2),
		.out_wire_0_3(horizontal_tile_13_9_to_tile_13_10_3),
		.in_wire_0_0(horizontal_tile_13_10_to_tile_13_9_0),
		.in_wire_0_1(horizontal_tile_13_10_to_tile_13_9_1),
		.in_wire_0_2(horizontal_tile_13_10_to_tile_13_9_2),
		.in_wire_0_3(horizontal_tile_13_10_to_tile_13_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(426)
	);

	pe_tile pe_tile_13_10(
		.out_wire_3_0(vertical_tile_13_10_to_tile_12_10_0),
		.out_wire_3_1(vertical_tile_13_10_to_tile_12_10_1),
		.out_wire_3_2(vertical_tile_13_10_to_tile_12_10_2),
		.out_wire_3_3(vertical_tile_13_10_to_tile_12_10_3),
		.in_wire_3_0(vertical_tile_12_10_to_tile_13_10_0),
		.in_wire_3_1(vertical_tile_12_10_to_tile_13_10_1),
		.in_wire_3_2(vertical_tile_12_10_to_tile_13_10_2),
		.in_wire_3_3(vertical_tile_12_10_to_tile_13_10_3),
		.out_wire_1_0(vertical_tile_13_10_to_tile_14_10_0),
		.out_wire_1_1(vertical_tile_13_10_to_tile_14_10_1),
		.out_wire_1_2(vertical_tile_13_10_to_tile_14_10_2),
		.out_wire_1_3(vertical_tile_13_10_to_tile_14_10_3),
		.in_wire_1_0(vertical_tile_14_10_to_tile_13_10_0),
		.in_wire_1_1(vertical_tile_14_10_to_tile_13_10_1),
		.in_wire_1_2(vertical_tile_14_10_to_tile_13_10_2),
		.in_wire_1_3(vertical_tile_14_10_to_tile_13_10_3),
		.out_wire_2_0(horizontal_tile_13_10_to_tile_13_9_0),
		.out_wire_2_1(horizontal_tile_13_10_to_tile_13_9_1),
		.out_wire_2_2(horizontal_tile_13_10_to_tile_13_9_2),
		.out_wire_2_3(horizontal_tile_13_10_to_tile_13_9_3),
		.in_wire_2_0(horizontal_tile_13_9_to_tile_13_10_0),
		.in_wire_2_1(horizontal_tile_13_9_to_tile_13_10_1),
		.in_wire_2_2(horizontal_tile_13_9_to_tile_13_10_2),
		.in_wire_2_3(horizontal_tile_13_9_to_tile_13_10_3),
		.out_wire_0_0(horizontal_tile_13_10_to_tile_13_11_0),
		.out_wire_0_1(horizontal_tile_13_10_to_tile_13_11_1),
		.out_wire_0_2(horizontal_tile_13_10_to_tile_13_11_2),
		.out_wire_0_3(horizontal_tile_13_10_to_tile_13_11_3),
		.in_wire_0_0(horizontal_tile_13_11_to_tile_13_10_0),
		.in_wire_0_1(horizontal_tile_13_11_to_tile_13_10_1),
		.in_wire_0_2(horizontal_tile_13_11_to_tile_13_10_2),
		.in_wire_0_3(horizontal_tile_13_11_to_tile_13_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(427)
	);

	pe_tile pe_tile_13_11(
		.out_wire_3_0(vertical_tile_13_11_to_tile_12_11_0),
		.out_wire_3_1(vertical_tile_13_11_to_tile_12_11_1),
		.out_wire_3_2(vertical_tile_13_11_to_tile_12_11_2),
		.out_wire_3_3(vertical_tile_13_11_to_tile_12_11_3),
		.in_wire_3_0(vertical_tile_12_11_to_tile_13_11_0),
		.in_wire_3_1(vertical_tile_12_11_to_tile_13_11_1),
		.in_wire_3_2(vertical_tile_12_11_to_tile_13_11_2),
		.in_wire_3_3(vertical_tile_12_11_to_tile_13_11_3),
		.out_wire_1_0(vertical_tile_13_11_to_tile_14_11_0),
		.out_wire_1_1(vertical_tile_13_11_to_tile_14_11_1),
		.out_wire_1_2(vertical_tile_13_11_to_tile_14_11_2),
		.out_wire_1_3(vertical_tile_13_11_to_tile_14_11_3),
		.in_wire_1_0(vertical_tile_14_11_to_tile_13_11_0),
		.in_wire_1_1(vertical_tile_14_11_to_tile_13_11_1),
		.in_wire_1_2(vertical_tile_14_11_to_tile_13_11_2),
		.in_wire_1_3(vertical_tile_14_11_to_tile_13_11_3),
		.out_wire_2_0(horizontal_tile_13_11_to_tile_13_10_0),
		.out_wire_2_1(horizontal_tile_13_11_to_tile_13_10_1),
		.out_wire_2_2(horizontal_tile_13_11_to_tile_13_10_2),
		.out_wire_2_3(horizontal_tile_13_11_to_tile_13_10_3),
		.in_wire_2_0(horizontal_tile_13_10_to_tile_13_11_0),
		.in_wire_2_1(horizontal_tile_13_10_to_tile_13_11_1),
		.in_wire_2_2(horizontal_tile_13_10_to_tile_13_11_2),
		.in_wire_2_3(horizontal_tile_13_10_to_tile_13_11_3),
		.out_wire_0_0(horizontal_tile_13_11_to_tile_13_12_0),
		.out_wire_0_1(horizontal_tile_13_11_to_tile_13_12_1),
		.out_wire_0_2(horizontal_tile_13_11_to_tile_13_12_2),
		.out_wire_0_3(horizontal_tile_13_11_to_tile_13_12_3),
		.in_wire_0_0(horizontal_tile_13_12_to_tile_13_11_0),
		.in_wire_0_1(horizontal_tile_13_12_to_tile_13_11_1),
		.in_wire_0_2(horizontal_tile_13_12_to_tile_13_11_2),
		.in_wire_0_3(horizontal_tile_13_12_to_tile_13_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(428)
	);

	pe_tile pe_tile_13_12(
		.out_wire_3_0(vertical_tile_13_12_to_tile_12_12_0),
		.out_wire_3_1(vertical_tile_13_12_to_tile_12_12_1),
		.out_wire_3_2(vertical_tile_13_12_to_tile_12_12_2),
		.out_wire_3_3(vertical_tile_13_12_to_tile_12_12_3),
		.in_wire_3_0(vertical_tile_12_12_to_tile_13_12_0),
		.in_wire_3_1(vertical_tile_12_12_to_tile_13_12_1),
		.in_wire_3_2(vertical_tile_12_12_to_tile_13_12_2),
		.in_wire_3_3(vertical_tile_12_12_to_tile_13_12_3),
		.out_wire_1_0(vertical_tile_13_12_to_tile_14_12_0),
		.out_wire_1_1(vertical_tile_13_12_to_tile_14_12_1),
		.out_wire_1_2(vertical_tile_13_12_to_tile_14_12_2),
		.out_wire_1_3(vertical_tile_13_12_to_tile_14_12_3),
		.in_wire_1_0(vertical_tile_14_12_to_tile_13_12_0),
		.in_wire_1_1(vertical_tile_14_12_to_tile_13_12_1),
		.in_wire_1_2(vertical_tile_14_12_to_tile_13_12_2),
		.in_wire_1_3(vertical_tile_14_12_to_tile_13_12_3),
		.out_wire_2_0(horizontal_tile_13_12_to_tile_13_11_0),
		.out_wire_2_1(horizontal_tile_13_12_to_tile_13_11_1),
		.out_wire_2_2(horizontal_tile_13_12_to_tile_13_11_2),
		.out_wire_2_3(horizontal_tile_13_12_to_tile_13_11_3),
		.in_wire_2_0(horizontal_tile_13_11_to_tile_13_12_0),
		.in_wire_2_1(horizontal_tile_13_11_to_tile_13_12_1),
		.in_wire_2_2(horizontal_tile_13_11_to_tile_13_12_2),
		.in_wire_2_3(horizontal_tile_13_11_to_tile_13_12_3),
		.out_wire_0_0(horizontal_tile_13_12_to_tile_13_13_0),
		.out_wire_0_1(horizontal_tile_13_12_to_tile_13_13_1),
		.out_wire_0_2(horizontal_tile_13_12_to_tile_13_13_2),
		.out_wire_0_3(horizontal_tile_13_12_to_tile_13_13_3),
		.in_wire_0_0(horizontal_tile_13_13_to_tile_13_12_0),
		.in_wire_0_1(horizontal_tile_13_13_to_tile_13_12_1),
		.in_wire_0_2(horizontal_tile_13_13_to_tile_13_12_2),
		.in_wire_0_3(horizontal_tile_13_13_to_tile_13_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(429)
	);

	pe_tile pe_tile_13_13(
		.out_wire_3_0(vertical_tile_13_13_to_tile_12_13_0),
		.out_wire_3_1(vertical_tile_13_13_to_tile_12_13_1),
		.out_wire_3_2(vertical_tile_13_13_to_tile_12_13_2),
		.out_wire_3_3(vertical_tile_13_13_to_tile_12_13_3),
		.in_wire_3_0(vertical_tile_12_13_to_tile_13_13_0),
		.in_wire_3_1(vertical_tile_12_13_to_tile_13_13_1),
		.in_wire_3_2(vertical_tile_12_13_to_tile_13_13_2),
		.in_wire_3_3(vertical_tile_12_13_to_tile_13_13_3),
		.out_wire_1_0(vertical_tile_13_13_to_tile_14_13_0),
		.out_wire_1_1(vertical_tile_13_13_to_tile_14_13_1),
		.out_wire_1_2(vertical_tile_13_13_to_tile_14_13_2),
		.out_wire_1_3(vertical_tile_13_13_to_tile_14_13_3),
		.in_wire_1_0(vertical_tile_14_13_to_tile_13_13_0),
		.in_wire_1_1(vertical_tile_14_13_to_tile_13_13_1),
		.in_wire_1_2(vertical_tile_14_13_to_tile_13_13_2),
		.in_wire_1_3(vertical_tile_14_13_to_tile_13_13_3),
		.out_wire_2_0(horizontal_tile_13_13_to_tile_13_12_0),
		.out_wire_2_1(horizontal_tile_13_13_to_tile_13_12_1),
		.out_wire_2_2(horizontal_tile_13_13_to_tile_13_12_2),
		.out_wire_2_3(horizontal_tile_13_13_to_tile_13_12_3),
		.in_wire_2_0(horizontal_tile_13_12_to_tile_13_13_0),
		.in_wire_2_1(horizontal_tile_13_12_to_tile_13_13_1),
		.in_wire_2_2(horizontal_tile_13_12_to_tile_13_13_2),
		.in_wire_2_3(horizontal_tile_13_12_to_tile_13_13_3),
		.out_wire_0_0(horizontal_tile_13_13_to_tile_13_14_0),
		.out_wire_0_1(horizontal_tile_13_13_to_tile_13_14_1),
		.out_wire_0_2(horizontal_tile_13_13_to_tile_13_14_2),
		.out_wire_0_3(horizontal_tile_13_13_to_tile_13_14_3),
		.in_wire_0_0(horizontal_tile_13_14_to_tile_13_13_0),
		.in_wire_0_1(horizontal_tile_13_14_to_tile_13_13_1),
		.in_wire_0_2(horizontal_tile_13_14_to_tile_13_13_2),
		.in_wire_0_3(horizontal_tile_13_14_to_tile_13_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(430)
	);

	pe_tile pe_tile_13_14(
		.out_wire_3_0(vertical_tile_13_14_to_tile_12_14_0),
		.out_wire_3_1(vertical_tile_13_14_to_tile_12_14_1),
		.out_wire_3_2(vertical_tile_13_14_to_tile_12_14_2),
		.out_wire_3_3(vertical_tile_13_14_to_tile_12_14_3),
		.in_wire_3_0(vertical_tile_12_14_to_tile_13_14_0),
		.in_wire_3_1(vertical_tile_12_14_to_tile_13_14_1),
		.in_wire_3_2(vertical_tile_12_14_to_tile_13_14_2),
		.in_wire_3_3(vertical_tile_12_14_to_tile_13_14_3),
		.out_wire_1_0(vertical_tile_13_14_to_tile_14_14_0),
		.out_wire_1_1(vertical_tile_13_14_to_tile_14_14_1),
		.out_wire_1_2(vertical_tile_13_14_to_tile_14_14_2),
		.out_wire_1_3(vertical_tile_13_14_to_tile_14_14_3),
		.in_wire_1_0(vertical_tile_14_14_to_tile_13_14_0),
		.in_wire_1_1(vertical_tile_14_14_to_tile_13_14_1),
		.in_wire_1_2(vertical_tile_14_14_to_tile_13_14_2),
		.in_wire_1_3(vertical_tile_14_14_to_tile_13_14_3),
		.out_wire_2_0(horizontal_tile_13_14_to_tile_13_13_0),
		.out_wire_2_1(horizontal_tile_13_14_to_tile_13_13_1),
		.out_wire_2_2(horizontal_tile_13_14_to_tile_13_13_2),
		.out_wire_2_3(horizontal_tile_13_14_to_tile_13_13_3),
		.in_wire_2_0(horizontal_tile_13_13_to_tile_13_14_0),
		.in_wire_2_1(horizontal_tile_13_13_to_tile_13_14_1),
		.in_wire_2_2(horizontal_tile_13_13_to_tile_13_14_2),
		.in_wire_2_3(horizontal_tile_13_13_to_tile_13_14_3),
		.out_wire_0_0(horizontal_tile_13_14_to_tile_13_15_0),
		.out_wire_0_1(horizontal_tile_13_14_to_tile_13_15_1),
		.out_wire_0_2(horizontal_tile_13_14_to_tile_13_15_2),
		.out_wire_0_3(horizontal_tile_13_14_to_tile_13_15_3),
		.in_wire_0_0(horizontal_tile_13_15_to_tile_13_14_0),
		.in_wire_0_1(horizontal_tile_13_15_to_tile_13_14_1),
		.in_wire_0_2(horizontal_tile_13_15_to_tile_13_14_2),
		.in_wire_0_3(horizontal_tile_13_15_to_tile_13_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(431)
	);

	pe_tile pe_tile_13_15(
		.out_wire_3_0(vertical_tile_13_15_to_tile_12_15_0),
		.out_wire_3_1(vertical_tile_13_15_to_tile_12_15_1),
		.out_wire_3_2(vertical_tile_13_15_to_tile_12_15_2),
		.out_wire_3_3(vertical_tile_13_15_to_tile_12_15_3),
		.in_wire_3_0(vertical_tile_12_15_to_tile_13_15_0),
		.in_wire_3_1(vertical_tile_12_15_to_tile_13_15_1),
		.in_wire_3_2(vertical_tile_12_15_to_tile_13_15_2),
		.in_wire_3_3(vertical_tile_12_15_to_tile_13_15_3),
		.out_wire_1_0(vertical_tile_13_15_to_tile_14_15_0),
		.out_wire_1_1(vertical_tile_13_15_to_tile_14_15_1),
		.out_wire_1_2(vertical_tile_13_15_to_tile_14_15_2),
		.out_wire_1_3(vertical_tile_13_15_to_tile_14_15_3),
		.in_wire_1_0(vertical_tile_14_15_to_tile_13_15_0),
		.in_wire_1_1(vertical_tile_14_15_to_tile_13_15_1),
		.in_wire_1_2(vertical_tile_14_15_to_tile_13_15_2),
		.in_wire_1_3(vertical_tile_14_15_to_tile_13_15_3),
		.out_wire_2_0(horizontal_tile_13_15_to_tile_13_14_0),
		.out_wire_2_1(horizontal_tile_13_15_to_tile_13_14_1),
		.out_wire_2_2(horizontal_tile_13_15_to_tile_13_14_2),
		.out_wire_2_3(horizontal_tile_13_15_to_tile_13_14_3),
		.in_wire_2_0(horizontal_tile_13_14_to_tile_13_15_0),
		.in_wire_2_1(horizontal_tile_13_14_to_tile_13_15_1),
		.in_wire_2_2(horizontal_tile_13_14_to_tile_13_15_2),
		.in_wire_2_3(horizontal_tile_13_14_to_tile_13_15_3),
		.out_wire_0_0(horizontal_tile_13_15_to_tile_13_16_0),
		.out_wire_0_1(horizontal_tile_13_15_to_tile_13_16_1),
		.out_wire_0_2(horizontal_tile_13_15_to_tile_13_16_2),
		.out_wire_0_3(horizontal_tile_13_15_to_tile_13_16_3),
		.in_wire_0_0(horizontal_tile_13_16_to_tile_13_15_0),
		.in_wire_0_1(horizontal_tile_13_16_to_tile_13_15_1),
		.in_wire_0_2(horizontal_tile_13_16_to_tile_13_15_2),
		.in_wire_0_3(horizontal_tile_13_16_to_tile_13_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(432)
	);

	pe_tile pe_tile_13_16(
		.out_wire_3_0(vertical_tile_13_16_to_tile_12_16_0),
		.out_wire_3_1(vertical_tile_13_16_to_tile_12_16_1),
		.out_wire_3_2(vertical_tile_13_16_to_tile_12_16_2),
		.out_wire_3_3(vertical_tile_13_16_to_tile_12_16_3),
		.in_wire_3_0(vertical_tile_12_16_to_tile_13_16_0),
		.in_wire_3_1(vertical_tile_12_16_to_tile_13_16_1),
		.in_wire_3_2(vertical_tile_12_16_to_tile_13_16_2),
		.in_wire_3_3(vertical_tile_12_16_to_tile_13_16_3),
		.out_wire_1_0(vertical_tile_13_16_to_tile_14_16_0),
		.out_wire_1_1(vertical_tile_13_16_to_tile_14_16_1),
		.out_wire_1_2(vertical_tile_13_16_to_tile_14_16_2),
		.out_wire_1_3(vertical_tile_13_16_to_tile_14_16_3),
		.in_wire_1_0(vertical_tile_14_16_to_tile_13_16_0),
		.in_wire_1_1(vertical_tile_14_16_to_tile_13_16_1),
		.in_wire_1_2(vertical_tile_14_16_to_tile_13_16_2),
		.in_wire_1_3(vertical_tile_14_16_to_tile_13_16_3),
		.out_wire_2_0(horizontal_tile_13_16_to_tile_13_15_0),
		.out_wire_2_1(horizontal_tile_13_16_to_tile_13_15_1),
		.out_wire_2_2(horizontal_tile_13_16_to_tile_13_15_2),
		.out_wire_2_3(horizontal_tile_13_16_to_tile_13_15_3),
		.in_wire_2_0(horizontal_tile_13_15_to_tile_13_16_0),
		.in_wire_2_1(horizontal_tile_13_15_to_tile_13_16_1),
		.in_wire_2_2(horizontal_tile_13_15_to_tile_13_16_2),
		.in_wire_2_3(horizontal_tile_13_15_to_tile_13_16_3),
		.out_wire_0_0(horizontal_tile_13_16_to_tile_13_17_0),
		.out_wire_0_1(horizontal_tile_13_16_to_tile_13_17_1),
		.out_wire_0_2(horizontal_tile_13_16_to_tile_13_17_2),
		.out_wire_0_3(horizontal_tile_13_16_to_tile_13_17_3),
		.in_wire_0_0(horizontal_tile_13_17_to_tile_13_16_0),
		.in_wire_0_1(horizontal_tile_13_17_to_tile_13_16_1),
		.in_wire_0_2(horizontal_tile_13_17_to_tile_13_16_2),
		.in_wire_0_3(horizontal_tile_13_17_to_tile_13_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(433)
	);

	pe_tile pe_tile_13_17(
		.out_wire_3_0(vertical_tile_13_17_to_tile_12_17_0),
		.out_wire_3_1(vertical_tile_13_17_to_tile_12_17_1),
		.out_wire_3_2(vertical_tile_13_17_to_tile_12_17_2),
		.out_wire_3_3(vertical_tile_13_17_to_tile_12_17_3),
		.in_wire_3_0(vertical_tile_12_17_to_tile_13_17_0),
		.in_wire_3_1(vertical_tile_12_17_to_tile_13_17_1),
		.in_wire_3_2(vertical_tile_12_17_to_tile_13_17_2),
		.in_wire_3_3(vertical_tile_12_17_to_tile_13_17_3),
		.out_wire_1_0(vertical_tile_13_17_to_tile_14_17_0),
		.out_wire_1_1(vertical_tile_13_17_to_tile_14_17_1),
		.out_wire_1_2(vertical_tile_13_17_to_tile_14_17_2),
		.out_wire_1_3(vertical_tile_13_17_to_tile_14_17_3),
		.in_wire_1_0(vertical_tile_14_17_to_tile_13_17_0),
		.in_wire_1_1(vertical_tile_14_17_to_tile_13_17_1),
		.in_wire_1_2(vertical_tile_14_17_to_tile_13_17_2),
		.in_wire_1_3(vertical_tile_14_17_to_tile_13_17_3),
		.out_wire_2_0(horizontal_tile_13_17_to_tile_13_16_0),
		.out_wire_2_1(horizontal_tile_13_17_to_tile_13_16_1),
		.out_wire_2_2(horizontal_tile_13_17_to_tile_13_16_2),
		.out_wire_2_3(horizontal_tile_13_17_to_tile_13_16_3),
		.in_wire_2_0(horizontal_tile_13_16_to_tile_13_17_0),
		.in_wire_2_1(horizontal_tile_13_16_to_tile_13_17_1),
		.in_wire_2_2(horizontal_tile_13_16_to_tile_13_17_2),
		.in_wire_2_3(horizontal_tile_13_16_to_tile_13_17_3),
		.out_wire_0_0(horizontal_tile_13_17_to_tile_13_18_0),
		.out_wire_0_1(horizontal_tile_13_17_to_tile_13_18_1),
		.out_wire_0_2(horizontal_tile_13_17_to_tile_13_18_2),
		.out_wire_0_3(horizontal_tile_13_17_to_tile_13_18_3),
		.in_wire_0_0(horizontal_tile_13_18_to_tile_13_17_0),
		.in_wire_0_1(horizontal_tile_13_18_to_tile_13_17_1),
		.in_wire_0_2(horizontal_tile_13_18_to_tile_13_17_2),
		.in_wire_0_3(horizontal_tile_13_18_to_tile_13_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(434)
	);

	pe_tile pe_tile_13_18(
		.out_wire_3_0(vertical_tile_13_18_to_tile_12_18_0),
		.out_wire_3_1(vertical_tile_13_18_to_tile_12_18_1),
		.out_wire_3_2(vertical_tile_13_18_to_tile_12_18_2),
		.out_wire_3_3(vertical_tile_13_18_to_tile_12_18_3),
		.in_wire_3_0(vertical_tile_12_18_to_tile_13_18_0),
		.in_wire_3_1(vertical_tile_12_18_to_tile_13_18_1),
		.in_wire_3_2(vertical_tile_12_18_to_tile_13_18_2),
		.in_wire_3_3(vertical_tile_12_18_to_tile_13_18_3),
		.out_wire_1_0(vertical_tile_13_18_to_tile_14_18_0),
		.out_wire_1_1(vertical_tile_13_18_to_tile_14_18_1),
		.out_wire_1_2(vertical_tile_13_18_to_tile_14_18_2),
		.out_wire_1_3(vertical_tile_13_18_to_tile_14_18_3),
		.in_wire_1_0(vertical_tile_14_18_to_tile_13_18_0),
		.in_wire_1_1(vertical_tile_14_18_to_tile_13_18_1),
		.in_wire_1_2(vertical_tile_14_18_to_tile_13_18_2),
		.in_wire_1_3(vertical_tile_14_18_to_tile_13_18_3),
		.out_wire_2_0(horizontal_tile_13_18_to_tile_13_17_0),
		.out_wire_2_1(horizontal_tile_13_18_to_tile_13_17_1),
		.out_wire_2_2(horizontal_tile_13_18_to_tile_13_17_2),
		.out_wire_2_3(horizontal_tile_13_18_to_tile_13_17_3),
		.in_wire_2_0(horizontal_tile_13_17_to_tile_13_18_0),
		.in_wire_2_1(horizontal_tile_13_17_to_tile_13_18_1),
		.in_wire_2_2(horizontal_tile_13_17_to_tile_13_18_2),
		.in_wire_2_3(horizontal_tile_13_17_to_tile_13_18_3),
		.out_wire_0_0(horizontal_tile_13_18_to_tile_13_19_0),
		.out_wire_0_1(horizontal_tile_13_18_to_tile_13_19_1),
		.out_wire_0_2(horizontal_tile_13_18_to_tile_13_19_2),
		.out_wire_0_3(horizontal_tile_13_18_to_tile_13_19_3),
		.in_wire_0_0(horizontal_tile_13_19_to_tile_13_18_0),
		.in_wire_0_1(horizontal_tile_13_19_to_tile_13_18_1),
		.in_wire_0_2(horizontal_tile_13_19_to_tile_13_18_2),
		.in_wire_0_3(horizontal_tile_13_19_to_tile_13_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(435)
	);

	pe_tile pe_tile_13_19(
		.out_wire_3_0(vertical_tile_13_19_to_tile_12_19_0),
		.out_wire_3_1(vertical_tile_13_19_to_tile_12_19_1),
		.out_wire_3_2(vertical_tile_13_19_to_tile_12_19_2),
		.out_wire_3_3(vertical_tile_13_19_to_tile_12_19_3),
		.in_wire_3_0(vertical_tile_12_19_to_tile_13_19_0),
		.in_wire_3_1(vertical_tile_12_19_to_tile_13_19_1),
		.in_wire_3_2(vertical_tile_12_19_to_tile_13_19_2),
		.in_wire_3_3(vertical_tile_12_19_to_tile_13_19_3),
		.out_wire_1_0(vertical_tile_13_19_to_tile_14_19_0),
		.out_wire_1_1(vertical_tile_13_19_to_tile_14_19_1),
		.out_wire_1_2(vertical_tile_13_19_to_tile_14_19_2),
		.out_wire_1_3(vertical_tile_13_19_to_tile_14_19_3),
		.in_wire_1_0(vertical_tile_14_19_to_tile_13_19_0),
		.in_wire_1_1(vertical_tile_14_19_to_tile_13_19_1),
		.in_wire_1_2(vertical_tile_14_19_to_tile_13_19_2),
		.in_wire_1_3(vertical_tile_14_19_to_tile_13_19_3),
		.out_wire_2_0(horizontal_tile_13_19_to_tile_13_18_0),
		.out_wire_2_1(horizontal_tile_13_19_to_tile_13_18_1),
		.out_wire_2_2(horizontal_tile_13_19_to_tile_13_18_2),
		.out_wire_2_3(horizontal_tile_13_19_to_tile_13_18_3),
		.in_wire_2_0(horizontal_tile_13_18_to_tile_13_19_0),
		.in_wire_2_1(horizontal_tile_13_18_to_tile_13_19_1),
		.in_wire_2_2(horizontal_tile_13_18_to_tile_13_19_2),
		.in_wire_2_3(horizontal_tile_13_18_to_tile_13_19_3),
		.out_wire_0_0(horizontal_tile_13_19_to_tile_13_20_0),
		.out_wire_0_1(horizontal_tile_13_19_to_tile_13_20_1),
		.out_wire_0_2(horizontal_tile_13_19_to_tile_13_20_2),
		.out_wire_0_3(horizontal_tile_13_19_to_tile_13_20_3),
		.in_wire_0_0(horizontal_tile_13_20_to_tile_13_19_0),
		.in_wire_0_1(horizontal_tile_13_20_to_tile_13_19_1),
		.in_wire_0_2(horizontal_tile_13_20_to_tile_13_19_2),
		.in_wire_0_3(horizontal_tile_13_20_to_tile_13_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(436)
	);

	pe_tile pe_tile_13_20(
		.out_wire_3_0(vertical_tile_13_20_to_tile_12_20_0),
		.out_wire_3_1(vertical_tile_13_20_to_tile_12_20_1),
		.out_wire_3_2(vertical_tile_13_20_to_tile_12_20_2),
		.out_wire_3_3(vertical_tile_13_20_to_tile_12_20_3),
		.in_wire_3_0(vertical_tile_12_20_to_tile_13_20_0),
		.in_wire_3_1(vertical_tile_12_20_to_tile_13_20_1),
		.in_wire_3_2(vertical_tile_12_20_to_tile_13_20_2),
		.in_wire_3_3(vertical_tile_12_20_to_tile_13_20_3),
		.out_wire_1_0(vertical_tile_13_20_to_tile_14_20_0),
		.out_wire_1_1(vertical_tile_13_20_to_tile_14_20_1),
		.out_wire_1_2(vertical_tile_13_20_to_tile_14_20_2),
		.out_wire_1_3(vertical_tile_13_20_to_tile_14_20_3),
		.in_wire_1_0(vertical_tile_14_20_to_tile_13_20_0),
		.in_wire_1_1(vertical_tile_14_20_to_tile_13_20_1),
		.in_wire_1_2(vertical_tile_14_20_to_tile_13_20_2),
		.in_wire_1_3(vertical_tile_14_20_to_tile_13_20_3),
		.out_wire_2_0(horizontal_tile_13_20_to_tile_13_19_0),
		.out_wire_2_1(horizontal_tile_13_20_to_tile_13_19_1),
		.out_wire_2_2(horizontal_tile_13_20_to_tile_13_19_2),
		.out_wire_2_3(horizontal_tile_13_20_to_tile_13_19_3),
		.in_wire_2_0(horizontal_tile_13_19_to_tile_13_20_0),
		.in_wire_2_1(horizontal_tile_13_19_to_tile_13_20_1),
		.in_wire_2_2(horizontal_tile_13_19_to_tile_13_20_2),
		.in_wire_2_3(horizontal_tile_13_19_to_tile_13_20_3),
		.out_wire_0_0(horizontal_tile_13_20_to_tile_13_21_0),
		.out_wire_0_1(horizontal_tile_13_20_to_tile_13_21_1),
		.out_wire_0_2(horizontal_tile_13_20_to_tile_13_21_2),
		.out_wire_0_3(horizontal_tile_13_20_to_tile_13_21_3),
		.in_wire_0_0(horizontal_tile_13_21_to_tile_13_20_0),
		.in_wire_0_1(horizontal_tile_13_21_to_tile_13_20_1),
		.in_wire_0_2(horizontal_tile_13_21_to_tile_13_20_2),
		.in_wire_0_3(horizontal_tile_13_21_to_tile_13_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(437)
	);

	pe_tile pe_tile_13_21(
		.out_wire_3_0(vertical_tile_13_21_to_tile_12_21_0),
		.out_wire_3_1(vertical_tile_13_21_to_tile_12_21_1),
		.out_wire_3_2(vertical_tile_13_21_to_tile_12_21_2),
		.out_wire_3_3(vertical_tile_13_21_to_tile_12_21_3),
		.in_wire_3_0(vertical_tile_12_21_to_tile_13_21_0),
		.in_wire_3_1(vertical_tile_12_21_to_tile_13_21_1),
		.in_wire_3_2(vertical_tile_12_21_to_tile_13_21_2),
		.in_wire_3_3(vertical_tile_12_21_to_tile_13_21_3),
		.out_wire_1_0(vertical_tile_13_21_to_tile_14_21_0),
		.out_wire_1_1(vertical_tile_13_21_to_tile_14_21_1),
		.out_wire_1_2(vertical_tile_13_21_to_tile_14_21_2),
		.out_wire_1_3(vertical_tile_13_21_to_tile_14_21_3),
		.in_wire_1_0(vertical_tile_14_21_to_tile_13_21_0),
		.in_wire_1_1(vertical_tile_14_21_to_tile_13_21_1),
		.in_wire_1_2(vertical_tile_14_21_to_tile_13_21_2),
		.in_wire_1_3(vertical_tile_14_21_to_tile_13_21_3),
		.out_wire_2_0(horizontal_tile_13_21_to_tile_13_20_0),
		.out_wire_2_1(horizontal_tile_13_21_to_tile_13_20_1),
		.out_wire_2_2(horizontal_tile_13_21_to_tile_13_20_2),
		.out_wire_2_3(horizontal_tile_13_21_to_tile_13_20_3),
		.in_wire_2_0(horizontal_tile_13_20_to_tile_13_21_0),
		.in_wire_2_1(horizontal_tile_13_20_to_tile_13_21_1),
		.in_wire_2_2(horizontal_tile_13_20_to_tile_13_21_2),
		.in_wire_2_3(horizontal_tile_13_20_to_tile_13_21_3),
		.out_wire_0_0(horizontal_tile_13_21_to_tile_13_22_0),
		.out_wire_0_1(horizontal_tile_13_21_to_tile_13_22_1),
		.out_wire_0_2(horizontal_tile_13_21_to_tile_13_22_2),
		.out_wire_0_3(horizontal_tile_13_21_to_tile_13_22_3),
		.in_wire_0_0(horizontal_tile_13_22_to_tile_13_21_0),
		.in_wire_0_1(horizontal_tile_13_22_to_tile_13_21_1),
		.in_wire_0_2(horizontal_tile_13_22_to_tile_13_21_2),
		.in_wire_0_3(horizontal_tile_13_22_to_tile_13_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(438)
	);

	pe_tile pe_tile_13_22(
		.out_wire_3_0(vertical_tile_13_22_to_tile_12_22_0),
		.out_wire_3_1(vertical_tile_13_22_to_tile_12_22_1),
		.out_wire_3_2(vertical_tile_13_22_to_tile_12_22_2),
		.out_wire_3_3(vertical_tile_13_22_to_tile_12_22_3),
		.in_wire_3_0(vertical_tile_12_22_to_tile_13_22_0),
		.in_wire_3_1(vertical_tile_12_22_to_tile_13_22_1),
		.in_wire_3_2(vertical_tile_12_22_to_tile_13_22_2),
		.in_wire_3_3(vertical_tile_12_22_to_tile_13_22_3),
		.out_wire_1_0(vertical_tile_13_22_to_tile_14_22_0),
		.out_wire_1_1(vertical_tile_13_22_to_tile_14_22_1),
		.out_wire_1_2(vertical_tile_13_22_to_tile_14_22_2),
		.out_wire_1_3(vertical_tile_13_22_to_tile_14_22_3),
		.in_wire_1_0(vertical_tile_14_22_to_tile_13_22_0),
		.in_wire_1_1(vertical_tile_14_22_to_tile_13_22_1),
		.in_wire_1_2(vertical_tile_14_22_to_tile_13_22_2),
		.in_wire_1_3(vertical_tile_14_22_to_tile_13_22_3),
		.out_wire_2_0(horizontal_tile_13_22_to_tile_13_21_0),
		.out_wire_2_1(horizontal_tile_13_22_to_tile_13_21_1),
		.out_wire_2_2(horizontal_tile_13_22_to_tile_13_21_2),
		.out_wire_2_3(horizontal_tile_13_22_to_tile_13_21_3),
		.in_wire_2_0(horizontal_tile_13_21_to_tile_13_22_0),
		.in_wire_2_1(horizontal_tile_13_21_to_tile_13_22_1),
		.in_wire_2_2(horizontal_tile_13_21_to_tile_13_22_2),
		.in_wire_2_3(horizontal_tile_13_21_to_tile_13_22_3),
		.out_wire_0_0(horizontal_tile_13_22_to_tile_13_23_0),
		.out_wire_0_1(horizontal_tile_13_22_to_tile_13_23_1),
		.out_wire_0_2(horizontal_tile_13_22_to_tile_13_23_2),
		.out_wire_0_3(horizontal_tile_13_22_to_tile_13_23_3),
		.in_wire_0_0(horizontal_tile_13_23_to_tile_13_22_0),
		.in_wire_0_1(horizontal_tile_13_23_to_tile_13_22_1),
		.in_wire_0_2(horizontal_tile_13_23_to_tile_13_22_2),
		.in_wire_0_3(horizontal_tile_13_23_to_tile_13_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(439)
	);

	pe_tile pe_tile_13_23(
		.out_wire_3_0(vertical_tile_13_23_to_tile_12_23_0),
		.out_wire_3_1(vertical_tile_13_23_to_tile_12_23_1),
		.out_wire_3_2(vertical_tile_13_23_to_tile_12_23_2),
		.out_wire_3_3(vertical_tile_13_23_to_tile_12_23_3),
		.in_wire_3_0(vertical_tile_12_23_to_tile_13_23_0),
		.in_wire_3_1(vertical_tile_12_23_to_tile_13_23_1),
		.in_wire_3_2(vertical_tile_12_23_to_tile_13_23_2),
		.in_wire_3_3(vertical_tile_12_23_to_tile_13_23_3),
		.out_wire_1_0(vertical_tile_13_23_to_tile_14_23_0),
		.out_wire_1_1(vertical_tile_13_23_to_tile_14_23_1),
		.out_wire_1_2(vertical_tile_13_23_to_tile_14_23_2),
		.out_wire_1_3(vertical_tile_13_23_to_tile_14_23_3),
		.in_wire_1_0(vertical_tile_14_23_to_tile_13_23_0),
		.in_wire_1_1(vertical_tile_14_23_to_tile_13_23_1),
		.in_wire_1_2(vertical_tile_14_23_to_tile_13_23_2),
		.in_wire_1_3(vertical_tile_14_23_to_tile_13_23_3),
		.out_wire_2_0(horizontal_tile_13_23_to_tile_13_22_0),
		.out_wire_2_1(horizontal_tile_13_23_to_tile_13_22_1),
		.out_wire_2_2(horizontal_tile_13_23_to_tile_13_22_2),
		.out_wire_2_3(horizontal_tile_13_23_to_tile_13_22_3),
		.in_wire_2_0(horizontal_tile_13_22_to_tile_13_23_0),
		.in_wire_2_1(horizontal_tile_13_22_to_tile_13_23_1),
		.in_wire_2_2(horizontal_tile_13_22_to_tile_13_23_2),
		.in_wire_2_3(horizontal_tile_13_22_to_tile_13_23_3),
		.out_wire_0_0(horizontal_tile_13_23_to_tile_13_24_0),
		.out_wire_0_1(horizontal_tile_13_23_to_tile_13_24_1),
		.out_wire_0_2(horizontal_tile_13_23_to_tile_13_24_2),
		.out_wire_0_3(horizontal_tile_13_23_to_tile_13_24_3),
		.in_wire_0_0(horizontal_tile_13_24_to_tile_13_23_0),
		.in_wire_0_1(horizontal_tile_13_24_to_tile_13_23_1),
		.in_wire_0_2(horizontal_tile_13_24_to_tile_13_23_2),
		.in_wire_0_3(horizontal_tile_13_24_to_tile_13_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(440)
	);

	pe_tile pe_tile_13_24(
		.out_wire_3_0(vertical_tile_13_24_to_tile_12_24_0),
		.out_wire_3_1(vertical_tile_13_24_to_tile_12_24_1),
		.out_wire_3_2(vertical_tile_13_24_to_tile_12_24_2),
		.out_wire_3_3(vertical_tile_13_24_to_tile_12_24_3),
		.in_wire_3_0(vertical_tile_12_24_to_tile_13_24_0),
		.in_wire_3_1(vertical_tile_12_24_to_tile_13_24_1),
		.in_wire_3_2(vertical_tile_12_24_to_tile_13_24_2),
		.in_wire_3_3(vertical_tile_12_24_to_tile_13_24_3),
		.out_wire_1_0(vertical_tile_13_24_to_tile_14_24_0),
		.out_wire_1_1(vertical_tile_13_24_to_tile_14_24_1),
		.out_wire_1_2(vertical_tile_13_24_to_tile_14_24_2),
		.out_wire_1_3(vertical_tile_13_24_to_tile_14_24_3),
		.in_wire_1_0(vertical_tile_14_24_to_tile_13_24_0),
		.in_wire_1_1(vertical_tile_14_24_to_tile_13_24_1),
		.in_wire_1_2(vertical_tile_14_24_to_tile_13_24_2),
		.in_wire_1_3(vertical_tile_14_24_to_tile_13_24_3),
		.out_wire_2_0(horizontal_tile_13_24_to_tile_13_23_0),
		.out_wire_2_1(horizontal_tile_13_24_to_tile_13_23_1),
		.out_wire_2_2(horizontal_tile_13_24_to_tile_13_23_2),
		.out_wire_2_3(horizontal_tile_13_24_to_tile_13_23_3),
		.in_wire_2_0(horizontal_tile_13_23_to_tile_13_24_0),
		.in_wire_2_1(horizontal_tile_13_23_to_tile_13_24_1),
		.in_wire_2_2(horizontal_tile_13_23_to_tile_13_24_2),
		.in_wire_2_3(horizontal_tile_13_23_to_tile_13_24_3),
		.out_wire_0_0(horizontal_tile_13_24_to_tile_13_25_0),
		.out_wire_0_1(horizontal_tile_13_24_to_tile_13_25_1),
		.out_wire_0_2(horizontal_tile_13_24_to_tile_13_25_2),
		.out_wire_0_3(horizontal_tile_13_24_to_tile_13_25_3),
		.in_wire_0_0(horizontal_tile_13_25_to_tile_13_24_0),
		.in_wire_0_1(horizontal_tile_13_25_to_tile_13_24_1),
		.in_wire_0_2(horizontal_tile_13_25_to_tile_13_24_2),
		.in_wire_0_3(horizontal_tile_13_25_to_tile_13_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(441)
	);

	pe_tile pe_tile_13_25(
		.out_wire_3_0(vertical_tile_13_25_to_tile_12_25_0),
		.out_wire_3_1(vertical_tile_13_25_to_tile_12_25_1),
		.out_wire_3_2(vertical_tile_13_25_to_tile_12_25_2),
		.out_wire_3_3(vertical_tile_13_25_to_tile_12_25_3),
		.in_wire_3_0(vertical_tile_12_25_to_tile_13_25_0),
		.in_wire_3_1(vertical_tile_12_25_to_tile_13_25_1),
		.in_wire_3_2(vertical_tile_12_25_to_tile_13_25_2),
		.in_wire_3_3(vertical_tile_12_25_to_tile_13_25_3),
		.out_wire_1_0(vertical_tile_13_25_to_tile_14_25_0),
		.out_wire_1_1(vertical_tile_13_25_to_tile_14_25_1),
		.out_wire_1_2(vertical_tile_13_25_to_tile_14_25_2),
		.out_wire_1_3(vertical_tile_13_25_to_tile_14_25_3),
		.in_wire_1_0(vertical_tile_14_25_to_tile_13_25_0),
		.in_wire_1_1(vertical_tile_14_25_to_tile_13_25_1),
		.in_wire_1_2(vertical_tile_14_25_to_tile_13_25_2),
		.in_wire_1_3(vertical_tile_14_25_to_tile_13_25_3),
		.out_wire_2_0(horizontal_tile_13_25_to_tile_13_24_0),
		.out_wire_2_1(horizontal_tile_13_25_to_tile_13_24_1),
		.out_wire_2_2(horizontal_tile_13_25_to_tile_13_24_2),
		.out_wire_2_3(horizontal_tile_13_25_to_tile_13_24_3),
		.in_wire_2_0(horizontal_tile_13_24_to_tile_13_25_0),
		.in_wire_2_1(horizontal_tile_13_24_to_tile_13_25_1),
		.in_wire_2_2(horizontal_tile_13_24_to_tile_13_25_2),
		.in_wire_2_3(horizontal_tile_13_24_to_tile_13_25_3),
		.out_wire_0_0(horizontal_tile_13_25_to_tile_13_26_0),
		.out_wire_0_1(horizontal_tile_13_25_to_tile_13_26_1),
		.out_wire_0_2(horizontal_tile_13_25_to_tile_13_26_2),
		.out_wire_0_3(horizontal_tile_13_25_to_tile_13_26_3),
		.in_wire_0_0(horizontal_tile_13_26_to_tile_13_25_0),
		.in_wire_0_1(horizontal_tile_13_26_to_tile_13_25_1),
		.in_wire_0_2(horizontal_tile_13_26_to_tile_13_25_2),
		.in_wire_0_3(horizontal_tile_13_26_to_tile_13_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(442)
	);

	pe_tile pe_tile_13_26(
		.out_wire_3_0(vertical_tile_13_26_to_tile_12_26_0),
		.out_wire_3_1(vertical_tile_13_26_to_tile_12_26_1),
		.out_wire_3_2(vertical_tile_13_26_to_tile_12_26_2),
		.out_wire_3_3(vertical_tile_13_26_to_tile_12_26_3),
		.in_wire_3_0(vertical_tile_12_26_to_tile_13_26_0),
		.in_wire_3_1(vertical_tile_12_26_to_tile_13_26_1),
		.in_wire_3_2(vertical_tile_12_26_to_tile_13_26_2),
		.in_wire_3_3(vertical_tile_12_26_to_tile_13_26_3),
		.out_wire_1_0(vertical_tile_13_26_to_tile_14_26_0),
		.out_wire_1_1(vertical_tile_13_26_to_tile_14_26_1),
		.out_wire_1_2(vertical_tile_13_26_to_tile_14_26_2),
		.out_wire_1_3(vertical_tile_13_26_to_tile_14_26_3),
		.in_wire_1_0(vertical_tile_14_26_to_tile_13_26_0),
		.in_wire_1_1(vertical_tile_14_26_to_tile_13_26_1),
		.in_wire_1_2(vertical_tile_14_26_to_tile_13_26_2),
		.in_wire_1_3(vertical_tile_14_26_to_tile_13_26_3),
		.out_wire_2_0(horizontal_tile_13_26_to_tile_13_25_0),
		.out_wire_2_1(horizontal_tile_13_26_to_tile_13_25_1),
		.out_wire_2_2(horizontal_tile_13_26_to_tile_13_25_2),
		.out_wire_2_3(horizontal_tile_13_26_to_tile_13_25_3),
		.in_wire_2_0(horizontal_tile_13_25_to_tile_13_26_0),
		.in_wire_2_1(horizontal_tile_13_25_to_tile_13_26_1),
		.in_wire_2_2(horizontal_tile_13_25_to_tile_13_26_2),
		.in_wire_2_3(horizontal_tile_13_25_to_tile_13_26_3),
		.out_wire_0_0(horizontal_tile_13_26_to_tile_13_27_0),
		.out_wire_0_1(horizontal_tile_13_26_to_tile_13_27_1),
		.out_wire_0_2(horizontal_tile_13_26_to_tile_13_27_2),
		.out_wire_0_3(horizontal_tile_13_26_to_tile_13_27_3),
		.in_wire_0_0(horizontal_tile_13_27_to_tile_13_26_0),
		.in_wire_0_1(horizontal_tile_13_27_to_tile_13_26_1),
		.in_wire_0_2(horizontal_tile_13_27_to_tile_13_26_2),
		.in_wire_0_3(horizontal_tile_13_27_to_tile_13_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(443)
	);

	pe_tile pe_tile_13_27(
		.out_wire_3_0(vertical_tile_13_27_to_tile_12_27_0),
		.out_wire_3_1(vertical_tile_13_27_to_tile_12_27_1),
		.out_wire_3_2(vertical_tile_13_27_to_tile_12_27_2),
		.out_wire_3_3(vertical_tile_13_27_to_tile_12_27_3),
		.in_wire_3_0(vertical_tile_12_27_to_tile_13_27_0),
		.in_wire_3_1(vertical_tile_12_27_to_tile_13_27_1),
		.in_wire_3_2(vertical_tile_12_27_to_tile_13_27_2),
		.in_wire_3_3(vertical_tile_12_27_to_tile_13_27_3),
		.out_wire_1_0(vertical_tile_13_27_to_tile_14_27_0),
		.out_wire_1_1(vertical_tile_13_27_to_tile_14_27_1),
		.out_wire_1_2(vertical_tile_13_27_to_tile_14_27_2),
		.out_wire_1_3(vertical_tile_13_27_to_tile_14_27_3),
		.in_wire_1_0(vertical_tile_14_27_to_tile_13_27_0),
		.in_wire_1_1(vertical_tile_14_27_to_tile_13_27_1),
		.in_wire_1_2(vertical_tile_14_27_to_tile_13_27_2),
		.in_wire_1_3(vertical_tile_14_27_to_tile_13_27_3),
		.out_wire_2_0(horizontal_tile_13_27_to_tile_13_26_0),
		.out_wire_2_1(horizontal_tile_13_27_to_tile_13_26_1),
		.out_wire_2_2(horizontal_tile_13_27_to_tile_13_26_2),
		.out_wire_2_3(horizontal_tile_13_27_to_tile_13_26_3),
		.in_wire_2_0(horizontal_tile_13_26_to_tile_13_27_0),
		.in_wire_2_1(horizontal_tile_13_26_to_tile_13_27_1),
		.in_wire_2_2(horizontal_tile_13_26_to_tile_13_27_2),
		.in_wire_2_3(horizontal_tile_13_26_to_tile_13_27_3),
		.out_wire_0_0(horizontal_tile_13_27_to_tile_13_28_0),
		.out_wire_0_1(horizontal_tile_13_27_to_tile_13_28_1),
		.out_wire_0_2(horizontal_tile_13_27_to_tile_13_28_2),
		.out_wire_0_3(horizontal_tile_13_27_to_tile_13_28_3),
		.in_wire_0_0(horizontal_tile_13_28_to_tile_13_27_0),
		.in_wire_0_1(horizontal_tile_13_28_to_tile_13_27_1),
		.in_wire_0_2(horizontal_tile_13_28_to_tile_13_27_2),
		.in_wire_0_3(horizontal_tile_13_28_to_tile_13_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(444)
	);

	pe_tile pe_tile_13_28(
		.out_wire_3_0(vertical_tile_13_28_to_tile_12_28_0),
		.out_wire_3_1(vertical_tile_13_28_to_tile_12_28_1),
		.out_wire_3_2(vertical_tile_13_28_to_tile_12_28_2),
		.out_wire_3_3(vertical_tile_13_28_to_tile_12_28_3),
		.in_wire_3_0(vertical_tile_12_28_to_tile_13_28_0),
		.in_wire_3_1(vertical_tile_12_28_to_tile_13_28_1),
		.in_wire_3_2(vertical_tile_12_28_to_tile_13_28_2),
		.in_wire_3_3(vertical_tile_12_28_to_tile_13_28_3),
		.out_wire_1_0(vertical_tile_13_28_to_tile_14_28_0),
		.out_wire_1_1(vertical_tile_13_28_to_tile_14_28_1),
		.out_wire_1_2(vertical_tile_13_28_to_tile_14_28_2),
		.out_wire_1_3(vertical_tile_13_28_to_tile_14_28_3),
		.in_wire_1_0(vertical_tile_14_28_to_tile_13_28_0),
		.in_wire_1_1(vertical_tile_14_28_to_tile_13_28_1),
		.in_wire_1_2(vertical_tile_14_28_to_tile_13_28_2),
		.in_wire_1_3(vertical_tile_14_28_to_tile_13_28_3),
		.out_wire_2_0(horizontal_tile_13_28_to_tile_13_27_0),
		.out_wire_2_1(horizontal_tile_13_28_to_tile_13_27_1),
		.out_wire_2_2(horizontal_tile_13_28_to_tile_13_27_2),
		.out_wire_2_3(horizontal_tile_13_28_to_tile_13_27_3),
		.in_wire_2_0(horizontal_tile_13_27_to_tile_13_28_0),
		.in_wire_2_1(horizontal_tile_13_27_to_tile_13_28_1),
		.in_wire_2_2(horizontal_tile_13_27_to_tile_13_28_2),
		.in_wire_2_3(horizontal_tile_13_27_to_tile_13_28_3),
		.out_wire_0_0(horizontal_tile_13_28_to_tile_13_29_0),
		.out_wire_0_1(horizontal_tile_13_28_to_tile_13_29_1),
		.out_wire_0_2(horizontal_tile_13_28_to_tile_13_29_2),
		.out_wire_0_3(horizontal_tile_13_28_to_tile_13_29_3),
		.in_wire_0_0(horizontal_tile_13_29_to_tile_13_28_0),
		.in_wire_0_1(horizontal_tile_13_29_to_tile_13_28_1),
		.in_wire_0_2(horizontal_tile_13_29_to_tile_13_28_2),
		.in_wire_0_3(horizontal_tile_13_29_to_tile_13_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(445)
	);

	pe_tile pe_tile_13_29(
		.out_wire_3_0(vertical_tile_13_29_to_tile_12_29_0),
		.out_wire_3_1(vertical_tile_13_29_to_tile_12_29_1),
		.out_wire_3_2(vertical_tile_13_29_to_tile_12_29_2),
		.out_wire_3_3(vertical_tile_13_29_to_tile_12_29_3),
		.in_wire_3_0(vertical_tile_12_29_to_tile_13_29_0),
		.in_wire_3_1(vertical_tile_12_29_to_tile_13_29_1),
		.in_wire_3_2(vertical_tile_12_29_to_tile_13_29_2),
		.in_wire_3_3(vertical_tile_12_29_to_tile_13_29_3),
		.out_wire_1_0(vertical_tile_13_29_to_tile_14_29_0),
		.out_wire_1_1(vertical_tile_13_29_to_tile_14_29_1),
		.out_wire_1_2(vertical_tile_13_29_to_tile_14_29_2),
		.out_wire_1_3(vertical_tile_13_29_to_tile_14_29_3),
		.in_wire_1_0(vertical_tile_14_29_to_tile_13_29_0),
		.in_wire_1_1(vertical_tile_14_29_to_tile_13_29_1),
		.in_wire_1_2(vertical_tile_14_29_to_tile_13_29_2),
		.in_wire_1_3(vertical_tile_14_29_to_tile_13_29_3),
		.out_wire_2_0(horizontal_tile_13_29_to_tile_13_28_0),
		.out_wire_2_1(horizontal_tile_13_29_to_tile_13_28_1),
		.out_wire_2_2(horizontal_tile_13_29_to_tile_13_28_2),
		.out_wire_2_3(horizontal_tile_13_29_to_tile_13_28_3),
		.in_wire_2_0(horizontal_tile_13_28_to_tile_13_29_0),
		.in_wire_2_1(horizontal_tile_13_28_to_tile_13_29_1),
		.in_wire_2_2(horizontal_tile_13_28_to_tile_13_29_2),
		.in_wire_2_3(horizontal_tile_13_28_to_tile_13_29_3),
		.out_wire_0_0(horizontal_tile_13_29_to_tile_13_30_0),
		.out_wire_0_1(horizontal_tile_13_29_to_tile_13_30_1),
		.out_wire_0_2(horizontal_tile_13_29_to_tile_13_30_2),
		.out_wire_0_3(horizontal_tile_13_29_to_tile_13_30_3),
		.in_wire_0_0(horizontal_tile_13_30_to_tile_13_29_0),
		.in_wire_0_1(horizontal_tile_13_30_to_tile_13_29_1),
		.in_wire_0_2(horizontal_tile_13_30_to_tile_13_29_2),
		.in_wire_0_3(horizontal_tile_13_30_to_tile_13_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(446)
	);

	pe_tile pe_tile_13_30(
		.out_wire_3_0(vertical_tile_13_30_to_tile_12_30_0),
		.out_wire_3_1(vertical_tile_13_30_to_tile_12_30_1),
		.out_wire_3_2(vertical_tile_13_30_to_tile_12_30_2),
		.out_wire_3_3(vertical_tile_13_30_to_tile_12_30_3),
		.in_wire_3_0(vertical_tile_12_30_to_tile_13_30_0),
		.in_wire_3_1(vertical_tile_12_30_to_tile_13_30_1),
		.in_wire_3_2(vertical_tile_12_30_to_tile_13_30_2),
		.in_wire_3_3(vertical_tile_12_30_to_tile_13_30_3),
		.out_wire_1_0(vertical_tile_13_30_to_tile_14_30_0),
		.out_wire_1_1(vertical_tile_13_30_to_tile_14_30_1),
		.out_wire_1_2(vertical_tile_13_30_to_tile_14_30_2),
		.out_wire_1_3(vertical_tile_13_30_to_tile_14_30_3),
		.in_wire_1_0(vertical_tile_14_30_to_tile_13_30_0),
		.in_wire_1_1(vertical_tile_14_30_to_tile_13_30_1),
		.in_wire_1_2(vertical_tile_14_30_to_tile_13_30_2),
		.in_wire_1_3(vertical_tile_14_30_to_tile_13_30_3),
		.out_wire_2_0(horizontal_tile_13_30_to_tile_13_29_0),
		.out_wire_2_1(horizontal_tile_13_30_to_tile_13_29_1),
		.out_wire_2_2(horizontal_tile_13_30_to_tile_13_29_2),
		.out_wire_2_3(horizontal_tile_13_30_to_tile_13_29_3),
		.in_wire_2_0(horizontal_tile_13_29_to_tile_13_30_0),
		.in_wire_2_1(horizontal_tile_13_29_to_tile_13_30_1),
		.in_wire_2_2(horizontal_tile_13_29_to_tile_13_30_2),
		.in_wire_2_3(horizontal_tile_13_29_to_tile_13_30_3),
		.out_wire_0_0(horizontal_tile_13_30_to_tile_13_31_0),
		.out_wire_0_1(horizontal_tile_13_30_to_tile_13_31_1),
		.out_wire_0_2(horizontal_tile_13_30_to_tile_13_31_2),
		.out_wire_0_3(horizontal_tile_13_30_to_tile_13_31_3),
		.in_wire_0_0(horizontal_tile_13_31_to_tile_13_30_0),
		.in_wire_0_1(horizontal_tile_13_31_to_tile_13_30_1),
		.in_wire_0_2(horizontal_tile_13_31_to_tile_13_30_2),
		.in_wire_0_3(horizontal_tile_13_31_to_tile_13_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(447)
	);

	pe_tile_right pe_tile_13_31(
		.out_wire_3_0(vertical_tile_13_31_to_tile_12_31_0),
		.out_wire_3_1(vertical_tile_13_31_to_tile_12_31_1),
		.out_wire_3_2(vertical_tile_13_31_to_tile_12_31_2),
		.out_wire_3_3(vertical_tile_13_31_to_tile_12_31_3),
		.in_wire_3_0(vertical_tile_12_31_to_tile_13_31_0),
		.in_wire_3_1(vertical_tile_12_31_to_tile_13_31_1),
		.in_wire_3_2(vertical_tile_12_31_to_tile_13_31_2),
		.in_wire_3_3(vertical_tile_12_31_to_tile_13_31_3),
		.out_wire_1_0(vertical_tile_13_31_to_tile_14_31_0),
		.out_wire_1_1(vertical_tile_13_31_to_tile_14_31_1),
		.out_wire_1_2(vertical_tile_13_31_to_tile_14_31_2),
		.out_wire_1_3(vertical_tile_13_31_to_tile_14_31_3),
		.in_wire_1_0(vertical_tile_14_31_to_tile_13_31_0),
		.in_wire_1_1(vertical_tile_14_31_to_tile_13_31_1),
		.in_wire_1_2(vertical_tile_14_31_to_tile_13_31_2),
		.in_wire_1_3(vertical_tile_14_31_to_tile_13_31_3),
		.out_wire_2_0(horizontal_tile_13_31_to_tile_13_30_0),
		.out_wire_2_1(horizontal_tile_13_31_to_tile_13_30_1),
		.out_wire_2_2(horizontal_tile_13_31_to_tile_13_30_2),
		.out_wire_2_3(horizontal_tile_13_31_to_tile_13_30_3),
		.in_wire_2_0(horizontal_tile_13_30_to_tile_13_31_0),
		.in_wire_2_1(horizontal_tile_13_30_to_tile_13_31_1),
		.in_wire_2_2(horizontal_tile_13_30_to_tile_13_31_2),
		.in_wire_2_3(horizontal_tile_13_30_to_tile_13_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(448)
	);

	pe_tile_left pe_tile_14_0(
		.out_wire_3_0(vertical_tile_14_0_to_tile_13_0_0),
		.out_wire_3_1(vertical_tile_14_0_to_tile_13_0_1),
		.out_wire_3_2(vertical_tile_14_0_to_tile_13_0_2),
		.out_wire_3_3(vertical_tile_14_0_to_tile_13_0_3),
		.in_wire_3_0(vertical_tile_13_0_to_tile_14_0_0),
		.in_wire_3_1(vertical_tile_13_0_to_tile_14_0_1),
		.in_wire_3_2(vertical_tile_13_0_to_tile_14_0_2),
		.in_wire_3_3(vertical_tile_13_0_to_tile_14_0_3),
		.out_wire_1_0(vertical_tile_14_0_to_tile_15_0_0),
		.out_wire_1_1(vertical_tile_14_0_to_tile_15_0_1),
		.out_wire_1_2(vertical_tile_14_0_to_tile_15_0_2),
		.out_wire_1_3(vertical_tile_14_0_to_tile_15_0_3),
		.in_wire_1_0(vertical_tile_15_0_to_tile_14_0_0),
		.in_wire_1_1(vertical_tile_15_0_to_tile_14_0_1),
		.in_wire_1_2(vertical_tile_15_0_to_tile_14_0_2),
		.in_wire_1_3(vertical_tile_15_0_to_tile_14_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_14_0_to_tile_14_1_0),
		.out_wire_0_1(horizontal_tile_14_0_to_tile_14_1_1),
		.out_wire_0_2(horizontal_tile_14_0_to_tile_14_1_2),
		.out_wire_0_3(horizontal_tile_14_0_to_tile_14_1_3),
		.in_wire_0_0(horizontal_tile_14_1_to_tile_14_0_0),
		.in_wire_0_1(horizontal_tile_14_1_to_tile_14_0_1),
		.in_wire_0_2(horizontal_tile_14_1_to_tile_14_0_2),
		.in_wire_0_3(horizontal_tile_14_1_to_tile_14_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(449)
	);

	pe_tile pe_tile_14_1(
		.out_wire_3_0(vertical_tile_14_1_to_tile_13_1_0),
		.out_wire_3_1(vertical_tile_14_1_to_tile_13_1_1),
		.out_wire_3_2(vertical_tile_14_1_to_tile_13_1_2),
		.out_wire_3_3(vertical_tile_14_1_to_tile_13_1_3),
		.in_wire_3_0(vertical_tile_13_1_to_tile_14_1_0),
		.in_wire_3_1(vertical_tile_13_1_to_tile_14_1_1),
		.in_wire_3_2(vertical_tile_13_1_to_tile_14_1_2),
		.in_wire_3_3(vertical_tile_13_1_to_tile_14_1_3),
		.out_wire_1_0(vertical_tile_14_1_to_tile_15_1_0),
		.out_wire_1_1(vertical_tile_14_1_to_tile_15_1_1),
		.out_wire_1_2(vertical_tile_14_1_to_tile_15_1_2),
		.out_wire_1_3(vertical_tile_14_1_to_tile_15_1_3),
		.in_wire_1_0(vertical_tile_15_1_to_tile_14_1_0),
		.in_wire_1_1(vertical_tile_15_1_to_tile_14_1_1),
		.in_wire_1_2(vertical_tile_15_1_to_tile_14_1_2),
		.in_wire_1_3(vertical_tile_15_1_to_tile_14_1_3),
		.out_wire_2_0(horizontal_tile_14_1_to_tile_14_0_0),
		.out_wire_2_1(horizontal_tile_14_1_to_tile_14_0_1),
		.out_wire_2_2(horizontal_tile_14_1_to_tile_14_0_2),
		.out_wire_2_3(horizontal_tile_14_1_to_tile_14_0_3),
		.in_wire_2_0(horizontal_tile_14_0_to_tile_14_1_0),
		.in_wire_2_1(horizontal_tile_14_0_to_tile_14_1_1),
		.in_wire_2_2(horizontal_tile_14_0_to_tile_14_1_2),
		.in_wire_2_3(horizontal_tile_14_0_to_tile_14_1_3),
		.out_wire_0_0(horizontal_tile_14_1_to_tile_14_2_0),
		.out_wire_0_1(horizontal_tile_14_1_to_tile_14_2_1),
		.out_wire_0_2(horizontal_tile_14_1_to_tile_14_2_2),
		.out_wire_0_3(horizontal_tile_14_1_to_tile_14_2_3),
		.in_wire_0_0(horizontal_tile_14_2_to_tile_14_1_0),
		.in_wire_0_1(horizontal_tile_14_2_to_tile_14_1_1),
		.in_wire_0_2(horizontal_tile_14_2_to_tile_14_1_2),
		.in_wire_0_3(horizontal_tile_14_2_to_tile_14_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(450)
	);

	pe_tile pe_tile_14_2(
		.out_wire_3_0(vertical_tile_14_2_to_tile_13_2_0),
		.out_wire_3_1(vertical_tile_14_2_to_tile_13_2_1),
		.out_wire_3_2(vertical_tile_14_2_to_tile_13_2_2),
		.out_wire_3_3(vertical_tile_14_2_to_tile_13_2_3),
		.in_wire_3_0(vertical_tile_13_2_to_tile_14_2_0),
		.in_wire_3_1(vertical_tile_13_2_to_tile_14_2_1),
		.in_wire_3_2(vertical_tile_13_2_to_tile_14_2_2),
		.in_wire_3_3(vertical_tile_13_2_to_tile_14_2_3),
		.out_wire_1_0(vertical_tile_14_2_to_tile_15_2_0),
		.out_wire_1_1(vertical_tile_14_2_to_tile_15_2_1),
		.out_wire_1_2(vertical_tile_14_2_to_tile_15_2_2),
		.out_wire_1_3(vertical_tile_14_2_to_tile_15_2_3),
		.in_wire_1_0(vertical_tile_15_2_to_tile_14_2_0),
		.in_wire_1_1(vertical_tile_15_2_to_tile_14_2_1),
		.in_wire_1_2(vertical_tile_15_2_to_tile_14_2_2),
		.in_wire_1_3(vertical_tile_15_2_to_tile_14_2_3),
		.out_wire_2_0(horizontal_tile_14_2_to_tile_14_1_0),
		.out_wire_2_1(horizontal_tile_14_2_to_tile_14_1_1),
		.out_wire_2_2(horizontal_tile_14_2_to_tile_14_1_2),
		.out_wire_2_3(horizontal_tile_14_2_to_tile_14_1_3),
		.in_wire_2_0(horizontal_tile_14_1_to_tile_14_2_0),
		.in_wire_2_1(horizontal_tile_14_1_to_tile_14_2_1),
		.in_wire_2_2(horizontal_tile_14_1_to_tile_14_2_2),
		.in_wire_2_3(horizontal_tile_14_1_to_tile_14_2_3),
		.out_wire_0_0(horizontal_tile_14_2_to_tile_14_3_0),
		.out_wire_0_1(horizontal_tile_14_2_to_tile_14_3_1),
		.out_wire_0_2(horizontal_tile_14_2_to_tile_14_3_2),
		.out_wire_0_3(horizontal_tile_14_2_to_tile_14_3_3),
		.in_wire_0_0(horizontal_tile_14_3_to_tile_14_2_0),
		.in_wire_0_1(horizontal_tile_14_3_to_tile_14_2_1),
		.in_wire_0_2(horizontal_tile_14_3_to_tile_14_2_2),
		.in_wire_0_3(horizontal_tile_14_3_to_tile_14_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(451)
	);

	pe_tile pe_tile_14_3(
		.out_wire_3_0(vertical_tile_14_3_to_tile_13_3_0),
		.out_wire_3_1(vertical_tile_14_3_to_tile_13_3_1),
		.out_wire_3_2(vertical_tile_14_3_to_tile_13_3_2),
		.out_wire_3_3(vertical_tile_14_3_to_tile_13_3_3),
		.in_wire_3_0(vertical_tile_13_3_to_tile_14_3_0),
		.in_wire_3_1(vertical_tile_13_3_to_tile_14_3_1),
		.in_wire_3_2(vertical_tile_13_3_to_tile_14_3_2),
		.in_wire_3_3(vertical_tile_13_3_to_tile_14_3_3),
		.out_wire_1_0(vertical_tile_14_3_to_tile_15_3_0),
		.out_wire_1_1(vertical_tile_14_3_to_tile_15_3_1),
		.out_wire_1_2(vertical_tile_14_3_to_tile_15_3_2),
		.out_wire_1_3(vertical_tile_14_3_to_tile_15_3_3),
		.in_wire_1_0(vertical_tile_15_3_to_tile_14_3_0),
		.in_wire_1_1(vertical_tile_15_3_to_tile_14_3_1),
		.in_wire_1_2(vertical_tile_15_3_to_tile_14_3_2),
		.in_wire_1_3(vertical_tile_15_3_to_tile_14_3_3),
		.out_wire_2_0(horizontal_tile_14_3_to_tile_14_2_0),
		.out_wire_2_1(horizontal_tile_14_3_to_tile_14_2_1),
		.out_wire_2_2(horizontal_tile_14_3_to_tile_14_2_2),
		.out_wire_2_3(horizontal_tile_14_3_to_tile_14_2_3),
		.in_wire_2_0(horizontal_tile_14_2_to_tile_14_3_0),
		.in_wire_2_1(horizontal_tile_14_2_to_tile_14_3_1),
		.in_wire_2_2(horizontal_tile_14_2_to_tile_14_3_2),
		.in_wire_2_3(horizontal_tile_14_2_to_tile_14_3_3),
		.out_wire_0_0(horizontal_tile_14_3_to_tile_14_4_0),
		.out_wire_0_1(horizontal_tile_14_3_to_tile_14_4_1),
		.out_wire_0_2(horizontal_tile_14_3_to_tile_14_4_2),
		.out_wire_0_3(horizontal_tile_14_3_to_tile_14_4_3),
		.in_wire_0_0(horizontal_tile_14_4_to_tile_14_3_0),
		.in_wire_0_1(horizontal_tile_14_4_to_tile_14_3_1),
		.in_wire_0_2(horizontal_tile_14_4_to_tile_14_3_2),
		.in_wire_0_3(horizontal_tile_14_4_to_tile_14_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(452)
	);

	pe_tile pe_tile_14_4(
		.out_wire_3_0(vertical_tile_14_4_to_tile_13_4_0),
		.out_wire_3_1(vertical_tile_14_4_to_tile_13_4_1),
		.out_wire_3_2(vertical_tile_14_4_to_tile_13_4_2),
		.out_wire_3_3(vertical_tile_14_4_to_tile_13_4_3),
		.in_wire_3_0(vertical_tile_13_4_to_tile_14_4_0),
		.in_wire_3_1(vertical_tile_13_4_to_tile_14_4_1),
		.in_wire_3_2(vertical_tile_13_4_to_tile_14_4_2),
		.in_wire_3_3(vertical_tile_13_4_to_tile_14_4_3),
		.out_wire_1_0(vertical_tile_14_4_to_tile_15_4_0),
		.out_wire_1_1(vertical_tile_14_4_to_tile_15_4_1),
		.out_wire_1_2(vertical_tile_14_4_to_tile_15_4_2),
		.out_wire_1_3(vertical_tile_14_4_to_tile_15_4_3),
		.in_wire_1_0(vertical_tile_15_4_to_tile_14_4_0),
		.in_wire_1_1(vertical_tile_15_4_to_tile_14_4_1),
		.in_wire_1_2(vertical_tile_15_4_to_tile_14_4_2),
		.in_wire_1_3(vertical_tile_15_4_to_tile_14_4_3),
		.out_wire_2_0(horizontal_tile_14_4_to_tile_14_3_0),
		.out_wire_2_1(horizontal_tile_14_4_to_tile_14_3_1),
		.out_wire_2_2(horizontal_tile_14_4_to_tile_14_3_2),
		.out_wire_2_3(horizontal_tile_14_4_to_tile_14_3_3),
		.in_wire_2_0(horizontal_tile_14_3_to_tile_14_4_0),
		.in_wire_2_1(horizontal_tile_14_3_to_tile_14_4_1),
		.in_wire_2_2(horizontal_tile_14_3_to_tile_14_4_2),
		.in_wire_2_3(horizontal_tile_14_3_to_tile_14_4_3),
		.out_wire_0_0(horizontal_tile_14_4_to_tile_14_5_0),
		.out_wire_0_1(horizontal_tile_14_4_to_tile_14_5_1),
		.out_wire_0_2(horizontal_tile_14_4_to_tile_14_5_2),
		.out_wire_0_3(horizontal_tile_14_4_to_tile_14_5_3),
		.in_wire_0_0(horizontal_tile_14_5_to_tile_14_4_0),
		.in_wire_0_1(horizontal_tile_14_5_to_tile_14_4_1),
		.in_wire_0_2(horizontal_tile_14_5_to_tile_14_4_2),
		.in_wire_0_3(horizontal_tile_14_5_to_tile_14_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(453)
	);

	pe_tile pe_tile_14_5(
		.out_wire_3_0(vertical_tile_14_5_to_tile_13_5_0),
		.out_wire_3_1(vertical_tile_14_5_to_tile_13_5_1),
		.out_wire_3_2(vertical_tile_14_5_to_tile_13_5_2),
		.out_wire_3_3(vertical_tile_14_5_to_tile_13_5_3),
		.in_wire_3_0(vertical_tile_13_5_to_tile_14_5_0),
		.in_wire_3_1(vertical_tile_13_5_to_tile_14_5_1),
		.in_wire_3_2(vertical_tile_13_5_to_tile_14_5_2),
		.in_wire_3_3(vertical_tile_13_5_to_tile_14_5_3),
		.out_wire_1_0(vertical_tile_14_5_to_tile_15_5_0),
		.out_wire_1_1(vertical_tile_14_5_to_tile_15_5_1),
		.out_wire_1_2(vertical_tile_14_5_to_tile_15_5_2),
		.out_wire_1_3(vertical_tile_14_5_to_tile_15_5_3),
		.in_wire_1_0(vertical_tile_15_5_to_tile_14_5_0),
		.in_wire_1_1(vertical_tile_15_5_to_tile_14_5_1),
		.in_wire_1_2(vertical_tile_15_5_to_tile_14_5_2),
		.in_wire_1_3(vertical_tile_15_5_to_tile_14_5_3),
		.out_wire_2_0(horizontal_tile_14_5_to_tile_14_4_0),
		.out_wire_2_1(horizontal_tile_14_5_to_tile_14_4_1),
		.out_wire_2_2(horizontal_tile_14_5_to_tile_14_4_2),
		.out_wire_2_3(horizontal_tile_14_5_to_tile_14_4_3),
		.in_wire_2_0(horizontal_tile_14_4_to_tile_14_5_0),
		.in_wire_2_1(horizontal_tile_14_4_to_tile_14_5_1),
		.in_wire_2_2(horizontal_tile_14_4_to_tile_14_5_2),
		.in_wire_2_3(horizontal_tile_14_4_to_tile_14_5_3),
		.out_wire_0_0(horizontal_tile_14_5_to_tile_14_6_0),
		.out_wire_0_1(horizontal_tile_14_5_to_tile_14_6_1),
		.out_wire_0_2(horizontal_tile_14_5_to_tile_14_6_2),
		.out_wire_0_3(horizontal_tile_14_5_to_tile_14_6_3),
		.in_wire_0_0(horizontal_tile_14_6_to_tile_14_5_0),
		.in_wire_0_1(horizontal_tile_14_6_to_tile_14_5_1),
		.in_wire_0_2(horizontal_tile_14_6_to_tile_14_5_2),
		.in_wire_0_3(horizontal_tile_14_6_to_tile_14_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(454)
	);

	pe_tile pe_tile_14_6(
		.out_wire_3_0(vertical_tile_14_6_to_tile_13_6_0),
		.out_wire_3_1(vertical_tile_14_6_to_tile_13_6_1),
		.out_wire_3_2(vertical_tile_14_6_to_tile_13_6_2),
		.out_wire_3_3(vertical_tile_14_6_to_tile_13_6_3),
		.in_wire_3_0(vertical_tile_13_6_to_tile_14_6_0),
		.in_wire_3_1(vertical_tile_13_6_to_tile_14_6_1),
		.in_wire_3_2(vertical_tile_13_6_to_tile_14_6_2),
		.in_wire_3_3(vertical_tile_13_6_to_tile_14_6_3),
		.out_wire_1_0(vertical_tile_14_6_to_tile_15_6_0),
		.out_wire_1_1(vertical_tile_14_6_to_tile_15_6_1),
		.out_wire_1_2(vertical_tile_14_6_to_tile_15_6_2),
		.out_wire_1_3(vertical_tile_14_6_to_tile_15_6_3),
		.in_wire_1_0(vertical_tile_15_6_to_tile_14_6_0),
		.in_wire_1_1(vertical_tile_15_6_to_tile_14_6_1),
		.in_wire_1_2(vertical_tile_15_6_to_tile_14_6_2),
		.in_wire_1_3(vertical_tile_15_6_to_tile_14_6_3),
		.out_wire_2_0(horizontal_tile_14_6_to_tile_14_5_0),
		.out_wire_2_1(horizontal_tile_14_6_to_tile_14_5_1),
		.out_wire_2_2(horizontal_tile_14_6_to_tile_14_5_2),
		.out_wire_2_3(horizontal_tile_14_6_to_tile_14_5_3),
		.in_wire_2_0(horizontal_tile_14_5_to_tile_14_6_0),
		.in_wire_2_1(horizontal_tile_14_5_to_tile_14_6_1),
		.in_wire_2_2(horizontal_tile_14_5_to_tile_14_6_2),
		.in_wire_2_3(horizontal_tile_14_5_to_tile_14_6_3),
		.out_wire_0_0(horizontal_tile_14_6_to_tile_14_7_0),
		.out_wire_0_1(horizontal_tile_14_6_to_tile_14_7_1),
		.out_wire_0_2(horizontal_tile_14_6_to_tile_14_7_2),
		.out_wire_0_3(horizontal_tile_14_6_to_tile_14_7_3),
		.in_wire_0_0(horizontal_tile_14_7_to_tile_14_6_0),
		.in_wire_0_1(horizontal_tile_14_7_to_tile_14_6_1),
		.in_wire_0_2(horizontal_tile_14_7_to_tile_14_6_2),
		.in_wire_0_3(horizontal_tile_14_7_to_tile_14_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(455)
	);

	pe_tile pe_tile_14_7(
		.out_wire_3_0(vertical_tile_14_7_to_tile_13_7_0),
		.out_wire_3_1(vertical_tile_14_7_to_tile_13_7_1),
		.out_wire_3_2(vertical_tile_14_7_to_tile_13_7_2),
		.out_wire_3_3(vertical_tile_14_7_to_tile_13_7_3),
		.in_wire_3_0(vertical_tile_13_7_to_tile_14_7_0),
		.in_wire_3_1(vertical_tile_13_7_to_tile_14_7_1),
		.in_wire_3_2(vertical_tile_13_7_to_tile_14_7_2),
		.in_wire_3_3(vertical_tile_13_7_to_tile_14_7_3),
		.out_wire_1_0(vertical_tile_14_7_to_tile_15_7_0),
		.out_wire_1_1(vertical_tile_14_7_to_tile_15_7_1),
		.out_wire_1_2(vertical_tile_14_7_to_tile_15_7_2),
		.out_wire_1_3(vertical_tile_14_7_to_tile_15_7_3),
		.in_wire_1_0(vertical_tile_15_7_to_tile_14_7_0),
		.in_wire_1_1(vertical_tile_15_7_to_tile_14_7_1),
		.in_wire_1_2(vertical_tile_15_7_to_tile_14_7_2),
		.in_wire_1_3(vertical_tile_15_7_to_tile_14_7_3),
		.out_wire_2_0(horizontal_tile_14_7_to_tile_14_6_0),
		.out_wire_2_1(horizontal_tile_14_7_to_tile_14_6_1),
		.out_wire_2_2(horizontal_tile_14_7_to_tile_14_6_2),
		.out_wire_2_3(horizontal_tile_14_7_to_tile_14_6_3),
		.in_wire_2_0(horizontal_tile_14_6_to_tile_14_7_0),
		.in_wire_2_1(horizontal_tile_14_6_to_tile_14_7_1),
		.in_wire_2_2(horizontal_tile_14_6_to_tile_14_7_2),
		.in_wire_2_3(horizontal_tile_14_6_to_tile_14_7_3),
		.out_wire_0_0(horizontal_tile_14_7_to_tile_14_8_0),
		.out_wire_0_1(horizontal_tile_14_7_to_tile_14_8_1),
		.out_wire_0_2(horizontal_tile_14_7_to_tile_14_8_2),
		.out_wire_0_3(horizontal_tile_14_7_to_tile_14_8_3),
		.in_wire_0_0(horizontal_tile_14_8_to_tile_14_7_0),
		.in_wire_0_1(horizontal_tile_14_8_to_tile_14_7_1),
		.in_wire_0_2(horizontal_tile_14_8_to_tile_14_7_2),
		.in_wire_0_3(horizontal_tile_14_8_to_tile_14_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(456)
	);

	pe_tile pe_tile_14_8(
		.out_wire_3_0(vertical_tile_14_8_to_tile_13_8_0),
		.out_wire_3_1(vertical_tile_14_8_to_tile_13_8_1),
		.out_wire_3_2(vertical_tile_14_8_to_tile_13_8_2),
		.out_wire_3_3(vertical_tile_14_8_to_tile_13_8_3),
		.in_wire_3_0(vertical_tile_13_8_to_tile_14_8_0),
		.in_wire_3_1(vertical_tile_13_8_to_tile_14_8_1),
		.in_wire_3_2(vertical_tile_13_8_to_tile_14_8_2),
		.in_wire_3_3(vertical_tile_13_8_to_tile_14_8_3),
		.out_wire_1_0(vertical_tile_14_8_to_tile_15_8_0),
		.out_wire_1_1(vertical_tile_14_8_to_tile_15_8_1),
		.out_wire_1_2(vertical_tile_14_8_to_tile_15_8_2),
		.out_wire_1_3(vertical_tile_14_8_to_tile_15_8_3),
		.in_wire_1_0(vertical_tile_15_8_to_tile_14_8_0),
		.in_wire_1_1(vertical_tile_15_8_to_tile_14_8_1),
		.in_wire_1_2(vertical_tile_15_8_to_tile_14_8_2),
		.in_wire_1_3(vertical_tile_15_8_to_tile_14_8_3),
		.out_wire_2_0(horizontal_tile_14_8_to_tile_14_7_0),
		.out_wire_2_1(horizontal_tile_14_8_to_tile_14_7_1),
		.out_wire_2_2(horizontal_tile_14_8_to_tile_14_7_2),
		.out_wire_2_3(horizontal_tile_14_8_to_tile_14_7_3),
		.in_wire_2_0(horizontal_tile_14_7_to_tile_14_8_0),
		.in_wire_2_1(horizontal_tile_14_7_to_tile_14_8_1),
		.in_wire_2_2(horizontal_tile_14_7_to_tile_14_8_2),
		.in_wire_2_3(horizontal_tile_14_7_to_tile_14_8_3),
		.out_wire_0_0(horizontal_tile_14_8_to_tile_14_9_0),
		.out_wire_0_1(horizontal_tile_14_8_to_tile_14_9_1),
		.out_wire_0_2(horizontal_tile_14_8_to_tile_14_9_2),
		.out_wire_0_3(horizontal_tile_14_8_to_tile_14_9_3),
		.in_wire_0_0(horizontal_tile_14_9_to_tile_14_8_0),
		.in_wire_0_1(horizontal_tile_14_9_to_tile_14_8_1),
		.in_wire_0_2(horizontal_tile_14_9_to_tile_14_8_2),
		.in_wire_0_3(horizontal_tile_14_9_to_tile_14_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(457)
	);

	pe_tile pe_tile_14_9(
		.out_wire_3_0(vertical_tile_14_9_to_tile_13_9_0),
		.out_wire_3_1(vertical_tile_14_9_to_tile_13_9_1),
		.out_wire_3_2(vertical_tile_14_9_to_tile_13_9_2),
		.out_wire_3_3(vertical_tile_14_9_to_tile_13_9_3),
		.in_wire_3_0(vertical_tile_13_9_to_tile_14_9_0),
		.in_wire_3_1(vertical_tile_13_9_to_tile_14_9_1),
		.in_wire_3_2(vertical_tile_13_9_to_tile_14_9_2),
		.in_wire_3_3(vertical_tile_13_9_to_tile_14_9_3),
		.out_wire_1_0(vertical_tile_14_9_to_tile_15_9_0),
		.out_wire_1_1(vertical_tile_14_9_to_tile_15_9_1),
		.out_wire_1_2(vertical_tile_14_9_to_tile_15_9_2),
		.out_wire_1_3(vertical_tile_14_9_to_tile_15_9_3),
		.in_wire_1_0(vertical_tile_15_9_to_tile_14_9_0),
		.in_wire_1_1(vertical_tile_15_9_to_tile_14_9_1),
		.in_wire_1_2(vertical_tile_15_9_to_tile_14_9_2),
		.in_wire_1_3(vertical_tile_15_9_to_tile_14_9_3),
		.out_wire_2_0(horizontal_tile_14_9_to_tile_14_8_0),
		.out_wire_2_1(horizontal_tile_14_9_to_tile_14_8_1),
		.out_wire_2_2(horizontal_tile_14_9_to_tile_14_8_2),
		.out_wire_2_3(horizontal_tile_14_9_to_tile_14_8_3),
		.in_wire_2_0(horizontal_tile_14_8_to_tile_14_9_0),
		.in_wire_2_1(horizontal_tile_14_8_to_tile_14_9_1),
		.in_wire_2_2(horizontal_tile_14_8_to_tile_14_9_2),
		.in_wire_2_3(horizontal_tile_14_8_to_tile_14_9_3),
		.out_wire_0_0(horizontal_tile_14_9_to_tile_14_10_0),
		.out_wire_0_1(horizontal_tile_14_9_to_tile_14_10_1),
		.out_wire_0_2(horizontal_tile_14_9_to_tile_14_10_2),
		.out_wire_0_3(horizontal_tile_14_9_to_tile_14_10_3),
		.in_wire_0_0(horizontal_tile_14_10_to_tile_14_9_0),
		.in_wire_0_1(horizontal_tile_14_10_to_tile_14_9_1),
		.in_wire_0_2(horizontal_tile_14_10_to_tile_14_9_2),
		.in_wire_0_3(horizontal_tile_14_10_to_tile_14_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(458)
	);

	pe_tile pe_tile_14_10(
		.out_wire_3_0(vertical_tile_14_10_to_tile_13_10_0),
		.out_wire_3_1(vertical_tile_14_10_to_tile_13_10_1),
		.out_wire_3_2(vertical_tile_14_10_to_tile_13_10_2),
		.out_wire_3_3(vertical_tile_14_10_to_tile_13_10_3),
		.in_wire_3_0(vertical_tile_13_10_to_tile_14_10_0),
		.in_wire_3_1(vertical_tile_13_10_to_tile_14_10_1),
		.in_wire_3_2(vertical_tile_13_10_to_tile_14_10_2),
		.in_wire_3_3(vertical_tile_13_10_to_tile_14_10_3),
		.out_wire_1_0(vertical_tile_14_10_to_tile_15_10_0),
		.out_wire_1_1(vertical_tile_14_10_to_tile_15_10_1),
		.out_wire_1_2(vertical_tile_14_10_to_tile_15_10_2),
		.out_wire_1_3(vertical_tile_14_10_to_tile_15_10_3),
		.in_wire_1_0(vertical_tile_15_10_to_tile_14_10_0),
		.in_wire_1_1(vertical_tile_15_10_to_tile_14_10_1),
		.in_wire_1_2(vertical_tile_15_10_to_tile_14_10_2),
		.in_wire_1_3(vertical_tile_15_10_to_tile_14_10_3),
		.out_wire_2_0(horizontal_tile_14_10_to_tile_14_9_0),
		.out_wire_2_1(horizontal_tile_14_10_to_tile_14_9_1),
		.out_wire_2_2(horizontal_tile_14_10_to_tile_14_9_2),
		.out_wire_2_3(horizontal_tile_14_10_to_tile_14_9_3),
		.in_wire_2_0(horizontal_tile_14_9_to_tile_14_10_0),
		.in_wire_2_1(horizontal_tile_14_9_to_tile_14_10_1),
		.in_wire_2_2(horizontal_tile_14_9_to_tile_14_10_2),
		.in_wire_2_3(horizontal_tile_14_9_to_tile_14_10_3),
		.out_wire_0_0(horizontal_tile_14_10_to_tile_14_11_0),
		.out_wire_0_1(horizontal_tile_14_10_to_tile_14_11_1),
		.out_wire_0_2(horizontal_tile_14_10_to_tile_14_11_2),
		.out_wire_0_3(horizontal_tile_14_10_to_tile_14_11_3),
		.in_wire_0_0(horizontal_tile_14_11_to_tile_14_10_0),
		.in_wire_0_1(horizontal_tile_14_11_to_tile_14_10_1),
		.in_wire_0_2(horizontal_tile_14_11_to_tile_14_10_2),
		.in_wire_0_3(horizontal_tile_14_11_to_tile_14_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(459)
	);

	pe_tile pe_tile_14_11(
		.out_wire_3_0(vertical_tile_14_11_to_tile_13_11_0),
		.out_wire_3_1(vertical_tile_14_11_to_tile_13_11_1),
		.out_wire_3_2(vertical_tile_14_11_to_tile_13_11_2),
		.out_wire_3_3(vertical_tile_14_11_to_tile_13_11_3),
		.in_wire_3_0(vertical_tile_13_11_to_tile_14_11_0),
		.in_wire_3_1(vertical_tile_13_11_to_tile_14_11_1),
		.in_wire_3_2(vertical_tile_13_11_to_tile_14_11_2),
		.in_wire_3_3(vertical_tile_13_11_to_tile_14_11_3),
		.out_wire_1_0(vertical_tile_14_11_to_tile_15_11_0),
		.out_wire_1_1(vertical_tile_14_11_to_tile_15_11_1),
		.out_wire_1_2(vertical_tile_14_11_to_tile_15_11_2),
		.out_wire_1_3(vertical_tile_14_11_to_tile_15_11_3),
		.in_wire_1_0(vertical_tile_15_11_to_tile_14_11_0),
		.in_wire_1_1(vertical_tile_15_11_to_tile_14_11_1),
		.in_wire_1_2(vertical_tile_15_11_to_tile_14_11_2),
		.in_wire_1_3(vertical_tile_15_11_to_tile_14_11_3),
		.out_wire_2_0(horizontal_tile_14_11_to_tile_14_10_0),
		.out_wire_2_1(horizontal_tile_14_11_to_tile_14_10_1),
		.out_wire_2_2(horizontal_tile_14_11_to_tile_14_10_2),
		.out_wire_2_3(horizontal_tile_14_11_to_tile_14_10_3),
		.in_wire_2_0(horizontal_tile_14_10_to_tile_14_11_0),
		.in_wire_2_1(horizontal_tile_14_10_to_tile_14_11_1),
		.in_wire_2_2(horizontal_tile_14_10_to_tile_14_11_2),
		.in_wire_2_3(horizontal_tile_14_10_to_tile_14_11_3),
		.out_wire_0_0(horizontal_tile_14_11_to_tile_14_12_0),
		.out_wire_0_1(horizontal_tile_14_11_to_tile_14_12_1),
		.out_wire_0_2(horizontal_tile_14_11_to_tile_14_12_2),
		.out_wire_0_3(horizontal_tile_14_11_to_tile_14_12_3),
		.in_wire_0_0(horizontal_tile_14_12_to_tile_14_11_0),
		.in_wire_0_1(horizontal_tile_14_12_to_tile_14_11_1),
		.in_wire_0_2(horizontal_tile_14_12_to_tile_14_11_2),
		.in_wire_0_3(horizontal_tile_14_12_to_tile_14_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(460)
	);

	pe_tile pe_tile_14_12(
		.out_wire_3_0(vertical_tile_14_12_to_tile_13_12_0),
		.out_wire_3_1(vertical_tile_14_12_to_tile_13_12_1),
		.out_wire_3_2(vertical_tile_14_12_to_tile_13_12_2),
		.out_wire_3_3(vertical_tile_14_12_to_tile_13_12_3),
		.in_wire_3_0(vertical_tile_13_12_to_tile_14_12_0),
		.in_wire_3_1(vertical_tile_13_12_to_tile_14_12_1),
		.in_wire_3_2(vertical_tile_13_12_to_tile_14_12_2),
		.in_wire_3_3(vertical_tile_13_12_to_tile_14_12_3),
		.out_wire_1_0(vertical_tile_14_12_to_tile_15_12_0),
		.out_wire_1_1(vertical_tile_14_12_to_tile_15_12_1),
		.out_wire_1_2(vertical_tile_14_12_to_tile_15_12_2),
		.out_wire_1_3(vertical_tile_14_12_to_tile_15_12_3),
		.in_wire_1_0(vertical_tile_15_12_to_tile_14_12_0),
		.in_wire_1_1(vertical_tile_15_12_to_tile_14_12_1),
		.in_wire_1_2(vertical_tile_15_12_to_tile_14_12_2),
		.in_wire_1_3(vertical_tile_15_12_to_tile_14_12_3),
		.out_wire_2_0(horizontal_tile_14_12_to_tile_14_11_0),
		.out_wire_2_1(horizontal_tile_14_12_to_tile_14_11_1),
		.out_wire_2_2(horizontal_tile_14_12_to_tile_14_11_2),
		.out_wire_2_3(horizontal_tile_14_12_to_tile_14_11_3),
		.in_wire_2_0(horizontal_tile_14_11_to_tile_14_12_0),
		.in_wire_2_1(horizontal_tile_14_11_to_tile_14_12_1),
		.in_wire_2_2(horizontal_tile_14_11_to_tile_14_12_2),
		.in_wire_2_3(horizontal_tile_14_11_to_tile_14_12_3),
		.out_wire_0_0(horizontal_tile_14_12_to_tile_14_13_0),
		.out_wire_0_1(horizontal_tile_14_12_to_tile_14_13_1),
		.out_wire_0_2(horizontal_tile_14_12_to_tile_14_13_2),
		.out_wire_0_3(horizontal_tile_14_12_to_tile_14_13_3),
		.in_wire_0_0(horizontal_tile_14_13_to_tile_14_12_0),
		.in_wire_0_1(horizontal_tile_14_13_to_tile_14_12_1),
		.in_wire_0_2(horizontal_tile_14_13_to_tile_14_12_2),
		.in_wire_0_3(horizontal_tile_14_13_to_tile_14_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(461)
	);

	pe_tile pe_tile_14_13(
		.out_wire_3_0(vertical_tile_14_13_to_tile_13_13_0),
		.out_wire_3_1(vertical_tile_14_13_to_tile_13_13_1),
		.out_wire_3_2(vertical_tile_14_13_to_tile_13_13_2),
		.out_wire_3_3(vertical_tile_14_13_to_tile_13_13_3),
		.in_wire_3_0(vertical_tile_13_13_to_tile_14_13_0),
		.in_wire_3_1(vertical_tile_13_13_to_tile_14_13_1),
		.in_wire_3_2(vertical_tile_13_13_to_tile_14_13_2),
		.in_wire_3_3(vertical_tile_13_13_to_tile_14_13_3),
		.out_wire_1_0(vertical_tile_14_13_to_tile_15_13_0),
		.out_wire_1_1(vertical_tile_14_13_to_tile_15_13_1),
		.out_wire_1_2(vertical_tile_14_13_to_tile_15_13_2),
		.out_wire_1_3(vertical_tile_14_13_to_tile_15_13_3),
		.in_wire_1_0(vertical_tile_15_13_to_tile_14_13_0),
		.in_wire_1_1(vertical_tile_15_13_to_tile_14_13_1),
		.in_wire_1_2(vertical_tile_15_13_to_tile_14_13_2),
		.in_wire_1_3(vertical_tile_15_13_to_tile_14_13_3),
		.out_wire_2_0(horizontal_tile_14_13_to_tile_14_12_0),
		.out_wire_2_1(horizontal_tile_14_13_to_tile_14_12_1),
		.out_wire_2_2(horizontal_tile_14_13_to_tile_14_12_2),
		.out_wire_2_3(horizontal_tile_14_13_to_tile_14_12_3),
		.in_wire_2_0(horizontal_tile_14_12_to_tile_14_13_0),
		.in_wire_2_1(horizontal_tile_14_12_to_tile_14_13_1),
		.in_wire_2_2(horizontal_tile_14_12_to_tile_14_13_2),
		.in_wire_2_3(horizontal_tile_14_12_to_tile_14_13_3),
		.out_wire_0_0(horizontal_tile_14_13_to_tile_14_14_0),
		.out_wire_0_1(horizontal_tile_14_13_to_tile_14_14_1),
		.out_wire_0_2(horizontal_tile_14_13_to_tile_14_14_2),
		.out_wire_0_3(horizontal_tile_14_13_to_tile_14_14_3),
		.in_wire_0_0(horizontal_tile_14_14_to_tile_14_13_0),
		.in_wire_0_1(horizontal_tile_14_14_to_tile_14_13_1),
		.in_wire_0_2(horizontal_tile_14_14_to_tile_14_13_2),
		.in_wire_0_3(horizontal_tile_14_14_to_tile_14_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(462)
	);

	pe_tile pe_tile_14_14(
		.out_wire_3_0(vertical_tile_14_14_to_tile_13_14_0),
		.out_wire_3_1(vertical_tile_14_14_to_tile_13_14_1),
		.out_wire_3_2(vertical_tile_14_14_to_tile_13_14_2),
		.out_wire_3_3(vertical_tile_14_14_to_tile_13_14_3),
		.in_wire_3_0(vertical_tile_13_14_to_tile_14_14_0),
		.in_wire_3_1(vertical_tile_13_14_to_tile_14_14_1),
		.in_wire_3_2(vertical_tile_13_14_to_tile_14_14_2),
		.in_wire_3_3(vertical_tile_13_14_to_tile_14_14_3),
		.out_wire_1_0(vertical_tile_14_14_to_tile_15_14_0),
		.out_wire_1_1(vertical_tile_14_14_to_tile_15_14_1),
		.out_wire_1_2(vertical_tile_14_14_to_tile_15_14_2),
		.out_wire_1_3(vertical_tile_14_14_to_tile_15_14_3),
		.in_wire_1_0(vertical_tile_15_14_to_tile_14_14_0),
		.in_wire_1_1(vertical_tile_15_14_to_tile_14_14_1),
		.in_wire_1_2(vertical_tile_15_14_to_tile_14_14_2),
		.in_wire_1_3(vertical_tile_15_14_to_tile_14_14_3),
		.out_wire_2_0(horizontal_tile_14_14_to_tile_14_13_0),
		.out_wire_2_1(horizontal_tile_14_14_to_tile_14_13_1),
		.out_wire_2_2(horizontal_tile_14_14_to_tile_14_13_2),
		.out_wire_2_3(horizontal_tile_14_14_to_tile_14_13_3),
		.in_wire_2_0(horizontal_tile_14_13_to_tile_14_14_0),
		.in_wire_2_1(horizontal_tile_14_13_to_tile_14_14_1),
		.in_wire_2_2(horizontal_tile_14_13_to_tile_14_14_2),
		.in_wire_2_3(horizontal_tile_14_13_to_tile_14_14_3),
		.out_wire_0_0(horizontal_tile_14_14_to_tile_14_15_0),
		.out_wire_0_1(horizontal_tile_14_14_to_tile_14_15_1),
		.out_wire_0_2(horizontal_tile_14_14_to_tile_14_15_2),
		.out_wire_0_3(horizontal_tile_14_14_to_tile_14_15_3),
		.in_wire_0_0(horizontal_tile_14_15_to_tile_14_14_0),
		.in_wire_0_1(horizontal_tile_14_15_to_tile_14_14_1),
		.in_wire_0_2(horizontal_tile_14_15_to_tile_14_14_2),
		.in_wire_0_3(horizontal_tile_14_15_to_tile_14_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(463)
	);

	pe_tile pe_tile_14_15(
		.out_wire_3_0(vertical_tile_14_15_to_tile_13_15_0),
		.out_wire_3_1(vertical_tile_14_15_to_tile_13_15_1),
		.out_wire_3_2(vertical_tile_14_15_to_tile_13_15_2),
		.out_wire_3_3(vertical_tile_14_15_to_tile_13_15_3),
		.in_wire_3_0(vertical_tile_13_15_to_tile_14_15_0),
		.in_wire_3_1(vertical_tile_13_15_to_tile_14_15_1),
		.in_wire_3_2(vertical_tile_13_15_to_tile_14_15_2),
		.in_wire_3_3(vertical_tile_13_15_to_tile_14_15_3),
		.out_wire_1_0(vertical_tile_14_15_to_tile_15_15_0),
		.out_wire_1_1(vertical_tile_14_15_to_tile_15_15_1),
		.out_wire_1_2(vertical_tile_14_15_to_tile_15_15_2),
		.out_wire_1_3(vertical_tile_14_15_to_tile_15_15_3),
		.in_wire_1_0(vertical_tile_15_15_to_tile_14_15_0),
		.in_wire_1_1(vertical_tile_15_15_to_tile_14_15_1),
		.in_wire_1_2(vertical_tile_15_15_to_tile_14_15_2),
		.in_wire_1_3(vertical_tile_15_15_to_tile_14_15_3),
		.out_wire_2_0(horizontal_tile_14_15_to_tile_14_14_0),
		.out_wire_2_1(horizontal_tile_14_15_to_tile_14_14_1),
		.out_wire_2_2(horizontal_tile_14_15_to_tile_14_14_2),
		.out_wire_2_3(horizontal_tile_14_15_to_tile_14_14_3),
		.in_wire_2_0(horizontal_tile_14_14_to_tile_14_15_0),
		.in_wire_2_1(horizontal_tile_14_14_to_tile_14_15_1),
		.in_wire_2_2(horizontal_tile_14_14_to_tile_14_15_2),
		.in_wire_2_3(horizontal_tile_14_14_to_tile_14_15_3),
		.out_wire_0_0(horizontal_tile_14_15_to_tile_14_16_0),
		.out_wire_0_1(horizontal_tile_14_15_to_tile_14_16_1),
		.out_wire_0_2(horizontal_tile_14_15_to_tile_14_16_2),
		.out_wire_0_3(horizontal_tile_14_15_to_tile_14_16_3),
		.in_wire_0_0(horizontal_tile_14_16_to_tile_14_15_0),
		.in_wire_0_1(horizontal_tile_14_16_to_tile_14_15_1),
		.in_wire_0_2(horizontal_tile_14_16_to_tile_14_15_2),
		.in_wire_0_3(horizontal_tile_14_16_to_tile_14_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(464)
	);

	pe_tile pe_tile_14_16(
		.out_wire_3_0(vertical_tile_14_16_to_tile_13_16_0),
		.out_wire_3_1(vertical_tile_14_16_to_tile_13_16_1),
		.out_wire_3_2(vertical_tile_14_16_to_tile_13_16_2),
		.out_wire_3_3(vertical_tile_14_16_to_tile_13_16_3),
		.in_wire_3_0(vertical_tile_13_16_to_tile_14_16_0),
		.in_wire_3_1(vertical_tile_13_16_to_tile_14_16_1),
		.in_wire_3_2(vertical_tile_13_16_to_tile_14_16_2),
		.in_wire_3_3(vertical_tile_13_16_to_tile_14_16_3),
		.out_wire_1_0(vertical_tile_14_16_to_tile_15_16_0),
		.out_wire_1_1(vertical_tile_14_16_to_tile_15_16_1),
		.out_wire_1_2(vertical_tile_14_16_to_tile_15_16_2),
		.out_wire_1_3(vertical_tile_14_16_to_tile_15_16_3),
		.in_wire_1_0(vertical_tile_15_16_to_tile_14_16_0),
		.in_wire_1_1(vertical_tile_15_16_to_tile_14_16_1),
		.in_wire_1_2(vertical_tile_15_16_to_tile_14_16_2),
		.in_wire_1_3(vertical_tile_15_16_to_tile_14_16_3),
		.out_wire_2_0(horizontal_tile_14_16_to_tile_14_15_0),
		.out_wire_2_1(horizontal_tile_14_16_to_tile_14_15_1),
		.out_wire_2_2(horizontal_tile_14_16_to_tile_14_15_2),
		.out_wire_2_3(horizontal_tile_14_16_to_tile_14_15_3),
		.in_wire_2_0(horizontal_tile_14_15_to_tile_14_16_0),
		.in_wire_2_1(horizontal_tile_14_15_to_tile_14_16_1),
		.in_wire_2_2(horizontal_tile_14_15_to_tile_14_16_2),
		.in_wire_2_3(horizontal_tile_14_15_to_tile_14_16_3),
		.out_wire_0_0(horizontal_tile_14_16_to_tile_14_17_0),
		.out_wire_0_1(horizontal_tile_14_16_to_tile_14_17_1),
		.out_wire_0_2(horizontal_tile_14_16_to_tile_14_17_2),
		.out_wire_0_3(horizontal_tile_14_16_to_tile_14_17_3),
		.in_wire_0_0(horizontal_tile_14_17_to_tile_14_16_0),
		.in_wire_0_1(horizontal_tile_14_17_to_tile_14_16_1),
		.in_wire_0_2(horizontal_tile_14_17_to_tile_14_16_2),
		.in_wire_0_3(horizontal_tile_14_17_to_tile_14_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(465)
	);

	pe_tile pe_tile_14_17(
		.out_wire_3_0(vertical_tile_14_17_to_tile_13_17_0),
		.out_wire_3_1(vertical_tile_14_17_to_tile_13_17_1),
		.out_wire_3_2(vertical_tile_14_17_to_tile_13_17_2),
		.out_wire_3_3(vertical_tile_14_17_to_tile_13_17_3),
		.in_wire_3_0(vertical_tile_13_17_to_tile_14_17_0),
		.in_wire_3_1(vertical_tile_13_17_to_tile_14_17_1),
		.in_wire_3_2(vertical_tile_13_17_to_tile_14_17_2),
		.in_wire_3_3(vertical_tile_13_17_to_tile_14_17_3),
		.out_wire_1_0(vertical_tile_14_17_to_tile_15_17_0),
		.out_wire_1_1(vertical_tile_14_17_to_tile_15_17_1),
		.out_wire_1_2(vertical_tile_14_17_to_tile_15_17_2),
		.out_wire_1_3(vertical_tile_14_17_to_tile_15_17_3),
		.in_wire_1_0(vertical_tile_15_17_to_tile_14_17_0),
		.in_wire_1_1(vertical_tile_15_17_to_tile_14_17_1),
		.in_wire_1_2(vertical_tile_15_17_to_tile_14_17_2),
		.in_wire_1_3(vertical_tile_15_17_to_tile_14_17_3),
		.out_wire_2_0(horizontal_tile_14_17_to_tile_14_16_0),
		.out_wire_2_1(horizontal_tile_14_17_to_tile_14_16_1),
		.out_wire_2_2(horizontal_tile_14_17_to_tile_14_16_2),
		.out_wire_2_3(horizontal_tile_14_17_to_tile_14_16_3),
		.in_wire_2_0(horizontal_tile_14_16_to_tile_14_17_0),
		.in_wire_2_1(horizontal_tile_14_16_to_tile_14_17_1),
		.in_wire_2_2(horizontal_tile_14_16_to_tile_14_17_2),
		.in_wire_2_3(horizontal_tile_14_16_to_tile_14_17_3),
		.out_wire_0_0(horizontal_tile_14_17_to_tile_14_18_0),
		.out_wire_0_1(horizontal_tile_14_17_to_tile_14_18_1),
		.out_wire_0_2(horizontal_tile_14_17_to_tile_14_18_2),
		.out_wire_0_3(horizontal_tile_14_17_to_tile_14_18_3),
		.in_wire_0_0(horizontal_tile_14_18_to_tile_14_17_0),
		.in_wire_0_1(horizontal_tile_14_18_to_tile_14_17_1),
		.in_wire_0_2(horizontal_tile_14_18_to_tile_14_17_2),
		.in_wire_0_3(horizontal_tile_14_18_to_tile_14_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(466)
	);

	pe_tile pe_tile_14_18(
		.out_wire_3_0(vertical_tile_14_18_to_tile_13_18_0),
		.out_wire_3_1(vertical_tile_14_18_to_tile_13_18_1),
		.out_wire_3_2(vertical_tile_14_18_to_tile_13_18_2),
		.out_wire_3_3(vertical_tile_14_18_to_tile_13_18_3),
		.in_wire_3_0(vertical_tile_13_18_to_tile_14_18_0),
		.in_wire_3_1(vertical_tile_13_18_to_tile_14_18_1),
		.in_wire_3_2(vertical_tile_13_18_to_tile_14_18_2),
		.in_wire_3_3(vertical_tile_13_18_to_tile_14_18_3),
		.out_wire_1_0(vertical_tile_14_18_to_tile_15_18_0),
		.out_wire_1_1(vertical_tile_14_18_to_tile_15_18_1),
		.out_wire_1_2(vertical_tile_14_18_to_tile_15_18_2),
		.out_wire_1_3(vertical_tile_14_18_to_tile_15_18_3),
		.in_wire_1_0(vertical_tile_15_18_to_tile_14_18_0),
		.in_wire_1_1(vertical_tile_15_18_to_tile_14_18_1),
		.in_wire_1_2(vertical_tile_15_18_to_tile_14_18_2),
		.in_wire_1_3(vertical_tile_15_18_to_tile_14_18_3),
		.out_wire_2_0(horizontal_tile_14_18_to_tile_14_17_0),
		.out_wire_2_1(horizontal_tile_14_18_to_tile_14_17_1),
		.out_wire_2_2(horizontal_tile_14_18_to_tile_14_17_2),
		.out_wire_2_3(horizontal_tile_14_18_to_tile_14_17_3),
		.in_wire_2_0(horizontal_tile_14_17_to_tile_14_18_0),
		.in_wire_2_1(horizontal_tile_14_17_to_tile_14_18_1),
		.in_wire_2_2(horizontal_tile_14_17_to_tile_14_18_2),
		.in_wire_2_3(horizontal_tile_14_17_to_tile_14_18_3),
		.out_wire_0_0(horizontal_tile_14_18_to_tile_14_19_0),
		.out_wire_0_1(horizontal_tile_14_18_to_tile_14_19_1),
		.out_wire_0_2(horizontal_tile_14_18_to_tile_14_19_2),
		.out_wire_0_3(horizontal_tile_14_18_to_tile_14_19_3),
		.in_wire_0_0(horizontal_tile_14_19_to_tile_14_18_0),
		.in_wire_0_1(horizontal_tile_14_19_to_tile_14_18_1),
		.in_wire_0_2(horizontal_tile_14_19_to_tile_14_18_2),
		.in_wire_0_3(horizontal_tile_14_19_to_tile_14_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(467)
	);

	pe_tile pe_tile_14_19(
		.out_wire_3_0(vertical_tile_14_19_to_tile_13_19_0),
		.out_wire_3_1(vertical_tile_14_19_to_tile_13_19_1),
		.out_wire_3_2(vertical_tile_14_19_to_tile_13_19_2),
		.out_wire_3_3(vertical_tile_14_19_to_tile_13_19_3),
		.in_wire_3_0(vertical_tile_13_19_to_tile_14_19_0),
		.in_wire_3_1(vertical_tile_13_19_to_tile_14_19_1),
		.in_wire_3_2(vertical_tile_13_19_to_tile_14_19_2),
		.in_wire_3_3(vertical_tile_13_19_to_tile_14_19_3),
		.out_wire_1_0(vertical_tile_14_19_to_tile_15_19_0),
		.out_wire_1_1(vertical_tile_14_19_to_tile_15_19_1),
		.out_wire_1_2(vertical_tile_14_19_to_tile_15_19_2),
		.out_wire_1_3(vertical_tile_14_19_to_tile_15_19_3),
		.in_wire_1_0(vertical_tile_15_19_to_tile_14_19_0),
		.in_wire_1_1(vertical_tile_15_19_to_tile_14_19_1),
		.in_wire_1_2(vertical_tile_15_19_to_tile_14_19_2),
		.in_wire_1_3(vertical_tile_15_19_to_tile_14_19_3),
		.out_wire_2_0(horizontal_tile_14_19_to_tile_14_18_0),
		.out_wire_2_1(horizontal_tile_14_19_to_tile_14_18_1),
		.out_wire_2_2(horizontal_tile_14_19_to_tile_14_18_2),
		.out_wire_2_3(horizontal_tile_14_19_to_tile_14_18_3),
		.in_wire_2_0(horizontal_tile_14_18_to_tile_14_19_0),
		.in_wire_2_1(horizontal_tile_14_18_to_tile_14_19_1),
		.in_wire_2_2(horizontal_tile_14_18_to_tile_14_19_2),
		.in_wire_2_3(horizontal_tile_14_18_to_tile_14_19_3),
		.out_wire_0_0(horizontal_tile_14_19_to_tile_14_20_0),
		.out_wire_0_1(horizontal_tile_14_19_to_tile_14_20_1),
		.out_wire_0_2(horizontal_tile_14_19_to_tile_14_20_2),
		.out_wire_0_3(horizontal_tile_14_19_to_tile_14_20_3),
		.in_wire_0_0(horizontal_tile_14_20_to_tile_14_19_0),
		.in_wire_0_1(horizontal_tile_14_20_to_tile_14_19_1),
		.in_wire_0_2(horizontal_tile_14_20_to_tile_14_19_2),
		.in_wire_0_3(horizontal_tile_14_20_to_tile_14_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(468)
	);

	pe_tile pe_tile_14_20(
		.out_wire_3_0(vertical_tile_14_20_to_tile_13_20_0),
		.out_wire_3_1(vertical_tile_14_20_to_tile_13_20_1),
		.out_wire_3_2(vertical_tile_14_20_to_tile_13_20_2),
		.out_wire_3_3(vertical_tile_14_20_to_tile_13_20_3),
		.in_wire_3_0(vertical_tile_13_20_to_tile_14_20_0),
		.in_wire_3_1(vertical_tile_13_20_to_tile_14_20_1),
		.in_wire_3_2(vertical_tile_13_20_to_tile_14_20_2),
		.in_wire_3_3(vertical_tile_13_20_to_tile_14_20_3),
		.out_wire_1_0(vertical_tile_14_20_to_tile_15_20_0),
		.out_wire_1_1(vertical_tile_14_20_to_tile_15_20_1),
		.out_wire_1_2(vertical_tile_14_20_to_tile_15_20_2),
		.out_wire_1_3(vertical_tile_14_20_to_tile_15_20_3),
		.in_wire_1_0(vertical_tile_15_20_to_tile_14_20_0),
		.in_wire_1_1(vertical_tile_15_20_to_tile_14_20_1),
		.in_wire_1_2(vertical_tile_15_20_to_tile_14_20_2),
		.in_wire_1_3(vertical_tile_15_20_to_tile_14_20_3),
		.out_wire_2_0(horizontal_tile_14_20_to_tile_14_19_0),
		.out_wire_2_1(horizontal_tile_14_20_to_tile_14_19_1),
		.out_wire_2_2(horizontal_tile_14_20_to_tile_14_19_2),
		.out_wire_2_3(horizontal_tile_14_20_to_tile_14_19_3),
		.in_wire_2_0(horizontal_tile_14_19_to_tile_14_20_0),
		.in_wire_2_1(horizontal_tile_14_19_to_tile_14_20_1),
		.in_wire_2_2(horizontal_tile_14_19_to_tile_14_20_2),
		.in_wire_2_3(horizontal_tile_14_19_to_tile_14_20_3),
		.out_wire_0_0(horizontal_tile_14_20_to_tile_14_21_0),
		.out_wire_0_1(horizontal_tile_14_20_to_tile_14_21_1),
		.out_wire_0_2(horizontal_tile_14_20_to_tile_14_21_2),
		.out_wire_0_3(horizontal_tile_14_20_to_tile_14_21_3),
		.in_wire_0_0(horizontal_tile_14_21_to_tile_14_20_0),
		.in_wire_0_1(horizontal_tile_14_21_to_tile_14_20_1),
		.in_wire_0_2(horizontal_tile_14_21_to_tile_14_20_2),
		.in_wire_0_3(horizontal_tile_14_21_to_tile_14_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(469)
	);

	pe_tile pe_tile_14_21(
		.out_wire_3_0(vertical_tile_14_21_to_tile_13_21_0),
		.out_wire_3_1(vertical_tile_14_21_to_tile_13_21_1),
		.out_wire_3_2(vertical_tile_14_21_to_tile_13_21_2),
		.out_wire_3_3(vertical_tile_14_21_to_tile_13_21_3),
		.in_wire_3_0(vertical_tile_13_21_to_tile_14_21_0),
		.in_wire_3_1(vertical_tile_13_21_to_tile_14_21_1),
		.in_wire_3_2(vertical_tile_13_21_to_tile_14_21_2),
		.in_wire_3_3(vertical_tile_13_21_to_tile_14_21_3),
		.out_wire_1_0(vertical_tile_14_21_to_tile_15_21_0),
		.out_wire_1_1(vertical_tile_14_21_to_tile_15_21_1),
		.out_wire_1_2(vertical_tile_14_21_to_tile_15_21_2),
		.out_wire_1_3(vertical_tile_14_21_to_tile_15_21_3),
		.in_wire_1_0(vertical_tile_15_21_to_tile_14_21_0),
		.in_wire_1_1(vertical_tile_15_21_to_tile_14_21_1),
		.in_wire_1_2(vertical_tile_15_21_to_tile_14_21_2),
		.in_wire_1_3(vertical_tile_15_21_to_tile_14_21_3),
		.out_wire_2_0(horizontal_tile_14_21_to_tile_14_20_0),
		.out_wire_2_1(horizontal_tile_14_21_to_tile_14_20_1),
		.out_wire_2_2(horizontal_tile_14_21_to_tile_14_20_2),
		.out_wire_2_3(horizontal_tile_14_21_to_tile_14_20_3),
		.in_wire_2_0(horizontal_tile_14_20_to_tile_14_21_0),
		.in_wire_2_1(horizontal_tile_14_20_to_tile_14_21_1),
		.in_wire_2_2(horizontal_tile_14_20_to_tile_14_21_2),
		.in_wire_2_3(horizontal_tile_14_20_to_tile_14_21_3),
		.out_wire_0_0(horizontal_tile_14_21_to_tile_14_22_0),
		.out_wire_0_1(horizontal_tile_14_21_to_tile_14_22_1),
		.out_wire_0_2(horizontal_tile_14_21_to_tile_14_22_2),
		.out_wire_0_3(horizontal_tile_14_21_to_tile_14_22_3),
		.in_wire_0_0(horizontal_tile_14_22_to_tile_14_21_0),
		.in_wire_0_1(horizontal_tile_14_22_to_tile_14_21_1),
		.in_wire_0_2(horizontal_tile_14_22_to_tile_14_21_2),
		.in_wire_0_3(horizontal_tile_14_22_to_tile_14_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(470)
	);

	pe_tile pe_tile_14_22(
		.out_wire_3_0(vertical_tile_14_22_to_tile_13_22_0),
		.out_wire_3_1(vertical_tile_14_22_to_tile_13_22_1),
		.out_wire_3_2(vertical_tile_14_22_to_tile_13_22_2),
		.out_wire_3_3(vertical_tile_14_22_to_tile_13_22_3),
		.in_wire_3_0(vertical_tile_13_22_to_tile_14_22_0),
		.in_wire_3_1(vertical_tile_13_22_to_tile_14_22_1),
		.in_wire_3_2(vertical_tile_13_22_to_tile_14_22_2),
		.in_wire_3_3(vertical_tile_13_22_to_tile_14_22_3),
		.out_wire_1_0(vertical_tile_14_22_to_tile_15_22_0),
		.out_wire_1_1(vertical_tile_14_22_to_tile_15_22_1),
		.out_wire_1_2(vertical_tile_14_22_to_tile_15_22_2),
		.out_wire_1_3(vertical_tile_14_22_to_tile_15_22_3),
		.in_wire_1_0(vertical_tile_15_22_to_tile_14_22_0),
		.in_wire_1_1(vertical_tile_15_22_to_tile_14_22_1),
		.in_wire_1_2(vertical_tile_15_22_to_tile_14_22_2),
		.in_wire_1_3(vertical_tile_15_22_to_tile_14_22_3),
		.out_wire_2_0(horizontal_tile_14_22_to_tile_14_21_0),
		.out_wire_2_1(horizontal_tile_14_22_to_tile_14_21_1),
		.out_wire_2_2(horizontal_tile_14_22_to_tile_14_21_2),
		.out_wire_2_3(horizontal_tile_14_22_to_tile_14_21_3),
		.in_wire_2_0(horizontal_tile_14_21_to_tile_14_22_0),
		.in_wire_2_1(horizontal_tile_14_21_to_tile_14_22_1),
		.in_wire_2_2(horizontal_tile_14_21_to_tile_14_22_2),
		.in_wire_2_3(horizontal_tile_14_21_to_tile_14_22_3),
		.out_wire_0_0(horizontal_tile_14_22_to_tile_14_23_0),
		.out_wire_0_1(horizontal_tile_14_22_to_tile_14_23_1),
		.out_wire_0_2(horizontal_tile_14_22_to_tile_14_23_2),
		.out_wire_0_3(horizontal_tile_14_22_to_tile_14_23_3),
		.in_wire_0_0(horizontal_tile_14_23_to_tile_14_22_0),
		.in_wire_0_1(horizontal_tile_14_23_to_tile_14_22_1),
		.in_wire_0_2(horizontal_tile_14_23_to_tile_14_22_2),
		.in_wire_0_3(horizontal_tile_14_23_to_tile_14_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(471)
	);

	pe_tile pe_tile_14_23(
		.out_wire_3_0(vertical_tile_14_23_to_tile_13_23_0),
		.out_wire_3_1(vertical_tile_14_23_to_tile_13_23_1),
		.out_wire_3_2(vertical_tile_14_23_to_tile_13_23_2),
		.out_wire_3_3(vertical_tile_14_23_to_tile_13_23_3),
		.in_wire_3_0(vertical_tile_13_23_to_tile_14_23_0),
		.in_wire_3_1(vertical_tile_13_23_to_tile_14_23_1),
		.in_wire_3_2(vertical_tile_13_23_to_tile_14_23_2),
		.in_wire_3_3(vertical_tile_13_23_to_tile_14_23_3),
		.out_wire_1_0(vertical_tile_14_23_to_tile_15_23_0),
		.out_wire_1_1(vertical_tile_14_23_to_tile_15_23_1),
		.out_wire_1_2(vertical_tile_14_23_to_tile_15_23_2),
		.out_wire_1_3(vertical_tile_14_23_to_tile_15_23_3),
		.in_wire_1_0(vertical_tile_15_23_to_tile_14_23_0),
		.in_wire_1_1(vertical_tile_15_23_to_tile_14_23_1),
		.in_wire_1_2(vertical_tile_15_23_to_tile_14_23_2),
		.in_wire_1_3(vertical_tile_15_23_to_tile_14_23_3),
		.out_wire_2_0(horizontal_tile_14_23_to_tile_14_22_0),
		.out_wire_2_1(horizontal_tile_14_23_to_tile_14_22_1),
		.out_wire_2_2(horizontal_tile_14_23_to_tile_14_22_2),
		.out_wire_2_3(horizontal_tile_14_23_to_tile_14_22_3),
		.in_wire_2_0(horizontal_tile_14_22_to_tile_14_23_0),
		.in_wire_2_1(horizontal_tile_14_22_to_tile_14_23_1),
		.in_wire_2_2(horizontal_tile_14_22_to_tile_14_23_2),
		.in_wire_2_3(horizontal_tile_14_22_to_tile_14_23_3),
		.out_wire_0_0(horizontal_tile_14_23_to_tile_14_24_0),
		.out_wire_0_1(horizontal_tile_14_23_to_tile_14_24_1),
		.out_wire_0_2(horizontal_tile_14_23_to_tile_14_24_2),
		.out_wire_0_3(horizontal_tile_14_23_to_tile_14_24_3),
		.in_wire_0_0(horizontal_tile_14_24_to_tile_14_23_0),
		.in_wire_0_1(horizontal_tile_14_24_to_tile_14_23_1),
		.in_wire_0_2(horizontal_tile_14_24_to_tile_14_23_2),
		.in_wire_0_3(horizontal_tile_14_24_to_tile_14_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(472)
	);

	pe_tile pe_tile_14_24(
		.out_wire_3_0(vertical_tile_14_24_to_tile_13_24_0),
		.out_wire_3_1(vertical_tile_14_24_to_tile_13_24_1),
		.out_wire_3_2(vertical_tile_14_24_to_tile_13_24_2),
		.out_wire_3_3(vertical_tile_14_24_to_tile_13_24_3),
		.in_wire_3_0(vertical_tile_13_24_to_tile_14_24_0),
		.in_wire_3_1(vertical_tile_13_24_to_tile_14_24_1),
		.in_wire_3_2(vertical_tile_13_24_to_tile_14_24_2),
		.in_wire_3_3(vertical_tile_13_24_to_tile_14_24_3),
		.out_wire_1_0(vertical_tile_14_24_to_tile_15_24_0),
		.out_wire_1_1(vertical_tile_14_24_to_tile_15_24_1),
		.out_wire_1_2(vertical_tile_14_24_to_tile_15_24_2),
		.out_wire_1_3(vertical_tile_14_24_to_tile_15_24_3),
		.in_wire_1_0(vertical_tile_15_24_to_tile_14_24_0),
		.in_wire_1_1(vertical_tile_15_24_to_tile_14_24_1),
		.in_wire_1_2(vertical_tile_15_24_to_tile_14_24_2),
		.in_wire_1_3(vertical_tile_15_24_to_tile_14_24_3),
		.out_wire_2_0(horizontal_tile_14_24_to_tile_14_23_0),
		.out_wire_2_1(horizontal_tile_14_24_to_tile_14_23_1),
		.out_wire_2_2(horizontal_tile_14_24_to_tile_14_23_2),
		.out_wire_2_3(horizontal_tile_14_24_to_tile_14_23_3),
		.in_wire_2_0(horizontal_tile_14_23_to_tile_14_24_0),
		.in_wire_2_1(horizontal_tile_14_23_to_tile_14_24_1),
		.in_wire_2_2(horizontal_tile_14_23_to_tile_14_24_2),
		.in_wire_2_3(horizontal_tile_14_23_to_tile_14_24_3),
		.out_wire_0_0(horizontal_tile_14_24_to_tile_14_25_0),
		.out_wire_0_1(horizontal_tile_14_24_to_tile_14_25_1),
		.out_wire_0_2(horizontal_tile_14_24_to_tile_14_25_2),
		.out_wire_0_3(horizontal_tile_14_24_to_tile_14_25_3),
		.in_wire_0_0(horizontal_tile_14_25_to_tile_14_24_0),
		.in_wire_0_1(horizontal_tile_14_25_to_tile_14_24_1),
		.in_wire_0_2(horizontal_tile_14_25_to_tile_14_24_2),
		.in_wire_0_3(horizontal_tile_14_25_to_tile_14_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(473)
	);

	pe_tile pe_tile_14_25(
		.out_wire_3_0(vertical_tile_14_25_to_tile_13_25_0),
		.out_wire_3_1(vertical_tile_14_25_to_tile_13_25_1),
		.out_wire_3_2(vertical_tile_14_25_to_tile_13_25_2),
		.out_wire_3_3(vertical_tile_14_25_to_tile_13_25_3),
		.in_wire_3_0(vertical_tile_13_25_to_tile_14_25_0),
		.in_wire_3_1(vertical_tile_13_25_to_tile_14_25_1),
		.in_wire_3_2(vertical_tile_13_25_to_tile_14_25_2),
		.in_wire_3_3(vertical_tile_13_25_to_tile_14_25_3),
		.out_wire_1_0(vertical_tile_14_25_to_tile_15_25_0),
		.out_wire_1_1(vertical_tile_14_25_to_tile_15_25_1),
		.out_wire_1_2(vertical_tile_14_25_to_tile_15_25_2),
		.out_wire_1_3(vertical_tile_14_25_to_tile_15_25_3),
		.in_wire_1_0(vertical_tile_15_25_to_tile_14_25_0),
		.in_wire_1_1(vertical_tile_15_25_to_tile_14_25_1),
		.in_wire_1_2(vertical_tile_15_25_to_tile_14_25_2),
		.in_wire_1_3(vertical_tile_15_25_to_tile_14_25_3),
		.out_wire_2_0(horizontal_tile_14_25_to_tile_14_24_0),
		.out_wire_2_1(horizontal_tile_14_25_to_tile_14_24_1),
		.out_wire_2_2(horizontal_tile_14_25_to_tile_14_24_2),
		.out_wire_2_3(horizontal_tile_14_25_to_tile_14_24_3),
		.in_wire_2_0(horizontal_tile_14_24_to_tile_14_25_0),
		.in_wire_2_1(horizontal_tile_14_24_to_tile_14_25_1),
		.in_wire_2_2(horizontal_tile_14_24_to_tile_14_25_2),
		.in_wire_2_3(horizontal_tile_14_24_to_tile_14_25_3),
		.out_wire_0_0(horizontal_tile_14_25_to_tile_14_26_0),
		.out_wire_0_1(horizontal_tile_14_25_to_tile_14_26_1),
		.out_wire_0_2(horizontal_tile_14_25_to_tile_14_26_2),
		.out_wire_0_3(horizontal_tile_14_25_to_tile_14_26_3),
		.in_wire_0_0(horizontal_tile_14_26_to_tile_14_25_0),
		.in_wire_0_1(horizontal_tile_14_26_to_tile_14_25_1),
		.in_wire_0_2(horizontal_tile_14_26_to_tile_14_25_2),
		.in_wire_0_3(horizontal_tile_14_26_to_tile_14_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(474)
	);

	pe_tile pe_tile_14_26(
		.out_wire_3_0(vertical_tile_14_26_to_tile_13_26_0),
		.out_wire_3_1(vertical_tile_14_26_to_tile_13_26_1),
		.out_wire_3_2(vertical_tile_14_26_to_tile_13_26_2),
		.out_wire_3_3(vertical_tile_14_26_to_tile_13_26_3),
		.in_wire_3_0(vertical_tile_13_26_to_tile_14_26_0),
		.in_wire_3_1(vertical_tile_13_26_to_tile_14_26_1),
		.in_wire_3_2(vertical_tile_13_26_to_tile_14_26_2),
		.in_wire_3_3(vertical_tile_13_26_to_tile_14_26_3),
		.out_wire_1_0(vertical_tile_14_26_to_tile_15_26_0),
		.out_wire_1_1(vertical_tile_14_26_to_tile_15_26_1),
		.out_wire_1_2(vertical_tile_14_26_to_tile_15_26_2),
		.out_wire_1_3(vertical_tile_14_26_to_tile_15_26_3),
		.in_wire_1_0(vertical_tile_15_26_to_tile_14_26_0),
		.in_wire_1_1(vertical_tile_15_26_to_tile_14_26_1),
		.in_wire_1_2(vertical_tile_15_26_to_tile_14_26_2),
		.in_wire_1_3(vertical_tile_15_26_to_tile_14_26_3),
		.out_wire_2_0(horizontal_tile_14_26_to_tile_14_25_0),
		.out_wire_2_1(horizontal_tile_14_26_to_tile_14_25_1),
		.out_wire_2_2(horizontal_tile_14_26_to_tile_14_25_2),
		.out_wire_2_3(horizontal_tile_14_26_to_tile_14_25_3),
		.in_wire_2_0(horizontal_tile_14_25_to_tile_14_26_0),
		.in_wire_2_1(horizontal_tile_14_25_to_tile_14_26_1),
		.in_wire_2_2(horizontal_tile_14_25_to_tile_14_26_2),
		.in_wire_2_3(horizontal_tile_14_25_to_tile_14_26_3),
		.out_wire_0_0(horizontal_tile_14_26_to_tile_14_27_0),
		.out_wire_0_1(horizontal_tile_14_26_to_tile_14_27_1),
		.out_wire_0_2(horizontal_tile_14_26_to_tile_14_27_2),
		.out_wire_0_3(horizontal_tile_14_26_to_tile_14_27_3),
		.in_wire_0_0(horizontal_tile_14_27_to_tile_14_26_0),
		.in_wire_0_1(horizontal_tile_14_27_to_tile_14_26_1),
		.in_wire_0_2(horizontal_tile_14_27_to_tile_14_26_2),
		.in_wire_0_3(horizontal_tile_14_27_to_tile_14_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(475)
	);

	pe_tile pe_tile_14_27(
		.out_wire_3_0(vertical_tile_14_27_to_tile_13_27_0),
		.out_wire_3_1(vertical_tile_14_27_to_tile_13_27_1),
		.out_wire_3_2(vertical_tile_14_27_to_tile_13_27_2),
		.out_wire_3_3(vertical_tile_14_27_to_tile_13_27_3),
		.in_wire_3_0(vertical_tile_13_27_to_tile_14_27_0),
		.in_wire_3_1(vertical_tile_13_27_to_tile_14_27_1),
		.in_wire_3_2(vertical_tile_13_27_to_tile_14_27_2),
		.in_wire_3_3(vertical_tile_13_27_to_tile_14_27_3),
		.out_wire_1_0(vertical_tile_14_27_to_tile_15_27_0),
		.out_wire_1_1(vertical_tile_14_27_to_tile_15_27_1),
		.out_wire_1_2(vertical_tile_14_27_to_tile_15_27_2),
		.out_wire_1_3(vertical_tile_14_27_to_tile_15_27_3),
		.in_wire_1_0(vertical_tile_15_27_to_tile_14_27_0),
		.in_wire_1_1(vertical_tile_15_27_to_tile_14_27_1),
		.in_wire_1_2(vertical_tile_15_27_to_tile_14_27_2),
		.in_wire_1_3(vertical_tile_15_27_to_tile_14_27_3),
		.out_wire_2_0(horizontal_tile_14_27_to_tile_14_26_0),
		.out_wire_2_1(horizontal_tile_14_27_to_tile_14_26_1),
		.out_wire_2_2(horizontal_tile_14_27_to_tile_14_26_2),
		.out_wire_2_3(horizontal_tile_14_27_to_tile_14_26_3),
		.in_wire_2_0(horizontal_tile_14_26_to_tile_14_27_0),
		.in_wire_2_1(horizontal_tile_14_26_to_tile_14_27_1),
		.in_wire_2_2(horizontal_tile_14_26_to_tile_14_27_2),
		.in_wire_2_3(horizontal_tile_14_26_to_tile_14_27_3),
		.out_wire_0_0(horizontal_tile_14_27_to_tile_14_28_0),
		.out_wire_0_1(horizontal_tile_14_27_to_tile_14_28_1),
		.out_wire_0_2(horizontal_tile_14_27_to_tile_14_28_2),
		.out_wire_0_3(horizontal_tile_14_27_to_tile_14_28_3),
		.in_wire_0_0(horizontal_tile_14_28_to_tile_14_27_0),
		.in_wire_0_1(horizontal_tile_14_28_to_tile_14_27_1),
		.in_wire_0_2(horizontal_tile_14_28_to_tile_14_27_2),
		.in_wire_0_3(horizontal_tile_14_28_to_tile_14_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(476)
	);

	pe_tile pe_tile_14_28(
		.out_wire_3_0(vertical_tile_14_28_to_tile_13_28_0),
		.out_wire_3_1(vertical_tile_14_28_to_tile_13_28_1),
		.out_wire_3_2(vertical_tile_14_28_to_tile_13_28_2),
		.out_wire_3_3(vertical_tile_14_28_to_tile_13_28_3),
		.in_wire_3_0(vertical_tile_13_28_to_tile_14_28_0),
		.in_wire_3_1(vertical_tile_13_28_to_tile_14_28_1),
		.in_wire_3_2(vertical_tile_13_28_to_tile_14_28_2),
		.in_wire_3_3(vertical_tile_13_28_to_tile_14_28_3),
		.out_wire_1_0(vertical_tile_14_28_to_tile_15_28_0),
		.out_wire_1_1(vertical_tile_14_28_to_tile_15_28_1),
		.out_wire_1_2(vertical_tile_14_28_to_tile_15_28_2),
		.out_wire_1_3(vertical_tile_14_28_to_tile_15_28_3),
		.in_wire_1_0(vertical_tile_15_28_to_tile_14_28_0),
		.in_wire_1_1(vertical_tile_15_28_to_tile_14_28_1),
		.in_wire_1_2(vertical_tile_15_28_to_tile_14_28_2),
		.in_wire_1_3(vertical_tile_15_28_to_tile_14_28_3),
		.out_wire_2_0(horizontal_tile_14_28_to_tile_14_27_0),
		.out_wire_2_1(horizontal_tile_14_28_to_tile_14_27_1),
		.out_wire_2_2(horizontal_tile_14_28_to_tile_14_27_2),
		.out_wire_2_3(horizontal_tile_14_28_to_tile_14_27_3),
		.in_wire_2_0(horizontal_tile_14_27_to_tile_14_28_0),
		.in_wire_2_1(horizontal_tile_14_27_to_tile_14_28_1),
		.in_wire_2_2(horizontal_tile_14_27_to_tile_14_28_2),
		.in_wire_2_3(horizontal_tile_14_27_to_tile_14_28_3),
		.out_wire_0_0(horizontal_tile_14_28_to_tile_14_29_0),
		.out_wire_0_1(horizontal_tile_14_28_to_tile_14_29_1),
		.out_wire_0_2(horizontal_tile_14_28_to_tile_14_29_2),
		.out_wire_0_3(horizontal_tile_14_28_to_tile_14_29_3),
		.in_wire_0_0(horizontal_tile_14_29_to_tile_14_28_0),
		.in_wire_0_1(horizontal_tile_14_29_to_tile_14_28_1),
		.in_wire_0_2(horizontal_tile_14_29_to_tile_14_28_2),
		.in_wire_0_3(horizontal_tile_14_29_to_tile_14_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(477)
	);

	pe_tile pe_tile_14_29(
		.out_wire_3_0(vertical_tile_14_29_to_tile_13_29_0),
		.out_wire_3_1(vertical_tile_14_29_to_tile_13_29_1),
		.out_wire_3_2(vertical_tile_14_29_to_tile_13_29_2),
		.out_wire_3_3(vertical_tile_14_29_to_tile_13_29_3),
		.in_wire_3_0(vertical_tile_13_29_to_tile_14_29_0),
		.in_wire_3_1(vertical_tile_13_29_to_tile_14_29_1),
		.in_wire_3_2(vertical_tile_13_29_to_tile_14_29_2),
		.in_wire_3_3(vertical_tile_13_29_to_tile_14_29_3),
		.out_wire_1_0(vertical_tile_14_29_to_tile_15_29_0),
		.out_wire_1_1(vertical_tile_14_29_to_tile_15_29_1),
		.out_wire_1_2(vertical_tile_14_29_to_tile_15_29_2),
		.out_wire_1_3(vertical_tile_14_29_to_tile_15_29_3),
		.in_wire_1_0(vertical_tile_15_29_to_tile_14_29_0),
		.in_wire_1_1(vertical_tile_15_29_to_tile_14_29_1),
		.in_wire_1_2(vertical_tile_15_29_to_tile_14_29_2),
		.in_wire_1_3(vertical_tile_15_29_to_tile_14_29_3),
		.out_wire_2_0(horizontal_tile_14_29_to_tile_14_28_0),
		.out_wire_2_1(horizontal_tile_14_29_to_tile_14_28_1),
		.out_wire_2_2(horizontal_tile_14_29_to_tile_14_28_2),
		.out_wire_2_3(horizontal_tile_14_29_to_tile_14_28_3),
		.in_wire_2_0(horizontal_tile_14_28_to_tile_14_29_0),
		.in_wire_2_1(horizontal_tile_14_28_to_tile_14_29_1),
		.in_wire_2_2(horizontal_tile_14_28_to_tile_14_29_2),
		.in_wire_2_3(horizontal_tile_14_28_to_tile_14_29_3),
		.out_wire_0_0(horizontal_tile_14_29_to_tile_14_30_0),
		.out_wire_0_1(horizontal_tile_14_29_to_tile_14_30_1),
		.out_wire_0_2(horizontal_tile_14_29_to_tile_14_30_2),
		.out_wire_0_3(horizontal_tile_14_29_to_tile_14_30_3),
		.in_wire_0_0(horizontal_tile_14_30_to_tile_14_29_0),
		.in_wire_0_1(horizontal_tile_14_30_to_tile_14_29_1),
		.in_wire_0_2(horizontal_tile_14_30_to_tile_14_29_2),
		.in_wire_0_3(horizontal_tile_14_30_to_tile_14_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(478)
	);

	pe_tile pe_tile_14_30(
		.out_wire_3_0(vertical_tile_14_30_to_tile_13_30_0),
		.out_wire_3_1(vertical_tile_14_30_to_tile_13_30_1),
		.out_wire_3_2(vertical_tile_14_30_to_tile_13_30_2),
		.out_wire_3_3(vertical_tile_14_30_to_tile_13_30_3),
		.in_wire_3_0(vertical_tile_13_30_to_tile_14_30_0),
		.in_wire_3_1(vertical_tile_13_30_to_tile_14_30_1),
		.in_wire_3_2(vertical_tile_13_30_to_tile_14_30_2),
		.in_wire_3_3(vertical_tile_13_30_to_tile_14_30_3),
		.out_wire_1_0(vertical_tile_14_30_to_tile_15_30_0),
		.out_wire_1_1(vertical_tile_14_30_to_tile_15_30_1),
		.out_wire_1_2(vertical_tile_14_30_to_tile_15_30_2),
		.out_wire_1_3(vertical_tile_14_30_to_tile_15_30_3),
		.in_wire_1_0(vertical_tile_15_30_to_tile_14_30_0),
		.in_wire_1_1(vertical_tile_15_30_to_tile_14_30_1),
		.in_wire_1_2(vertical_tile_15_30_to_tile_14_30_2),
		.in_wire_1_3(vertical_tile_15_30_to_tile_14_30_3),
		.out_wire_2_0(horizontal_tile_14_30_to_tile_14_29_0),
		.out_wire_2_1(horizontal_tile_14_30_to_tile_14_29_1),
		.out_wire_2_2(horizontal_tile_14_30_to_tile_14_29_2),
		.out_wire_2_3(horizontal_tile_14_30_to_tile_14_29_3),
		.in_wire_2_0(horizontal_tile_14_29_to_tile_14_30_0),
		.in_wire_2_1(horizontal_tile_14_29_to_tile_14_30_1),
		.in_wire_2_2(horizontal_tile_14_29_to_tile_14_30_2),
		.in_wire_2_3(horizontal_tile_14_29_to_tile_14_30_3),
		.out_wire_0_0(horizontal_tile_14_30_to_tile_14_31_0),
		.out_wire_0_1(horizontal_tile_14_30_to_tile_14_31_1),
		.out_wire_0_2(horizontal_tile_14_30_to_tile_14_31_2),
		.out_wire_0_3(horizontal_tile_14_30_to_tile_14_31_3),
		.in_wire_0_0(horizontal_tile_14_31_to_tile_14_30_0),
		.in_wire_0_1(horizontal_tile_14_31_to_tile_14_30_1),
		.in_wire_0_2(horizontal_tile_14_31_to_tile_14_30_2),
		.in_wire_0_3(horizontal_tile_14_31_to_tile_14_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(479)
	);

	pe_tile_right pe_tile_14_31(
		.out_wire_3_0(vertical_tile_14_31_to_tile_13_31_0),
		.out_wire_3_1(vertical_tile_14_31_to_tile_13_31_1),
		.out_wire_3_2(vertical_tile_14_31_to_tile_13_31_2),
		.out_wire_3_3(vertical_tile_14_31_to_tile_13_31_3),
		.in_wire_3_0(vertical_tile_13_31_to_tile_14_31_0),
		.in_wire_3_1(vertical_tile_13_31_to_tile_14_31_1),
		.in_wire_3_2(vertical_tile_13_31_to_tile_14_31_2),
		.in_wire_3_3(vertical_tile_13_31_to_tile_14_31_3),
		.out_wire_1_0(vertical_tile_14_31_to_tile_15_31_0),
		.out_wire_1_1(vertical_tile_14_31_to_tile_15_31_1),
		.out_wire_1_2(vertical_tile_14_31_to_tile_15_31_2),
		.out_wire_1_3(vertical_tile_14_31_to_tile_15_31_3),
		.in_wire_1_0(vertical_tile_15_31_to_tile_14_31_0),
		.in_wire_1_1(vertical_tile_15_31_to_tile_14_31_1),
		.in_wire_1_2(vertical_tile_15_31_to_tile_14_31_2),
		.in_wire_1_3(vertical_tile_15_31_to_tile_14_31_3),
		.out_wire_2_0(horizontal_tile_14_31_to_tile_14_30_0),
		.out_wire_2_1(horizontal_tile_14_31_to_tile_14_30_1),
		.out_wire_2_2(horizontal_tile_14_31_to_tile_14_30_2),
		.out_wire_2_3(horizontal_tile_14_31_to_tile_14_30_3),
		.in_wire_2_0(horizontal_tile_14_30_to_tile_14_31_0),
		.in_wire_2_1(horizontal_tile_14_30_to_tile_14_31_1),
		.in_wire_2_2(horizontal_tile_14_30_to_tile_14_31_2),
		.in_wire_2_3(horizontal_tile_14_30_to_tile_14_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(480)
	);

	pe_tile_left pe_tile_15_0(
		.out_wire_3_0(vertical_tile_15_0_to_tile_14_0_0),
		.out_wire_3_1(vertical_tile_15_0_to_tile_14_0_1),
		.out_wire_3_2(vertical_tile_15_0_to_tile_14_0_2),
		.out_wire_3_3(vertical_tile_15_0_to_tile_14_0_3),
		.in_wire_3_0(vertical_tile_14_0_to_tile_15_0_0),
		.in_wire_3_1(vertical_tile_14_0_to_tile_15_0_1),
		.in_wire_3_2(vertical_tile_14_0_to_tile_15_0_2),
		.in_wire_3_3(vertical_tile_14_0_to_tile_15_0_3),
		.out_wire_1_0(vertical_tile_15_0_to_tile_16_0_0),
		.out_wire_1_1(vertical_tile_15_0_to_tile_16_0_1),
		.out_wire_1_2(vertical_tile_15_0_to_tile_16_0_2),
		.out_wire_1_3(vertical_tile_15_0_to_tile_16_0_3),
		.in_wire_1_0(vertical_tile_16_0_to_tile_15_0_0),
		.in_wire_1_1(vertical_tile_16_0_to_tile_15_0_1),
		.in_wire_1_2(vertical_tile_16_0_to_tile_15_0_2),
		.in_wire_1_3(vertical_tile_16_0_to_tile_15_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_15_0_to_tile_15_1_0),
		.out_wire_0_1(horizontal_tile_15_0_to_tile_15_1_1),
		.out_wire_0_2(horizontal_tile_15_0_to_tile_15_1_2),
		.out_wire_0_3(horizontal_tile_15_0_to_tile_15_1_3),
		.in_wire_0_0(horizontal_tile_15_1_to_tile_15_0_0),
		.in_wire_0_1(horizontal_tile_15_1_to_tile_15_0_1),
		.in_wire_0_2(horizontal_tile_15_1_to_tile_15_0_2),
		.in_wire_0_3(horizontal_tile_15_1_to_tile_15_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(481)
	);

	pe_tile pe_tile_15_1(
		.out_wire_3_0(vertical_tile_15_1_to_tile_14_1_0),
		.out_wire_3_1(vertical_tile_15_1_to_tile_14_1_1),
		.out_wire_3_2(vertical_tile_15_1_to_tile_14_1_2),
		.out_wire_3_3(vertical_tile_15_1_to_tile_14_1_3),
		.in_wire_3_0(vertical_tile_14_1_to_tile_15_1_0),
		.in_wire_3_1(vertical_tile_14_1_to_tile_15_1_1),
		.in_wire_3_2(vertical_tile_14_1_to_tile_15_1_2),
		.in_wire_3_3(vertical_tile_14_1_to_tile_15_1_3),
		.out_wire_1_0(vertical_tile_15_1_to_tile_16_1_0),
		.out_wire_1_1(vertical_tile_15_1_to_tile_16_1_1),
		.out_wire_1_2(vertical_tile_15_1_to_tile_16_1_2),
		.out_wire_1_3(vertical_tile_15_1_to_tile_16_1_3),
		.in_wire_1_0(vertical_tile_16_1_to_tile_15_1_0),
		.in_wire_1_1(vertical_tile_16_1_to_tile_15_1_1),
		.in_wire_1_2(vertical_tile_16_1_to_tile_15_1_2),
		.in_wire_1_3(vertical_tile_16_1_to_tile_15_1_3),
		.out_wire_2_0(horizontal_tile_15_1_to_tile_15_0_0),
		.out_wire_2_1(horizontal_tile_15_1_to_tile_15_0_1),
		.out_wire_2_2(horizontal_tile_15_1_to_tile_15_0_2),
		.out_wire_2_3(horizontal_tile_15_1_to_tile_15_0_3),
		.in_wire_2_0(horizontal_tile_15_0_to_tile_15_1_0),
		.in_wire_2_1(horizontal_tile_15_0_to_tile_15_1_1),
		.in_wire_2_2(horizontal_tile_15_0_to_tile_15_1_2),
		.in_wire_2_3(horizontal_tile_15_0_to_tile_15_1_3),
		.out_wire_0_0(horizontal_tile_15_1_to_tile_15_2_0),
		.out_wire_0_1(horizontal_tile_15_1_to_tile_15_2_1),
		.out_wire_0_2(horizontal_tile_15_1_to_tile_15_2_2),
		.out_wire_0_3(horizontal_tile_15_1_to_tile_15_2_3),
		.in_wire_0_0(horizontal_tile_15_2_to_tile_15_1_0),
		.in_wire_0_1(horizontal_tile_15_2_to_tile_15_1_1),
		.in_wire_0_2(horizontal_tile_15_2_to_tile_15_1_2),
		.in_wire_0_3(horizontal_tile_15_2_to_tile_15_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(482)
	);

	pe_tile pe_tile_15_2(
		.out_wire_3_0(vertical_tile_15_2_to_tile_14_2_0),
		.out_wire_3_1(vertical_tile_15_2_to_tile_14_2_1),
		.out_wire_3_2(vertical_tile_15_2_to_tile_14_2_2),
		.out_wire_3_3(vertical_tile_15_2_to_tile_14_2_3),
		.in_wire_3_0(vertical_tile_14_2_to_tile_15_2_0),
		.in_wire_3_1(vertical_tile_14_2_to_tile_15_2_1),
		.in_wire_3_2(vertical_tile_14_2_to_tile_15_2_2),
		.in_wire_3_3(vertical_tile_14_2_to_tile_15_2_3),
		.out_wire_1_0(vertical_tile_15_2_to_tile_16_2_0),
		.out_wire_1_1(vertical_tile_15_2_to_tile_16_2_1),
		.out_wire_1_2(vertical_tile_15_2_to_tile_16_2_2),
		.out_wire_1_3(vertical_tile_15_2_to_tile_16_2_3),
		.in_wire_1_0(vertical_tile_16_2_to_tile_15_2_0),
		.in_wire_1_1(vertical_tile_16_2_to_tile_15_2_1),
		.in_wire_1_2(vertical_tile_16_2_to_tile_15_2_2),
		.in_wire_1_3(vertical_tile_16_2_to_tile_15_2_3),
		.out_wire_2_0(horizontal_tile_15_2_to_tile_15_1_0),
		.out_wire_2_1(horizontal_tile_15_2_to_tile_15_1_1),
		.out_wire_2_2(horizontal_tile_15_2_to_tile_15_1_2),
		.out_wire_2_3(horizontal_tile_15_2_to_tile_15_1_3),
		.in_wire_2_0(horizontal_tile_15_1_to_tile_15_2_0),
		.in_wire_2_1(horizontal_tile_15_1_to_tile_15_2_1),
		.in_wire_2_2(horizontal_tile_15_1_to_tile_15_2_2),
		.in_wire_2_3(horizontal_tile_15_1_to_tile_15_2_3),
		.out_wire_0_0(horizontal_tile_15_2_to_tile_15_3_0),
		.out_wire_0_1(horizontal_tile_15_2_to_tile_15_3_1),
		.out_wire_0_2(horizontal_tile_15_2_to_tile_15_3_2),
		.out_wire_0_3(horizontal_tile_15_2_to_tile_15_3_3),
		.in_wire_0_0(horizontal_tile_15_3_to_tile_15_2_0),
		.in_wire_0_1(horizontal_tile_15_3_to_tile_15_2_1),
		.in_wire_0_2(horizontal_tile_15_3_to_tile_15_2_2),
		.in_wire_0_3(horizontal_tile_15_3_to_tile_15_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(483)
	);

	pe_tile pe_tile_15_3(
		.out_wire_3_0(vertical_tile_15_3_to_tile_14_3_0),
		.out_wire_3_1(vertical_tile_15_3_to_tile_14_3_1),
		.out_wire_3_2(vertical_tile_15_3_to_tile_14_3_2),
		.out_wire_3_3(vertical_tile_15_3_to_tile_14_3_3),
		.in_wire_3_0(vertical_tile_14_3_to_tile_15_3_0),
		.in_wire_3_1(vertical_tile_14_3_to_tile_15_3_1),
		.in_wire_3_2(vertical_tile_14_3_to_tile_15_3_2),
		.in_wire_3_3(vertical_tile_14_3_to_tile_15_3_3),
		.out_wire_1_0(vertical_tile_15_3_to_tile_16_3_0),
		.out_wire_1_1(vertical_tile_15_3_to_tile_16_3_1),
		.out_wire_1_2(vertical_tile_15_3_to_tile_16_3_2),
		.out_wire_1_3(vertical_tile_15_3_to_tile_16_3_3),
		.in_wire_1_0(vertical_tile_16_3_to_tile_15_3_0),
		.in_wire_1_1(vertical_tile_16_3_to_tile_15_3_1),
		.in_wire_1_2(vertical_tile_16_3_to_tile_15_3_2),
		.in_wire_1_3(vertical_tile_16_3_to_tile_15_3_3),
		.out_wire_2_0(horizontal_tile_15_3_to_tile_15_2_0),
		.out_wire_2_1(horizontal_tile_15_3_to_tile_15_2_1),
		.out_wire_2_2(horizontal_tile_15_3_to_tile_15_2_2),
		.out_wire_2_3(horizontal_tile_15_3_to_tile_15_2_3),
		.in_wire_2_0(horizontal_tile_15_2_to_tile_15_3_0),
		.in_wire_2_1(horizontal_tile_15_2_to_tile_15_3_1),
		.in_wire_2_2(horizontal_tile_15_2_to_tile_15_3_2),
		.in_wire_2_3(horizontal_tile_15_2_to_tile_15_3_3),
		.out_wire_0_0(horizontal_tile_15_3_to_tile_15_4_0),
		.out_wire_0_1(horizontal_tile_15_3_to_tile_15_4_1),
		.out_wire_0_2(horizontal_tile_15_3_to_tile_15_4_2),
		.out_wire_0_3(horizontal_tile_15_3_to_tile_15_4_3),
		.in_wire_0_0(horizontal_tile_15_4_to_tile_15_3_0),
		.in_wire_0_1(horizontal_tile_15_4_to_tile_15_3_1),
		.in_wire_0_2(horizontal_tile_15_4_to_tile_15_3_2),
		.in_wire_0_3(horizontal_tile_15_4_to_tile_15_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(484)
	);

	pe_tile pe_tile_15_4(
		.out_wire_3_0(vertical_tile_15_4_to_tile_14_4_0),
		.out_wire_3_1(vertical_tile_15_4_to_tile_14_4_1),
		.out_wire_3_2(vertical_tile_15_4_to_tile_14_4_2),
		.out_wire_3_3(vertical_tile_15_4_to_tile_14_4_3),
		.in_wire_3_0(vertical_tile_14_4_to_tile_15_4_0),
		.in_wire_3_1(vertical_tile_14_4_to_tile_15_4_1),
		.in_wire_3_2(vertical_tile_14_4_to_tile_15_4_2),
		.in_wire_3_3(vertical_tile_14_4_to_tile_15_4_3),
		.out_wire_1_0(vertical_tile_15_4_to_tile_16_4_0),
		.out_wire_1_1(vertical_tile_15_4_to_tile_16_4_1),
		.out_wire_1_2(vertical_tile_15_4_to_tile_16_4_2),
		.out_wire_1_3(vertical_tile_15_4_to_tile_16_4_3),
		.in_wire_1_0(vertical_tile_16_4_to_tile_15_4_0),
		.in_wire_1_1(vertical_tile_16_4_to_tile_15_4_1),
		.in_wire_1_2(vertical_tile_16_4_to_tile_15_4_2),
		.in_wire_1_3(vertical_tile_16_4_to_tile_15_4_3),
		.out_wire_2_0(horizontal_tile_15_4_to_tile_15_3_0),
		.out_wire_2_1(horizontal_tile_15_4_to_tile_15_3_1),
		.out_wire_2_2(horizontal_tile_15_4_to_tile_15_3_2),
		.out_wire_2_3(horizontal_tile_15_4_to_tile_15_3_3),
		.in_wire_2_0(horizontal_tile_15_3_to_tile_15_4_0),
		.in_wire_2_1(horizontal_tile_15_3_to_tile_15_4_1),
		.in_wire_2_2(horizontal_tile_15_3_to_tile_15_4_2),
		.in_wire_2_3(horizontal_tile_15_3_to_tile_15_4_3),
		.out_wire_0_0(horizontal_tile_15_4_to_tile_15_5_0),
		.out_wire_0_1(horizontal_tile_15_4_to_tile_15_5_1),
		.out_wire_0_2(horizontal_tile_15_4_to_tile_15_5_2),
		.out_wire_0_3(horizontal_tile_15_4_to_tile_15_5_3),
		.in_wire_0_0(horizontal_tile_15_5_to_tile_15_4_0),
		.in_wire_0_1(horizontal_tile_15_5_to_tile_15_4_1),
		.in_wire_0_2(horizontal_tile_15_5_to_tile_15_4_2),
		.in_wire_0_3(horizontal_tile_15_5_to_tile_15_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(485)
	);

	pe_tile pe_tile_15_5(
		.out_wire_3_0(vertical_tile_15_5_to_tile_14_5_0),
		.out_wire_3_1(vertical_tile_15_5_to_tile_14_5_1),
		.out_wire_3_2(vertical_tile_15_5_to_tile_14_5_2),
		.out_wire_3_3(vertical_tile_15_5_to_tile_14_5_3),
		.in_wire_3_0(vertical_tile_14_5_to_tile_15_5_0),
		.in_wire_3_1(vertical_tile_14_5_to_tile_15_5_1),
		.in_wire_3_2(vertical_tile_14_5_to_tile_15_5_2),
		.in_wire_3_3(vertical_tile_14_5_to_tile_15_5_3),
		.out_wire_1_0(vertical_tile_15_5_to_tile_16_5_0),
		.out_wire_1_1(vertical_tile_15_5_to_tile_16_5_1),
		.out_wire_1_2(vertical_tile_15_5_to_tile_16_5_2),
		.out_wire_1_3(vertical_tile_15_5_to_tile_16_5_3),
		.in_wire_1_0(vertical_tile_16_5_to_tile_15_5_0),
		.in_wire_1_1(vertical_tile_16_5_to_tile_15_5_1),
		.in_wire_1_2(vertical_tile_16_5_to_tile_15_5_2),
		.in_wire_1_3(vertical_tile_16_5_to_tile_15_5_3),
		.out_wire_2_0(horizontal_tile_15_5_to_tile_15_4_0),
		.out_wire_2_1(horizontal_tile_15_5_to_tile_15_4_1),
		.out_wire_2_2(horizontal_tile_15_5_to_tile_15_4_2),
		.out_wire_2_3(horizontal_tile_15_5_to_tile_15_4_3),
		.in_wire_2_0(horizontal_tile_15_4_to_tile_15_5_0),
		.in_wire_2_1(horizontal_tile_15_4_to_tile_15_5_1),
		.in_wire_2_2(horizontal_tile_15_4_to_tile_15_5_2),
		.in_wire_2_3(horizontal_tile_15_4_to_tile_15_5_3),
		.out_wire_0_0(horizontal_tile_15_5_to_tile_15_6_0),
		.out_wire_0_1(horizontal_tile_15_5_to_tile_15_6_1),
		.out_wire_0_2(horizontal_tile_15_5_to_tile_15_6_2),
		.out_wire_0_3(horizontal_tile_15_5_to_tile_15_6_3),
		.in_wire_0_0(horizontal_tile_15_6_to_tile_15_5_0),
		.in_wire_0_1(horizontal_tile_15_6_to_tile_15_5_1),
		.in_wire_0_2(horizontal_tile_15_6_to_tile_15_5_2),
		.in_wire_0_3(horizontal_tile_15_6_to_tile_15_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(486)
	);

	pe_tile pe_tile_15_6(
		.out_wire_3_0(vertical_tile_15_6_to_tile_14_6_0),
		.out_wire_3_1(vertical_tile_15_6_to_tile_14_6_1),
		.out_wire_3_2(vertical_tile_15_6_to_tile_14_6_2),
		.out_wire_3_3(vertical_tile_15_6_to_tile_14_6_3),
		.in_wire_3_0(vertical_tile_14_6_to_tile_15_6_0),
		.in_wire_3_1(vertical_tile_14_6_to_tile_15_6_1),
		.in_wire_3_2(vertical_tile_14_6_to_tile_15_6_2),
		.in_wire_3_3(vertical_tile_14_6_to_tile_15_6_3),
		.out_wire_1_0(vertical_tile_15_6_to_tile_16_6_0),
		.out_wire_1_1(vertical_tile_15_6_to_tile_16_6_1),
		.out_wire_1_2(vertical_tile_15_6_to_tile_16_6_2),
		.out_wire_1_3(vertical_tile_15_6_to_tile_16_6_3),
		.in_wire_1_0(vertical_tile_16_6_to_tile_15_6_0),
		.in_wire_1_1(vertical_tile_16_6_to_tile_15_6_1),
		.in_wire_1_2(vertical_tile_16_6_to_tile_15_6_2),
		.in_wire_1_3(vertical_tile_16_6_to_tile_15_6_3),
		.out_wire_2_0(horizontal_tile_15_6_to_tile_15_5_0),
		.out_wire_2_1(horizontal_tile_15_6_to_tile_15_5_1),
		.out_wire_2_2(horizontal_tile_15_6_to_tile_15_5_2),
		.out_wire_2_3(horizontal_tile_15_6_to_tile_15_5_3),
		.in_wire_2_0(horizontal_tile_15_5_to_tile_15_6_0),
		.in_wire_2_1(horizontal_tile_15_5_to_tile_15_6_1),
		.in_wire_2_2(horizontal_tile_15_5_to_tile_15_6_2),
		.in_wire_2_3(horizontal_tile_15_5_to_tile_15_6_3),
		.out_wire_0_0(horizontal_tile_15_6_to_tile_15_7_0),
		.out_wire_0_1(horizontal_tile_15_6_to_tile_15_7_1),
		.out_wire_0_2(horizontal_tile_15_6_to_tile_15_7_2),
		.out_wire_0_3(horizontal_tile_15_6_to_tile_15_7_3),
		.in_wire_0_0(horizontal_tile_15_7_to_tile_15_6_0),
		.in_wire_0_1(horizontal_tile_15_7_to_tile_15_6_1),
		.in_wire_0_2(horizontal_tile_15_7_to_tile_15_6_2),
		.in_wire_0_3(horizontal_tile_15_7_to_tile_15_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(487)
	);

	pe_tile pe_tile_15_7(
		.out_wire_3_0(vertical_tile_15_7_to_tile_14_7_0),
		.out_wire_3_1(vertical_tile_15_7_to_tile_14_7_1),
		.out_wire_3_2(vertical_tile_15_7_to_tile_14_7_2),
		.out_wire_3_3(vertical_tile_15_7_to_tile_14_7_3),
		.in_wire_3_0(vertical_tile_14_7_to_tile_15_7_0),
		.in_wire_3_1(vertical_tile_14_7_to_tile_15_7_1),
		.in_wire_3_2(vertical_tile_14_7_to_tile_15_7_2),
		.in_wire_3_3(vertical_tile_14_7_to_tile_15_7_3),
		.out_wire_1_0(vertical_tile_15_7_to_tile_16_7_0),
		.out_wire_1_1(vertical_tile_15_7_to_tile_16_7_1),
		.out_wire_1_2(vertical_tile_15_7_to_tile_16_7_2),
		.out_wire_1_3(vertical_tile_15_7_to_tile_16_7_3),
		.in_wire_1_0(vertical_tile_16_7_to_tile_15_7_0),
		.in_wire_1_1(vertical_tile_16_7_to_tile_15_7_1),
		.in_wire_1_2(vertical_tile_16_7_to_tile_15_7_2),
		.in_wire_1_3(vertical_tile_16_7_to_tile_15_7_3),
		.out_wire_2_0(horizontal_tile_15_7_to_tile_15_6_0),
		.out_wire_2_1(horizontal_tile_15_7_to_tile_15_6_1),
		.out_wire_2_2(horizontal_tile_15_7_to_tile_15_6_2),
		.out_wire_2_3(horizontal_tile_15_7_to_tile_15_6_3),
		.in_wire_2_0(horizontal_tile_15_6_to_tile_15_7_0),
		.in_wire_2_1(horizontal_tile_15_6_to_tile_15_7_1),
		.in_wire_2_2(horizontal_tile_15_6_to_tile_15_7_2),
		.in_wire_2_3(horizontal_tile_15_6_to_tile_15_7_3),
		.out_wire_0_0(horizontal_tile_15_7_to_tile_15_8_0),
		.out_wire_0_1(horizontal_tile_15_7_to_tile_15_8_1),
		.out_wire_0_2(horizontal_tile_15_7_to_tile_15_8_2),
		.out_wire_0_3(horizontal_tile_15_7_to_tile_15_8_3),
		.in_wire_0_0(horizontal_tile_15_8_to_tile_15_7_0),
		.in_wire_0_1(horizontal_tile_15_8_to_tile_15_7_1),
		.in_wire_0_2(horizontal_tile_15_8_to_tile_15_7_2),
		.in_wire_0_3(horizontal_tile_15_8_to_tile_15_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(488)
	);

	pe_tile pe_tile_15_8(
		.out_wire_3_0(vertical_tile_15_8_to_tile_14_8_0),
		.out_wire_3_1(vertical_tile_15_8_to_tile_14_8_1),
		.out_wire_3_2(vertical_tile_15_8_to_tile_14_8_2),
		.out_wire_3_3(vertical_tile_15_8_to_tile_14_8_3),
		.in_wire_3_0(vertical_tile_14_8_to_tile_15_8_0),
		.in_wire_3_1(vertical_tile_14_8_to_tile_15_8_1),
		.in_wire_3_2(vertical_tile_14_8_to_tile_15_8_2),
		.in_wire_3_3(vertical_tile_14_8_to_tile_15_8_3),
		.out_wire_1_0(vertical_tile_15_8_to_tile_16_8_0),
		.out_wire_1_1(vertical_tile_15_8_to_tile_16_8_1),
		.out_wire_1_2(vertical_tile_15_8_to_tile_16_8_2),
		.out_wire_1_3(vertical_tile_15_8_to_tile_16_8_3),
		.in_wire_1_0(vertical_tile_16_8_to_tile_15_8_0),
		.in_wire_1_1(vertical_tile_16_8_to_tile_15_8_1),
		.in_wire_1_2(vertical_tile_16_8_to_tile_15_8_2),
		.in_wire_1_3(vertical_tile_16_8_to_tile_15_8_3),
		.out_wire_2_0(horizontal_tile_15_8_to_tile_15_7_0),
		.out_wire_2_1(horizontal_tile_15_8_to_tile_15_7_1),
		.out_wire_2_2(horizontal_tile_15_8_to_tile_15_7_2),
		.out_wire_2_3(horizontal_tile_15_8_to_tile_15_7_3),
		.in_wire_2_0(horizontal_tile_15_7_to_tile_15_8_0),
		.in_wire_2_1(horizontal_tile_15_7_to_tile_15_8_1),
		.in_wire_2_2(horizontal_tile_15_7_to_tile_15_8_2),
		.in_wire_2_3(horizontal_tile_15_7_to_tile_15_8_3),
		.out_wire_0_0(horizontal_tile_15_8_to_tile_15_9_0),
		.out_wire_0_1(horizontal_tile_15_8_to_tile_15_9_1),
		.out_wire_0_2(horizontal_tile_15_8_to_tile_15_9_2),
		.out_wire_0_3(horizontal_tile_15_8_to_tile_15_9_3),
		.in_wire_0_0(horizontal_tile_15_9_to_tile_15_8_0),
		.in_wire_0_1(horizontal_tile_15_9_to_tile_15_8_1),
		.in_wire_0_2(horizontal_tile_15_9_to_tile_15_8_2),
		.in_wire_0_3(horizontal_tile_15_9_to_tile_15_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(489)
	);

	pe_tile pe_tile_15_9(
		.out_wire_3_0(vertical_tile_15_9_to_tile_14_9_0),
		.out_wire_3_1(vertical_tile_15_9_to_tile_14_9_1),
		.out_wire_3_2(vertical_tile_15_9_to_tile_14_9_2),
		.out_wire_3_3(vertical_tile_15_9_to_tile_14_9_3),
		.in_wire_3_0(vertical_tile_14_9_to_tile_15_9_0),
		.in_wire_3_1(vertical_tile_14_9_to_tile_15_9_1),
		.in_wire_3_2(vertical_tile_14_9_to_tile_15_9_2),
		.in_wire_3_3(vertical_tile_14_9_to_tile_15_9_3),
		.out_wire_1_0(vertical_tile_15_9_to_tile_16_9_0),
		.out_wire_1_1(vertical_tile_15_9_to_tile_16_9_1),
		.out_wire_1_2(vertical_tile_15_9_to_tile_16_9_2),
		.out_wire_1_3(vertical_tile_15_9_to_tile_16_9_3),
		.in_wire_1_0(vertical_tile_16_9_to_tile_15_9_0),
		.in_wire_1_1(vertical_tile_16_9_to_tile_15_9_1),
		.in_wire_1_2(vertical_tile_16_9_to_tile_15_9_2),
		.in_wire_1_3(vertical_tile_16_9_to_tile_15_9_3),
		.out_wire_2_0(horizontal_tile_15_9_to_tile_15_8_0),
		.out_wire_2_1(horizontal_tile_15_9_to_tile_15_8_1),
		.out_wire_2_2(horizontal_tile_15_9_to_tile_15_8_2),
		.out_wire_2_3(horizontal_tile_15_9_to_tile_15_8_3),
		.in_wire_2_0(horizontal_tile_15_8_to_tile_15_9_0),
		.in_wire_2_1(horizontal_tile_15_8_to_tile_15_9_1),
		.in_wire_2_2(horizontal_tile_15_8_to_tile_15_9_2),
		.in_wire_2_3(horizontal_tile_15_8_to_tile_15_9_3),
		.out_wire_0_0(horizontal_tile_15_9_to_tile_15_10_0),
		.out_wire_0_1(horizontal_tile_15_9_to_tile_15_10_1),
		.out_wire_0_2(horizontal_tile_15_9_to_tile_15_10_2),
		.out_wire_0_3(horizontal_tile_15_9_to_tile_15_10_3),
		.in_wire_0_0(horizontal_tile_15_10_to_tile_15_9_0),
		.in_wire_0_1(horizontal_tile_15_10_to_tile_15_9_1),
		.in_wire_0_2(horizontal_tile_15_10_to_tile_15_9_2),
		.in_wire_0_3(horizontal_tile_15_10_to_tile_15_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(490)
	);

	pe_tile pe_tile_15_10(
		.out_wire_3_0(vertical_tile_15_10_to_tile_14_10_0),
		.out_wire_3_1(vertical_tile_15_10_to_tile_14_10_1),
		.out_wire_3_2(vertical_tile_15_10_to_tile_14_10_2),
		.out_wire_3_3(vertical_tile_15_10_to_tile_14_10_3),
		.in_wire_3_0(vertical_tile_14_10_to_tile_15_10_0),
		.in_wire_3_1(vertical_tile_14_10_to_tile_15_10_1),
		.in_wire_3_2(vertical_tile_14_10_to_tile_15_10_2),
		.in_wire_3_3(vertical_tile_14_10_to_tile_15_10_3),
		.out_wire_1_0(vertical_tile_15_10_to_tile_16_10_0),
		.out_wire_1_1(vertical_tile_15_10_to_tile_16_10_1),
		.out_wire_1_2(vertical_tile_15_10_to_tile_16_10_2),
		.out_wire_1_3(vertical_tile_15_10_to_tile_16_10_3),
		.in_wire_1_0(vertical_tile_16_10_to_tile_15_10_0),
		.in_wire_1_1(vertical_tile_16_10_to_tile_15_10_1),
		.in_wire_1_2(vertical_tile_16_10_to_tile_15_10_2),
		.in_wire_1_3(vertical_tile_16_10_to_tile_15_10_3),
		.out_wire_2_0(horizontal_tile_15_10_to_tile_15_9_0),
		.out_wire_2_1(horizontal_tile_15_10_to_tile_15_9_1),
		.out_wire_2_2(horizontal_tile_15_10_to_tile_15_9_2),
		.out_wire_2_3(horizontal_tile_15_10_to_tile_15_9_3),
		.in_wire_2_0(horizontal_tile_15_9_to_tile_15_10_0),
		.in_wire_2_1(horizontal_tile_15_9_to_tile_15_10_1),
		.in_wire_2_2(horizontal_tile_15_9_to_tile_15_10_2),
		.in_wire_2_3(horizontal_tile_15_9_to_tile_15_10_3),
		.out_wire_0_0(horizontal_tile_15_10_to_tile_15_11_0),
		.out_wire_0_1(horizontal_tile_15_10_to_tile_15_11_1),
		.out_wire_0_2(horizontal_tile_15_10_to_tile_15_11_2),
		.out_wire_0_3(horizontal_tile_15_10_to_tile_15_11_3),
		.in_wire_0_0(horizontal_tile_15_11_to_tile_15_10_0),
		.in_wire_0_1(horizontal_tile_15_11_to_tile_15_10_1),
		.in_wire_0_2(horizontal_tile_15_11_to_tile_15_10_2),
		.in_wire_0_3(horizontal_tile_15_11_to_tile_15_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(491)
	);

	pe_tile pe_tile_15_11(
		.out_wire_3_0(vertical_tile_15_11_to_tile_14_11_0),
		.out_wire_3_1(vertical_tile_15_11_to_tile_14_11_1),
		.out_wire_3_2(vertical_tile_15_11_to_tile_14_11_2),
		.out_wire_3_3(vertical_tile_15_11_to_tile_14_11_3),
		.in_wire_3_0(vertical_tile_14_11_to_tile_15_11_0),
		.in_wire_3_1(vertical_tile_14_11_to_tile_15_11_1),
		.in_wire_3_2(vertical_tile_14_11_to_tile_15_11_2),
		.in_wire_3_3(vertical_tile_14_11_to_tile_15_11_3),
		.out_wire_1_0(vertical_tile_15_11_to_tile_16_11_0),
		.out_wire_1_1(vertical_tile_15_11_to_tile_16_11_1),
		.out_wire_1_2(vertical_tile_15_11_to_tile_16_11_2),
		.out_wire_1_3(vertical_tile_15_11_to_tile_16_11_3),
		.in_wire_1_0(vertical_tile_16_11_to_tile_15_11_0),
		.in_wire_1_1(vertical_tile_16_11_to_tile_15_11_1),
		.in_wire_1_2(vertical_tile_16_11_to_tile_15_11_2),
		.in_wire_1_3(vertical_tile_16_11_to_tile_15_11_3),
		.out_wire_2_0(horizontal_tile_15_11_to_tile_15_10_0),
		.out_wire_2_1(horizontal_tile_15_11_to_tile_15_10_1),
		.out_wire_2_2(horizontal_tile_15_11_to_tile_15_10_2),
		.out_wire_2_3(horizontal_tile_15_11_to_tile_15_10_3),
		.in_wire_2_0(horizontal_tile_15_10_to_tile_15_11_0),
		.in_wire_2_1(horizontal_tile_15_10_to_tile_15_11_1),
		.in_wire_2_2(horizontal_tile_15_10_to_tile_15_11_2),
		.in_wire_2_3(horizontal_tile_15_10_to_tile_15_11_3),
		.out_wire_0_0(horizontal_tile_15_11_to_tile_15_12_0),
		.out_wire_0_1(horizontal_tile_15_11_to_tile_15_12_1),
		.out_wire_0_2(horizontal_tile_15_11_to_tile_15_12_2),
		.out_wire_0_3(horizontal_tile_15_11_to_tile_15_12_3),
		.in_wire_0_0(horizontal_tile_15_12_to_tile_15_11_0),
		.in_wire_0_1(horizontal_tile_15_12_to_tile_15_11_1),
		.in_wire_0_2(horizontal_tile_15_12_to_tile_15_11_2),
		.in_wire_0_3(horizontal_tile_15_12_to_tile_15_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(492)
	);

	pe_tile pe_tile_15_12(
		.out_wire_3_0(vertical_tile_15_12_to_tile_14_12_0),
		.out_wire_3_1(vertical_tile_15_12_to_tile_14_12_1),
		.out_wire_3_2(vertical_tile_15_12_to_tile_14_12_2),
		.out_wire_3_3(vertical_tile_15_12_to_tile_14_12_3),
		.in_wire_3_0(vertical_tile_14_12_to_tile_15_12_0),
		.in_wire_3_1(vertical_tile_14_12_to_tile_15_12_1),
		.in_wire_3_2(vertical_tile_14_12_to_tile_15_12_2),
		.in_wire_3_3(vertical_tile_14_12_to_tile_15_12_3),
		.out_wire_1_0(vertical_tile_15_12_to_tile_16_12_0),
		.out_wire_1_1(vertical_tile_15_12_to_tile_16_12_1),
		.out_wire_1_2(vertical_tile_15_12_to_tile_16_12_2),
		.out_wire_1_3(vertical_tile_15_12_to_tile_16_12_3),
		.in_wire_1_0(vertical_tile_16_12_to_tile_15_12_0),
		.in_wire_1_1(vertical_tile_16_12_to_tile_15_12_1),
		.in_wire_1_2(vertical_tile_16_12_to_tile_15_12_2),
		.in_wire_1_3(vertical_tile_16_12_to_tile_15_12_3),
		.out_wire_2_0(horizontal_tile_15_12_to_tile_15_11_0),
		.out_wire_2_1(horizontal_tile_15_12_to_tile_15_11_1),
		.out_wire_2_2(horizontal_tile_15_12_to_tile_15_11_2),
		.out_wire_2_3(horizontal_tile_15_12_to_tile_15_11_3),
		.in_wire_2_0(horizontal_tile_15_11_to_tile_15_12_0),
		.in_wire_2_1(horizontal_tile_15_11_to_tile_15_12_1),
		.in_wire_2_2(horizontal_tile_15_11_to_tile_15_12_2),
		.in_wire_2_3(horizontal_tile_15_11_to_tile_15_12_3),
		.out_wire_0_0(horizontal_tile_15_12_to_tile_15_13_0),
		.out_wire_0_1(horizontal_tile_15_12_to_tile_15_13_1),
		.out_wire_0_2(horizontal_tile_15_12_to_tile_15_13_2),
		.out_wire_0_3(horizontal_tile_15_12_to_tile_15_13_3),
		.in_wire_0_0(horizontal_tile_15_13_to_tile_15_12_0),
		.in_wire_0_1(horizontal_tile_15_13_to_tile_15_12_1),
		.in_wire_0_2(horizontal_tile_15_13_to_tile_15_12_2),
		.in_wire_0_3(horizontal_tile_15_13_to_tile_15_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(493)
	);

	pe_tile pe_tile_15_13(
		.out_wire_3_0(vertical_tile_15_13_to_tile_14_13_0),
		.out_wire_3_1(vertical_tile_15_13_to_tile_14_13_1),
		.out_wire_3_2(vertical_tile_15_13_to_tile_14_13_2),
		.out_wire_3_3(vertical_tile_15_13_to_tile_14_13_3),
		.in_wire_3_0(vertical_tile_14_13_to_tile_15_13_0),
		.in_wire_3_1(vertical_tile_14_13_to_tile_15_13_1),
		.in_wire_3_2(vertical_tile_14_13_to_tile_15_13_2),
		.in_wire_3_3(vertical_tile_14_13_to_tile_15_13_3),
		.out_wire_1_0(vertical_tile_15_13_to_tile_16_13_0),
		.out_wire_1_1(vertical_tile_15_13_to_tile_16_13_1),
		.out_wire_1_2(vertical_tile_15_13_to_tile_16_13_2),
		.out_wire_1_3(vertical_tile_15_13_to_tile_16_13_3),
		.in_wire_1_0(vertical_tile_16_13_to_tile_15_13_0),
		.in_wire_1_1(vertical_tile_16_13_to_tile_15_13_1),
		.in_wire_1_2(vertical_tile_16_13_to_tile_15_13_2),
		.in_wire_1_3(vertical_tile_16_13_to_tile_15_13_3),
		.out_wire_2_0(horizontal_tile_15_13_to_tile_15_12_0),
		.out_wire_2_1(horizontal_tile_15_13_to_tile_15_12_1),
		.out_wire_2_2(horizontal_tile_15_13_to_tile_15_12_2),
		.out_wire_2_3(horizontal_tile_15_13_to_tile_15_12_3),
		.in_wire_2_0(horizontal_tile_15_12_to_tile_15_13_0),
		.in_wire_2_1(horizontal_tile_15_12_to_tile_15_13_1),
		.in_wire_2_2(horizontal_tile_15_12_to_tile_15_13_2),
		.in_wire_2_3(horizontal_tile_15_12_to_tile_15_13_3),
		.out_wire_0_0(horizontal_tile_15_13_to_tile_15_14_0),
		.out_wire_0_1(horizontal_tile_15_13_to_tile_15_14_1),
		.out_wire_0_2(horizontal_tile_15_13_to_tile_15_14_2),
		.out_wire_0_3(horizontal_tile_15_13_to_tile_15_14_3),
		.in_wire_0_0(horizontal_tile_15_14_to_tile_15_13_0),
		.in_wire_0_1(horizontal_tile_15_14_to_tile_15_13_1),
		.in_wire_0_2(horizontal_tile_15_14_to_tile_15_13_2),
		.in_wire_0_3(horizontal_tile_15_14_to_tile_15_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(494)
	);

	pe_tile pe_tile_15_14(
		.out_wire_3_0(vertical_tile_15_14_to_tile_14_14_0),
		.out_wire_3_1(vertical_tile_15_14_to_tile_14_14_1),
		.out_wire_3_2(vertical_tile_15_14_to_tile_14_14_2),
		.out_wire_3_3(vertical_tile_15_14_to_tile_14_14_3),
		.in_wire_3_0(vertical_tile_14_14_to_tile_15_14_0),
		.in_wire_3_1(vertical_tile_14_14_to_tile_15_14_1),
		.in_wire_3_2(vertical_tile_14_14_to_tile_15_14_2),
		.in_wire_3_3(vertical_tile_14_14_to_tile_15_14_3),
		.out_wire_1_0(vertical_tile_15_14_to_tile_16_14_0),
		.out_wire_1_1(vertical_tile_15_14_to_tile_16_14_1),
		.out_wire_1_2(vertical_tile_15_14_to_tile_16_14_2),
		.out_wire_1_3(vertical_tile_15_14_to_tile_16_14_3),
		.in_wire_1_0(vertical_tile_16_14_to_tile_15_14_0),
		.in_wire_1_1(vertical_tile_16_14_to_tile_15_14_1),
		.in_wire_1_2(vertical_tile_16_14_to_tile_15_14_2),
		.in_wire_1_3(vertical_tile_16_14_to_tile_15_14_3),
		.out_wire_2_0(horizontal_tile_15_14_to_tile_15_13_0),
		.out_wire_2_1(horizontal_tile_15_14_to_tile_15_13_1),
		.out_wire_2_2(horizontal_tile_15_14_to_tile_15_13_2),
		.out_wire_2_3(horizontal_tile_15_14_to_tile_15_13_3),
		.in_wire_2_0(horizontal_tile_15_13_to_tile_15_14_0),
		.in_wire_2_1(horizontal_tile_15_13_to_tile_15_14_1),
		.in_wire_2_2(horizontal_tile_15_13_to_tile_15_14_2),
		.in_wire_2_3(horizontal_tile_15_13_to_tile_15_14_3),
		.out_wire_0_0(horizontal_tile_15_14_to_tile_15_15_0),
		.out_wire_0_1(horizontal_tile_15_14_to_tile_15_15_1),
		.out_wire_0_2(horizontal_tile_15_14_to_tile_15_15_2),
		.out_wire_0_3(horizontal_tile_15_14_to_tile_15_15_3),
		.in_wire_0_0(horizontal_tile_15_15_to_tile_15_14_0),
		.in_wire_0_1(horizontal_tile_15_15_to_tile_15_14_1),
		.in_wire_0_2(horizontal_tile_15_15_to_tile_15_14_2),
		.in_wire_0_3(horizontal_tile_15_15_to_tile_15_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(495)
	);

	pe_tile pe_tile_15_15(
		.out_wire_3_0(vertical_tile_15_15_to_tile_14_15_0),
		.out_wire_3_1(vertical_tile_15_15_to_tile_14_15_1),
		.out_wire_3_2(vertical_tile_15_15_to_tile_14_15_2),
		.out_wire_3_3(vertical_tile_15_15_to_tile_14_15_3),
		.in_wire_3_0(vertical_tile_14_15_to_tile_15_15_0),
		.in_wire_3_1(vertical_tile_14_15_to_tile_15_15_1),
		.in_wire_3_2(vertical_tile_14_15_to_tile_15_15_2),
		.in_wire_3_3(vertical_tile_14_15_to_tile_15_15_3),
		.out_wire_1_0(vertical_tile_15_15_to_tile_16_15_0),
		.out_wire_1_1(vertical_tile_15_15_to_tile_16_15_1),
		.out_wire_1_2(vertical_tile_15_15_to_tile_16_15_2),
		.out_wire_1_3(vertical_tile_15_15_to_tile_16_15_3),
		.in_wire_1_0(vertical_tile_16_15_to_tile_15_15_0),
		.in_wire_1_1(vertical_tile_16_15_to_tile_15_15_1),
		.in_wire_1_2(vertical_tile_16_15_to_tile_15_15_2),
		.in_wire_1_3(vertical_tile_16_15_to_tile_15_15_3),
		.out_wire_2_0(horizontal_tile_15_15_to_tile_15_14_0),
		.out_wire_2_1(horizontal_tile_15_15_to_tile_15_14_1),
		.out_wire_2_2(horizontal_tile_15_15_to_tile_15_14_2),
		.out_wire_2_3(horizontal_tile_15_15_to_tile_15_14_3),
		.in_wire_2_0(horizontal_tile_15_14_to_tile_15_15_0),
		.in_wire_2_1(horizontal_tile_15_14_to_tile_15_15_1),
		.in_wire_2_2(horizontal_tile_15_14_to_tile_15_15_2),
		.in_wire_2_3(horizontal_tile_15_14_to_tile_15_15_3),
		.out_wire_0_0(horizontal_tile_15_15_to_tile_15_16_0),
		.out_wire_0_1(horizontal_tile_15_15_to_tile_15_16_1),
		.out_wire_0_2(horizontal_tile_15_15_to_tile_15_16_2),
		.out_wire_0_3(horizontal_tile_15_15_to_tile_15_16_3),
		.in_wire_0_0(horizontal_tile_15_16_to_tile_15_15_0),
		.in_wire_0_1(horizontal_tile_15_16_to_tile_15_15_1),
		.in_wire_0_2(horizontal_tile_15_16_to_tile_15_15_2),
		.in_wire_0_3(horizontal_tile_15_16_to_tile_15_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(496)
	);

	pe_tile pe_tile_15_16(
		.out_wire_3_0(vertical_tile_15_16_to_tile_14_16_0),
		.out_wire_3_1(vertical_tile_15_16_to_tile_14_16_1),
		.out_wire_3_2(vertical_tile_15_16_to_tile_14_16_2),
		.out_wire_3_3(vertical_tile_15_16_to_tile_14_16_3),
		.in_wire_3_0(vertical_tile_14_16_to_tile_15_16_0),
		.in_wire_3_1(vertical_tile_14_16_to_tile_15_16_1),
		.in_wire_3_2(vertical_tile_14_16_to_tile_15_16_2),
		.in_wire_3_3(vertical_tile_14_16_to_tile_15_16_3),
		.out_wire_1_0(vertical_tile_15_16_to_tile_16_16_0),
		.out_wire_1_1(vertical_tile_15_16_to_tile_16_16_1),
		.out_wire_1_2(vertical_tile_15_16_to_tile_16_16_2),
		.out_wire_1_3(vertical_tile_15_16_to_tile_16_16_3),
		.in_wire_1_0(vertical_tile_16_16_to_tile_15_16_0),
		.in_wire_1_1(vertical_tile_16_16_to_tile_15_16_1),
		.in_wire_1_2(vertical_tile_16_16_to_tile_15_16_2),
		.in_wire_1_3(vertical_tile_16_16_to_tile_15_16_3),
		.out_wire_2_0(horizontal_tile_15_16_to_tile_15_15_0),
		.out_wire_2_1(horizontal_tile_15_16_to_tile_15_15_1),
		.out_wire_2_2(horizontal_tile_15_16_to_tile_15_15_2),
		.out_wire_2_3(horizontal_tile_15_16_to_tile_15_15_3),
		.in_wire_2_0(horizontal_tile_15_15_to_tile_15_16_0),
		.in_wire_2_1(horizontal_tile_15_15_to_tile_15_16_1),
		.in_wire_2_2(horizontal_tile_15_15_to_tile_15_16_2),
		.in_wire_2_3(horizontal_tile_15_15_to_tile_15_16_3),
		.out_wire_0_0(horizontal_tile_15_16_to_tile_15_17_0),
		.out_wire_0_1(horizontal_tile_15_16_to_tile_15_17_1),
		.out_wire_0_2(horizontal_tile_15_16_to_tile_15_17_2),
		.out_wire_0_3(horizontal_tile_15_16_to_tile_15_17_3),
		.in_wire_0_0(horizontal_tile_15_17_to_tile_15_16_0),
		.in_wire_0_1(horizontal_tile_15_17_to_tile_15_16_1),
		.in_wire_0_2(horizontal_tile_15_17_to_tile_15_16_2),
		.in_wire_0_3(horizontal_tile_15_17_to_tile_15_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(497)
	);

	pe_tile pe_tile_15_17(
		.out_wire_3_0(vertical_tile_15_17_to_tile_14_17_0),
		.out_wire_3_1(vertical_tile_15_17_to_tile_14_17_1),
		.out_wire_3_2(vertical_tile_15_17_to_tile_14_17_2),
		.out_wire_3_3(vertical_tile_15_17_to_tile_14_17_3),
		.in_wire_3_0(vertical_tile_14_17_to_tile_15_17_0),
		.in_wire_3_1(vertical_tile_14_17_to_tile_15_17_1),
		.in_wire_3_2(vertical_tile_14_17_to_tile_15_17_2),
		.in_wire_3_3(vertical_tile_14_17_to_tile_15_17_3),
		.out_wire_1_0(vertical_tile_15_17_to_tile_16_17_0),
		.out_wire_1_1(vertical_tile_15_17_to_tile_16_17_1),
		.out_wire_1_2(vertical_tile_15_17_to_tile_16_17_2),
		.out_wire_1_3(vertical_tile_15_17_to_tile_16_17_3),
		.in_wire_1_0(vertical_tile_16_17_to_tile_15_17_0),
		.in_wire_1_1(vertical_tile_16_17_to_tile_15_17_1),
		.in_wire_1_2(vertical_tile_16_17_to_tile_15_17_2),
		.in_wire_1_3(vertical_tile_16_17_to_tile_15_17_3),
		.out_wire_2_0(horizontal_tile_15_17_to_tile_15_16_0),
		.out_wire_2_1(horizontal_tile_15_17_to_tile_15_16_1),
		.out_wire_2_2(horizontal_tile_15_17_to_tile_15_16_2),
		.out_wire_2_3(horizontal_tile_15_17_to_tile_15_16_3),
		.in_wire_2_0(horizontal_tile_15_16_to_tile_15_17_0),
		.in_wire_2_1(horizontal_tile_15_16_to_tile_15_17_1),
		.in_wire_2_2(horizontal_tile_15_16_to_tile_15_17_2),
		.in_wire_2_3(horizontal_tile_15_16_to_tile_15_17_3),
		.out_wire_0_0(horizontal_tile_15_17_to_tile_15_18_0),
		.out_wire_0_1(horizontal_tile_15_17_to_tile_15_18_1),
		.out_wire_0_2(horizontal_tile_15_17_to_tile_15_18_2),
		.out_wire_0_3(horizontal_tile_15_17_to_tile_15_18_3),
		.in_wire_0_0(horizontal_tile_15_18_to_tile_15_17_0),
		.in_wire_0_1(horizontal_tile_15_18_to_tile_15_17_1),
		.in_wire_0_2(horizontal_tile_15_18_to_tile_15_17_2),
		.in_wire_0_3(horizontal_tile_15_18_to_tile_15_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(498)
	);

	pe_tile pe_tile_15_18(
		.out_wire_3_0(vertical_tile_15_18_to_tile_14_18_0),
		.out_wire_3_1(vertical_tile_15_18_to_tile_14_18_1),
		.out_wire_3_2(vertical_tile_15_18_to_tile_14_18_2),
		.out_wire_3_3(vertical_tile_15_18_to_tile_14_18_3),
		.in_wire_3_0(vertical_tile_14_18_to_tile_15_18_0),
		.in_wire_3_1(vertical_tile_14_18_to_tile_15_18_1),
		.in_wire_3_2(vertical_tile_14_18_to_tile_15_18_2),
		.in_wire_3_3(vertical_tile_14_18_to_tile_15_18_3),
		.out_wire_1_0(vertical_tile_15_18_to_tile_16_18_0),
		.out_wire_1_1(vertical_tile_15_18_to_tile_16_18_1),
		.out_wire_1_2(vertical_tile_15_18_to_tile_16_18_2),
		.out_wire_1_3(vertical_tile_15_18_to_tile_16_18_3),
		.in_wire_1_0(vertical_tile_16_18_to_tile_15_18_0),
		.in_wire_1_1(vertical_tile_16_18_to_tile_15_18_1),
		.in_wire_1_2(vertical_tile_16_18_to_tile_15_18_2),
		.in_wire_1_3(vertical_tile_16_18_to_tile_15_18_3),
		.out_wire_2_0(horizontal_tile_15_18_to_tile_15_17_0),
		.out_wire_2_1(horizontal_tile_15_18_to_tile_15_17_1),
		.out_wire_2_2(horizontal_tile_15_18_to_tile_15_17_2),
		.out_wire_2_3(horizontal_tile_15_18_to_tile_15_17_3),
		.in_wire_2_0(horizontal_tile_15_17_to_tile_15_18_0),
		.in_wire_2_1(horizontal_tile_15_17_to_tile_15_18_1),
		.in_wire_2_2(horizontal_tile_15_17_to_tile_15_18_2),
		.in_wire_2_3(horizontal_tile_15_17_to_tile_15_18_3),
		.out_wire_0_0(horizontal_tile_15_18_to_tile_15_19_0),
		.out_wire_0_1(horizontal_tile_15_18_to_tile_15_19_1),
		.out_wire_0_2(horizontal_tile_15_18_to_tile_15_19_2),
		.out_wire_0_3(horizontal_tile_15_18_to_tile_15_19_3),
		.in_wire_0_0(horizontal_tile_15_19_to_tile_15_18_0),
		.in_wire_0_1(horizontal_tile_15_19_to_tile_15_18_1),
		.in_wire_0_2(horizontal_tile_15_19_to_tile_15_18_2),
		.in_wire_0_3(horizontal_tile_15_19_to_tile_15_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(499)
	);

	pe_tile pe_tile_15_19(
		.out_wire_3_0(vertical_tile_15_19_to_tile_14_19_0),
		.out_wire_3_1(vertical_tile_15_19_to_tile_14_19_1),
		.out_wire_3_2(vertical_tile_15_19_to_tile_14_19_2),
		.out_wire_3_3(vertical_tile_15_19_to_tile_14_19_3),
		.in_wire_3_0(vertical_tile_14_19_to_tile_15_19_0),
		.in_wire_3_1(vertical_tile_14_19_to_tile_15_19_1),
		.in_wire_3_2(vertical_tile_14_19_to_tile_15_19_2),
		.in_wire_3_3(vertical_tile_14_19_to_tile_15_19_3),
		.out_wire_1_0(vertical_tile_15_19_to_tile_16_19_0),
		.out_wire_1_1(vertical_tile_15_19_to_tile_16_19_1),
		.out_wire_1_2(vertical_tile_15_19_to_tile_16_19_2),
		.out_wire_1_3(vertical_tile_15_19_to_tile_16_19_3),
		.in_wire_1_0(vertical_tile_16_19_to_tile_15_19_0),
		.in_wire_1_1(vertical_tile_16_19_to_tile_15_19_1),
		.in_wire_1_2(vertical_tile_16_19_to_tile_15_19_2),
		.in_wire_1_3(vertical_tile_16_19_to_tile_15_19_3),
		.out_wire_2_0(horizontal_tile_15_19_to_tile_15_18_0),
		.out_wire_2_1(horizontal_tile_15_19_to_tile_15_18_1),
		.out_wire_2_2(horizontal_tile_15_19_to_tile_15_18_2),
		.out_wire_2_3(horizontal_tile_15_19_to_tile_15_18_3),
		.in_wire_2_0(horizontal_tile_15_18_to_tile_15_19_0),
		.in_wire_2_1(horizontal_tile_15_18_to_tile_15_19_1),
		.in_wire_2_2(horizontal_tile_15_18_to_tile_15_19_2),
		.in_wire_2_3(horizontal_tile_15_18_to_tile_15_19_3),
		.out_wire_0_0(horizontal_tile_15_19_to_tile_15_20_0),
		.out_wire_0_1(horizontal_tile_15_19_to_tile_15_20_1),
		.out_wire_0_2(horizontal_tile_15_19_to_tile_15_20_2),
		.out_wire_0_3(horizontal_tile_15_19_to_tile_15_20_3),
		.in_wire_0_0(horizontal_tile_15_20_to_tile_15_19_0),
		.in_wire_0_1(horizontal_tile_15_20_to_tile_15_19_1),
		.in_wire_0_2(horizontal_tile_15_20_to_tile_15_19_2),
		.in_wire_0_3(horizontal_tile_15_20_to_tile_15_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(500)
	);

	pe_tile pe_tile_15_20(
		.out_wire_3_0(vertical_tile_15_20_to_tile_14_20_0),
		.out_wire_3_1(vertical_tile_15_20_to_tile_14_20_1),
		.out_wire_3_2(vertical_tile_15_20_to_tile_14_20_2),
		.out_wire_3_3(vertical_tile_15_20_to_tile_14_20_3),
		.in_wire_3_0(vertical_tile_14_20_to_tile_15_20_0),
		.in_wire_3_1(vertical_tile_14_20_to_tile_15_20_1),
		.in_wire_3_2(vertical_tile_14_20_to_tile_15_20_2),
		.in_wire_3_3(vertical_tile_14_20_to_tile_15_20_3),
		.out_wire_1_0(vertical_tile_15_20_to_tile_16_20_0),
		.out_wire_1_1(vertical_tile_15_20_to_tile_16_20_1),
		.out_wire_1_2(vertical_tile_15_20_to_tile_16_20_2),
		.out_wire_1_3(vertical_tile_15_20_to_tile_16_20_3),
		.in_wire_1_0(vertical_tile_16_20_to_tile_15_20_0),
		.in_wire_1_1(vertical_tile_16_20_to_tile_15_20_1),
		.in_wire_1_2(vertical_tile_16_20_to_tile_15_20_2),
		.in_wire_1_3(vertical_tile_16_20_to_tile_15_20_3),
		.out_wire_2_0(horizontal_tile_15_20_to_tile_15_19_0),
		.out_wire_2_1(horizontal_tile_15_20_to_tile_15_19_1),
		.out_wire_2_2(horizontal_tile_15_20_to_tile_15_19_2),
		.out_wire_2_3(horizontal_tile_15_20_to_tile_15_19_3),
		.in_wire_2_0(horizontal_tile_15_19_to_tile_15_20_0),
		.in_wire_2_1(horizontal_tile_15_19_to_tile_15_20_1),
		.in_wire_2_2(horizontal_tile_15_19_to_tile_15_20_2),
		.in_wire_2_3(horizontal_tile_15_19_to_tile_15_20_3),
		.out_wire_0_0(horizontal_tile_15_20_to_tile_15_21_0),
		.out_wire_0_1(horizontal_tile_15_20_to_tile_15_21_1),
		.out_wire_0_2(horizontal_tile_15_20_to_tile_15_21_2),
		.out_wire_0_3(horizontal_tile_15_20_to_tile_15_21_3),
		.in_wire_0_0(horizontal_tile_15_21_to_tile_15_20_0),
		.in_wire_0_1(horizontal_tile_15_21_to_tile_15_20_1),
		.in_wire_0_2(horizontal_tile_15_21_to_tile_15_20_2),
		.in_wire_0_3(horizontal_tile_15_21_to_tile_15_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(501)
	);

	pe_tile pe_tile_15_21(
		.out_wire_3_0(vertical_tile_15_21_to_tile_14_21_0),
		.out_wire_3_1(vertical_tile_15_21_to_tile_14_21_1),
		.out_wire_3_2(vertical_tile_15_21_to_tile_14_21_2),
		.out_wire_3_3(vertical_tile_15_21_to_tile_14_21_3),
		.in_wire_3_0(vertical_tile_14_21_to_tile_15_21_0),
		.in_wire_3_1(vertical_tile_14_21_to_tile_15_21_1),
		.in_wire_3_2(vertical_tile_14_21_to_tile_15_21_2),
		.in_wire_3_3(vertical_tile_14_21_to_tile_15_21_3),
		.out_wire_1_0(vertical_tile_15_21_to_tile_16_21_0),
		.out_wire_1_1(vertical_tile_15_21_to_tile_16_21_1),
		.out_wire_1_2(vertical_tile_15_21_to_tile_16_21_2),
		.out_wire_1_3(vertical_tile_15_21_to_tile_16_21_3),
		.in_wire_1_0(vertical_tile_16_21_to_tile_15_21_0),
		.in_wire_1_1(vertical_tile_16_21_to_tile_15_21_1),
		.in_wire_1_2(vertical_tile_16_21_to_tile_15_21_2),
		.in_wire_1_3(vertical_tile_16_21_to_tile_15_21_3),
		.out_wire_2_0(horizontal_tile_15_21_to_tile_15_20_0),
		.out_wire_2_1(horizontal_tile_15_21_to_tile_15_20_1),
		.out_wire_2_2(horizontal_tile_15_21_to_tile_15_20_2),
		.out_wire_2_3(horizontal_tile_15_21_to_tile_15_20_3),
		.in_wire_2_0(horizontal_tile_15_20_to_tile_15_21_0),
		.in_wire_2_1(horizontal_tile_15_20_to_tile_15_21_1),
		.in_wire_2_2(horizontal_tile_15_20_to_tile_15_21_2),
		.in_wire_2_3(horizontal_tile_15_20_to_tile_15_21_3),
		.out_wire_0_0(horizontal_tile_15_21_to_tile_15_22_0),
		.out_wire_0_1(horizontal_tile_15_21_to_tile_15_22_1),
		.out_wire_0_2(horizontal_tile_15_21_to_tile_15_22_2),
		.out_wire_0_3(horizontal_tile_15_21_to_tile_15_22_3),
		.in_wire_0_0(horizontal_tile_15_22_to_tile_15_21_0),
		.in_wire_0_1(horizontal_tile_15_22_to_tile_15_21_1),
		.in_wire_0_2(horizontal_tile_15_22_to_tile_15_21_2),
		.in_wire_0_3(horizontal_tile_15_22_to_tile_15_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(502)
	);

	pe_tile pe_tile_15_22(
		.out_wire_3_0(vertical_tile_15_22_to_tile_14_22_0),
		.out_wire_3_1(vertical_tile_15_22_to_tile_14_22_1),
		.out_wire_3_2(vertical_tile_15_22_to_tile_14_22_2),
		.out_wire_3_3(vertical_tile_15_22_to_tile_14_22_3),
		.in_wire_3_0(vertical_tile_14_22_to_tile_15_22_0),
		.in_wire_3_1(vertical_tile_14_22_to_tile_15_22_1),
		.in_wire_3_2(vertical_tile_14_22_to_tile_15_22_2),
		.in_wire_3_3(vertical_tile_14_22_to_tile_15_22_3),
		.out_wire_1_0(vertical_tile_15_22_to_tile_16_22_0),
		.out_wire_1_1(vertical_tile_15_22_to_tile_16_22_1),
		.out_wire_1_2(vertical_tile_15_22_to_tile_16_22_2),
		.out_wire_1_3(vertical_tile_15_22_to_tile_16_22_3),
		.in_wire_1_0(vertical_tile_16_22_to_tile_15_22_0),
		.in_wire_1_1(vertical_tile_16_22_to_tile_15_22_1),
		.in_wire_1_2(vertical_tile_16_22_to_tile_15_22_2),
		.in_wire_1_3(vertical_tile_16_22_to_tile_15_22_3),
		.out_wire_2_0(horizontal_tile_15_22_to_tile_15_21_0),
		.out_wire_2_1(horizontal_tile_15_22_to_tile_15_21_1),
		.out_wire_2_2(horizontal_tile_15_22_to_tile_15_21_2),
		.out_wire_2_3(horizontal_tile_15_22_to_tile_15_21_3),
		.in_wire_2_0(horizontal_tile_15_21_to_tile_15_22_0),
		.in_wire_2_1(horizontal_tile_15_21_to_tile_15_22_1),
		.in_wire_2_2(horizontal_tile_15_21_to_tile_15_22_2),
		.in_wire_2_3(horizontal_tile_15_21_to_tile_15_22_3),
		.out_wire_0_0(horizontal_tile_15_22_to_tile_15_23_0),
		.out_wire_0_1(horizontal_tile_15_22_to_tile_15_23_1),
		.out_wire_0_2(horizontal_tile_15_22_to_tile_15_23_2),
		.out_wire_0_3(horizontal_tile_15_22_to_tile_15_23_3),
		.in_wire_0_0(horizontal_tile_15_23_to_tile_15_22_0),
		.in_wire_0_1(horizontal_tile_15_23_to_tile_15_22_1),
		.in_wire_0_2(horizontal_tile_15_23_to_tile_15_22_2),
		.in_wire_0_3(horizontal_tile_15_23_to_tile_15_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(503)
	);

	pe_tile pe_tile_15_23(
		.out_wire_3_0(vertical_tile_15_23_to_tile_14_23_0),
		.out_wire_3_1(vertical_tile_15_23_to_tile_14_23_1),
		.out_wire_3_2(vertical_tile_15_23_to_tile_14_23_2),
		.out_wire_3_3(vertical_tile_15_23_to_tile_14_23_3),
		.in_wire_3_0(vertical_tile_14_23_to_tile_15_23_0),
		.in_wire_3_1(vertical_tile_14_23_to_tile_15_23_1),
		.in_wire_3_2(vertical_tile_14_23_to_tile_15_23_2),
		.in_wire_3_3(vertical_tile_14_23_to_tile_15_23_3),
		.out_wire_1_0(vertical_tile_15_23_to_tile_16_23_0),
		.out_wire_1_1(vertical_tile_15_23_to_tile_16_23_1),
		.out_wire_1_2(vertical_tile_15_23_to_tile_16_23_2),
		.out_wire_1_3(vertical_tile_15_23_to_tile_16_23_3),
		.in_wire_1_0(vertical_tile_16_23_to_tile_15_23_0),
		.in_wire_1_1(vertical_tile_16_23_to_tile_15_23_1),
		.in_wire_1_2(vertical_tile_16_23_to_tile_15_23_2),
		.in_wire_1_3(vertical_tile_16_23_to_tile_15_23_3),
		.out_wire_2_0(horizontal_tile_15_23_to_tile_15_22_0),
		.out_wire_2_1(horizontal_tile_15_23_to_tile_15_22_1),
		.out_wire_2_2(horizontal_tile_15_23_to_tile_15_22_2),
		.out_wire_2_3(horizontal_tile_15_23_to_tile_15_22_3),
		.in_wire_2_0(horizontal_tile_15_22_to_tile_15_23_0),
		.in_wire_2_1(horizontal_tile_15_22_to_tile_15_23_1),
		.in_wire_2_2(horizontal_tile_15_22_to_tile_15_23_2),
		.in_wire_2_3(horizontal_tile_15_22_to_tile_15_23_3),
		.out_wire_0_0(horizontal_tile_15_23_to_tile_15_24_0),
		.out_wire_0_1(horizontal_tile_15_23_to_tile_15_24_1),
		.out_wire_0_2(horizontal_tile_15_23_to_tile_15_24_2),
		.out_wire_0_3(horizontal_tile_15_23_to_tile_15_24_3),
		.in_wire_0_0(horizontal_tile_15_24_to_tile_15_23_0),
		.in_wire_0_1(horizontal_tile_15_24_to_tile_15_23_1),
		.in_wire_0_2(horizontal_tile_15_24_to_tile_15_23_2),
		.in_wire_0_3(horizontal_tile_15_24_to_tile_15_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(504)
	);

	pe_tile pe_tile_15_24(
		.out_wire_3_0(vertical_tile_15_24_to_tile_14_24_0),
		.out_wire_3_1(vertical_tile_15_24_to_tile_14_24_1),
		.out_wire_3_2(vertical_tile_15_24_to_tile_14_24_2),
		.out_wire_3_3(vertical_tile_15_24_to_tile_14_24_3),
		.in_wire_3_0(vertical_tile_14_24_to_tile_15_24_0),
		.in_wire_3_1(vertical_tile_14_24_to_tile_15_24_1),
		.in_wire_3_2(vertical_tile_14_24_to_tile_15_24_2),
		.in_wire_3_3(vertical_tile_14_24_to_tile_15_24_3),
		.out_wire_1_0(vertical_tile_15_24_to_tile_16_24_0),
		.out_wire_1_1(vertical_tile_15_24_to_tile_16_24_1),
		.out_wire_1_2(vertical_tile_15_24_to_tile_16_24_2),
		.out_wire_1_3(vertical_tile_15_24_to_tile_16_24_3),
		.in_wire_1_0(vertical_tile_16_24_to_tile_15_24_0),
		.in_wire_1_1(vertical_tile_16_24_to_tile_15_24_1),
		.in_wire_1_2(vertical_tile_16_24_to_tile_15_24_2),
		.in_wire_1_3(vertical_tile_16_24_to_tile_15_24_3),
		.out_wire_2_0(horizontal_tile_15_24_to_tile_15_23_0),
		.out_wire_2_1(horizontal_tile_15_24_to_tile_15_23_1),
		.out_wire_2_2(horizontal_tile_15_24_to_tile_15_23_2),
		.out_wire_2_3(horizontal_tile_15_24_to_tile_15_23_3),
		.in_wire_2_0(horizontal_tile_15_23_to_tile_15_24_0),
		.in_wire_2_1(horizontal_tile_15_23_to_tile_15_24_1),
		.in_wire_2_2(horizontal_tile_15_23_to_tile_15_24_2),
		.in_wire_2_3(horizontal_tile_15_23_to_tile_15_24_3),
		.out_wire_0_0(horizontal_tile_15_24_to_tile_15_25_0),
		.out_wire_0_1(horizontal_tile_15_24_to_tile_15_25_1),
		.out_wire_0_2(horizontal_tile_15_24_to_tile_15_25_2),
		.out_wire_0_3(horizontal_tile_15_24_to_tile_15_25_3),
		.in_wire_0_0(horizontal_tile_15_25_to_tile_15_24_0),
		.in_wire_0_1(horizontal_tile_15_25_to_tile_15_24_1),
		.in_wire_0_2(horizontal_tile_15_25_to_tile_15_24_2),
		.in_wire_0_3(horizontal_tile_15_25_to_tile_15_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(505)
	);

	pe_tile pe_tile_15_25(
		.out_wire_3_0(vertical_tile_15_25_to_tile_14_25_0),
		.out_wire_3_1(vertical_tile_15_25_to_tile_14_25_1),
		.out_wire_3_2(vertical_tile_15_25_to_tile_14_25_2),
		.out_wire_3_3(vertical_tile_15_25_to_tile_14_25_3),
		.in_wire_3_0(vertical_tile_14_25_to_tile_15_25_0),
		.in_wire_3_1(vertical_tile_14_25_to_tile_15_25_1),
		.in_wire_3_2(vertical_tile_14_25_to_tile_15_25_2),
		.in_wire_3_3(vertical_tile_14_25_to_tile_15_25_3),
		.out_wire_1_0(vertical_tile_15_25_to_tile_16_25_0),
		.out_wire_1_1(vertical_tile_15_25_to_tile_16_25_1),
		.out_wire_1_2(vertical_tile_15_25_to_tile_16_25_2),
		.out_wire_1_3(vertical_tile_15_25_to_tile_16_25_3),
		.in_wire_1_0(vertical_tile_16_25_to_tile_15_25_0),
		.in_wire_1_1(vertical_tile_16_25_to_tile_15_25_1),
		.in_wire_1_2(vertical_tile_16_25_to_tile_15_25_2),
		.in_wire_1_3(vertical_tile_16_25_to_tile_15_25_3),
		.out_wire_2_0(horizontal_tile_15_25_to_tile_15_24_0),
		.out_wire_2_1(horizontal_tile_15_25_to_tile_15_24_1),
		.out_wire_2_2(horizontal_tile_15_25_to_tile_15_24_2),
		.out_wire_2_3(horizontal_tile_15_25_to_tile_15_24_3),
		.in_wire_2_0(horizontal_tile_15_24_to_tile_15_25_0),
		.in_wire_2_1(horizontal_tile_15_24_to_tile_15_25_1),
		.in_wire_2_2(horizontal_tile_15_24_to_tile_15_25_2),
		.in_wire_2_3(horizontal_tile_15_24_to_tile_15_25_3),
		.out_wire_0_0(horizontal_tile_15_25_to_tile_15_26_0),
		.out_wire_0_1(horizontal_tile_15_25_to_tile_15_26_1),
		.out_wire_0_2(horizontal_tile_15_25_to_tile_15_26_2),
		.out_wire_0_3(horizontal_tile_15_25_to_tile_15_26_3),
		.in_wire_0_0(horizontal_tile_15_26_to_tile_15_25_0),
		.in_wire_0_1(horizontal_tile_15_26_to_tile_15_25_1),
		.in_wire_0_2(horizontal_tile_15_26_to_tile_15_25_2),
		.in_wire_0_3(horizontal_tile_15_26_to_tile_15_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(506)
	);

	pe_tile pe_tile_15_26(
		.out_wire_3_0(vertical_tile_15_26_to_tile_14_26_0),
		.out_wire_3_1(vertical_tile_15_26_to_tile_14_26_1),
		.out_wire_3_2(vertical_tile_15_26_to_tile_14_26_2),
		.out_wire_3_3(vertical_tile_15_26_to_tile_14_26_3),
		.in_wire_3_0(vertical_tile_14_26_to_tile_15_26_0),
		.in_wire_3_1(vertical_tile_14_26_to_tile_15_26_1),
		.in_wire_3_2(vertical_tile_14_26_to_tile_15_26_2),
		.in_wire_3_3(vertical_tile_14_26_to_tile_15_26_3),
		.out_wire_1_0(vertical_tile_15_26_to_tile_16_26_0),
		.out_wire_1_1(vertical_tile_15_26_to_tile_16_26_1),
		.out_wire_1_2(vertical_tile_15_26_to_tile_16_26_2),
		.out_wire_1_3(vertical_tile_15_26_to_tile_16_26_3),
		.in_wire_1_0(vertical_tile_16_26_to_tile_15_26_0),
		.in_wire_1_1(vertical_tile_16_26_to_tile_15_26_1),
		.in_wire_1_2(vertical_tile_16_26_to_tile_15_26_2),
		.in_wire_1_3(vertical_tile_16_26_to_tile_15_26_3),
		.out_wire_2_0(horizontal_tile_15_26_to_tile_15_25_0),
		.out_wire_2_1(horizontal_tile_15_26_to_tile_15_25_1),
		.out_wire_2_2(horizontal_tile_15_26_to_tile_15_25_2),
		.out_wire_2_3(horizontal_tile_15_26_to_tile_15_25_3),
		.in_wire_2_0(horizontal_tile_15_25_to_tile_15_26_0),
		.in_wire_2_1(horizontal_tile_15_25_to_tile_15_26_1),
		.in_wire_2_2(horizontal_tile_15_25_to_tile_15_26_2),
		.in_wire_2_3(horizontal_tile_15_25_to_tile_15_26_3),
		.out_wire_0_0(horizontal_tile_15_26_to_tile_15_27_0),
		.out_wire_0_1(horizontal_tile_15_26_to_tile_15_27_1),
		.out_wire_0_2(horizontal_tile_15_26_to_tile_15_27_2),
		.out_wire_0_3(horizontal_tile_15_26_to_tile_15_27_3),
		.in_wire_0_0(horizontal_tile_15_27_to_tile_15_26_0),
		.in_wire_0_1(horizontal_tile_15_27_to_tile_15_26_1),
		.in_wire_0_2(horizontal_tile_15_27_to_tile_15_26_2),
		.in_wire_0_3(horizontal_tile_15_27_to_tile_15_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(507)
	);

	pe_tile pe_tile_15_27(
		.out_wire_3_0(vertical_tile_15_27_to_tile_14_27_0),
		.out_wire_3_1(vertical_tile_15_27_to_tile_14_27_1),
		.out_wire_3_2(vertical_tile_15_27_to_tile_14_27_2),
		.out_wire_3_3(vertical_tile_15_27_to_tile_14_27_3),
		.in_wire_3_0(vertical_tile_14_27_to_tile_15_27_0),
		.in_wire_3_1(vertical_tile_14_27_to_tile_15_27_1),
		.in_wire_3_2(vertical_tile_14_27_to_tile_15_27_2),
		.in_wire_3_3(vertical_tile_14_27_to_tile_15_27_3),
		.out_wire_1_0(vertical_tile_15_27_to_tile_16_27_0),
		.out_wire_1_1(vertical_tile_15_27_to_tile_16_27_1),
		.out_wire_1_2(vertical_tile_15_27_to_tile_16_27_2),
		.out_wire_1_3(vertical_tile_15_27_to_tile_16_27_3),
		.in_wire_1_0(vertical_tile_16_27_to_tile_15_27_0),
		.in_wire_1_1(vertical_tile_16_27_to_tile_15_27_1),
		.in_wire_1_2(vertical_tile_16_27_to_tile_15_27_2),
		.in_wire_1_3(vertical_tile_16_27_to_tile_15_27_3),
		.out_wire_2_0(horizontal_tile_15_27_to_tile_15_26_0),
		.out_wire_2_1(horizontal_tile_15_27_to_tile_15_26_1),
		.out_wire_2_2(horizontal_tile_15_27_to_tile_15_26_2),
		.out_wire_2_3(horizontal_tile_15_27_to_tile_15_26_3),
		.in_wire_2_0(horizontal_tile_15_26_to_tile_15_27_0),
		.in_wire_2_1(horizontal_tile_15_26_to_tile_15_27_1),
		.in_wire_2_2(horizontal_tile_15_26_to_tile_15_27_2),
		.in_wire_2_3(horizontal_tile_15_26_to_tile_15_27_3),
		.out_wire_0_0(horizontal_tile_15_27_to_tile_15_28_0),
		.out_wire_0_1(horizontal_tile_15_27_to_tile_15_28_1),
		.out_wire_0_2(horizontal_tile_15_27_to_tile_15_28_2),
		.out_wire_0_3(horizontal_tile_15_27_to_tile_15_28_3),
		.in_wire_0_0(horizontal_tile_15_28_to_tile_15_27_0),
		.in_wire_0_1(horizontal_tile_15_28_to_tile_15_27_1),
		.in_wire_0_2(horizontal_tile_15_28_to_tile_15_27_2),
		.in_wire_0_3(horizontal_tile_15_28_to_tile_15_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(508)
	);

	pe_tile pe_tile_15_28(
		.out_wire_3_0(vertical_tile_15_28_to_tile_14_28_0),
		.out_wire_3_1(vertical_tile_15_28_to_tile_14_28_1),
		.out_wire_3_2(vertical_tile_15_28_to_tile_14_28_2),
		.out_wire_3_3(vertical_tile_15_28_to_tile_14_28_3),
		.in_wire_3_0(vertical_tile_14_28_to_tile_15_28_0),
		.in_wire_3_1(vertical_tile_14_28_to_tile_15_28_1),
		.in_wire_3_2(vertical_tile_14_28_to_tile_15_28_2),
		.in_wire_3_3(vertical_tile_14_28_to_tile_15_28_3),
		.out_wire_1_0(vertical_tile_15_28_to_tile_16_28_0),
		.out_wire_1_1(vertical_tile_15_28_to_tile_16_28_1),
		.out_wire_1_2(vertical_tile_15_28_to_tile_16_28_2),
		.out_wire_1_3(vertical_tile_15_28_to_tile_16_28_3),
		.in_wire_1_0(vertical_tile_16_28_to_tile_15_28_0),
		.in_wire_1_1(vertical_tile_16_28_to_tile_15_28_1),
		.in_wire_1_2(vertical_tile_16_28_to_tile_15_28_2),
		.in_wire_1_3(vertical_tile_16_28_to_tile_15_28_3),
		.out_wire_2_0(horizontal_tile_15_28_to_tile_15_27_0),
		.out_wire_2_1(horizontal_tile_15_28_to_tile_15_27_1),
		.out_wire_2_2(horizontal_tile_15_28_to_tile_15_27_2),
		.out_wire_2_3(horizontal_tile_15_28_to_tile_15_27_3),
		.in_wire_2_0(horizontal_tile_15_27_to_tile_15_28_0),
		.in_wire_2_1(horizontal_tile_15_27_to_tile_15_28_1),
		.in_wire_2_2(horizontal_tile_15_27_to_tile_15_28_2),
		.in_wire_2_3(horizontal_tile_15_27_to_tile_15_28_3),
		.out_wire_0_0(horizontal_tile_15_28_to_tile_15_29_0),
		.out_wire_0_1(horizontal_tile_15_28_to_tile_15_29_1),
		.out_wire_0_2(horizontal_tile_15_28_to_tile_15_29_2),
		.out_wire_0_3(horizontal_tile_15_28_to_tile_15_29_3),
		.in_wire_0_0(horizontal_tile_15_29_to_tile_15_28_0),
		.in_wire_0_1(horizontal_tile_15_29_to_tile_15_28_1),
		.in_wire_0_2(horizontal_tile_15_29_to_tile_15_28_2),
		.in_wire_0_3(horizontal_tile_15_29_to_tile_15_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(509)
	);

	pe_tile pe_tile_15_29(
		.out_wire_3_0(vertical_tile_15_29_to_tile_14_29_0),
		.out_wire_3_1(vertical_tile_15_29_to_tile_14_29_1),
		.out_wire_3_2(vertical_tile_15_29_to_tile_14_29_2),
		.out_wire_3_3(vertical_tile_15_29_to_tile_14_29_3),
		.in_wire_3_0(vertical_tile_14_29_to_tile_15_29_0),
		.in_wire_3_1(vertical_tile_14_29_to_tile_15_29_1),
		.in_wire_3_2(vertical_tile_14_29_to_tile_15_29_2),
		.in_wire_3_3(vertical_tile_14_29_to_tile_15_29_3),
		.out_wire_1_0(vertical_tile_15_29_to_tile_16_29_0),
		.out_wire_1_1(vertical_tile_15_29_to_tile_16_29_1),
		.out_wire_1_2(vertical_tile_15_29_to_tile_16_29_2),
		.out_wire_1_3(vertical_tile_15_29_to_tile_16_29_3),
		.in_wire_1_0(vertical_tile_16_29_to_tile_15_29_0),
		.in_wire_1_1(vertical_tile_16_29_to_tile_15_29_1),
		.in_wire_1_2(vertical_tile_16_29_to_tile_15_29_2),
		.in_wire_1_3(vertical_tile_16_29_to_tile_15_29_3),
		.out_wire_2_0(horizontal_tile_15_29_to_tile_15_28_0),
		.out_wire_2_1(horizontal_tile_15_29_to_tile_15_28_1),
		.out_wire_2_2(horizontal_tile_15_29_to_tile_15_28_2),
		.out_wire_2_3(horizontal_tile_15_29_to_tile_15_28_3),
		.in_wire_2_0(horizontal_tile_15_28_to_tile_15_29_0),
		.in_wire_2_1(horizontal_tile_15_28_to_tile_15_29_1),
		.in_wire_2_2(horizontal_tile_15_28_to_tile_15_29_2),
		.in_wire_2_3(horizontal_tile_15_28_to_tile_15_29_3),
		.out_wire_0_0(horizontal_tile_15_29_to_tile_15_30_0),
		.out_wire_0_1(horizontal_tile_15_29_to_tile_15_30_1),
		.out_wire_0_2(horizontal_tile_15_29_to_tile_15_30_2),
		.out_wire_0_3(horizontal_tile_15_29_to_tile_15_30_3),
		.in_wire_0_0(horizontal_tile_15_30_to_tile_15_29_0),
		.in_wire_0_1(horizontal_tile_15_30_to_tile_15_29_1),
		.in_wire_0_2(horizontal_tile_15_30_to_tile_15_29_2),
		.in_wire_0_3(horizontal_tile_15_30_to_tile_15_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(510)
	);

	pe_tile pe_tile_15_30(
		.out_wire_3_0(vertical_tile_15_30_to_tile_14_30_0),
		.out_wire_3_1(vertical_tile_15_30_to_tile_14_30_1),
		.out_wire_3_2(vertical_tile_15_30_to_tile_14_30_2),
		.out_wire_3_3(vertical_tile_15_30_to_tile_14_30_3),
		.in_wire_3_0(vertical_tile_14_30_to_tile_15_30_0),
		.in_wire_3_1(vertical_tile_14_30_to_tile_15_30_1),
		.in_wire_3_2(vertical_tile_14_30_to_tile_15_30_2),
		.in_wire_3_3(vertical_tile_14_30_to_tile_15_30_3),
		.out_wire_1_0(vertical_tile_15_30_to_tile_16_30_0),
		.out_wire_1_1(vertical_tile_15_30_to_tile_16_30_1),
		.out_wire_1_2(vertical_tile_15_30_to_tile_16_30_2),
		.out_wire_1_3(vertical_tile_15_30_to_tile_16_30_3),
		.in_wire_1_0(vertical_tile_16_30_to_tile_15_30_0),
		.in_wire_1_1(vertical_tile_16_30_to_tile_15_30_1),
		.in_wire_1_2(vertical_tile_16_30_to_tile_15_30_2),
		.in_wire_1_3(vertical_tile_16_30_to_tile_15_30_3),
		.out_wire_2_0(horizontal_tile_15_30_to_tile_15_29_0),
		.out_wire_2_1(horizontal_tile_15_30_to_tile_15_29_1),
		.out_wire_2_2(horizontal_tile_15_30_to_tile_15_29_2),
		.out_wire_2_3(horizontal_tile_15_30_to_tile_15_29_3),
		.in_wire_2_0(horizontal_tile_15_29_to_tile_15_30_0),
		.in_wire_2_1(horizontal_tile_15_29_to_tile_15_30_1),
		.in_wire_2_2(horizontal_tile_15_29_to_tile_15_30_2),
		.in_wire_2_3(horizontal_tile_15_29_to_tile_15_30_3),
		.out_wire_0_0(horizontal_tile_15_30_to_tile_15_31_0),
		.out_wire_0_1(horizontal_tile_15_30_to_tile_15_31_1),
		.out_wire_0_2(horizontal_tile_15_30_to_tile_15_31_2),
		.out_wire_0_3(horizontal_tile_15_30_to_tile_15_31_3),
		.in_wire_0_0(horizontal_tile_15_31_to_tile_15_30_0),
		.in_wire_0_1(horizontal_tile_15_31_to_tile_15_30_1),
		.in_wire_0_2(horizontal_tile_15_31_to_tile_15_30_2),
		.in_wire_0_3(horizontal_tile_15_31_to_tile_15_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(511)
	);

	pe_tile_right pe_tile_15_31(
		.out_wire_3_0(vertical_tile_15_31_to_tile_14_31_0),
		.out_wire_3_1(vertical_tile_15_31_to_tile_14_31_1),
		.out_wire_3_2(vertical_tile_15_31_to_tile_14_31_2),
		.out_wire_3_3(vertical_tile_15_31_to_tile_14_31_3),
		.in_wire_3_0(vertical_tile_14_31_to_tile_15_31_0),
		.in_wire_3_1(vertical_tile_14_31_to_tile_15_31_1),
		.in_wire_3_2(vertical_tile_14_31_to_tile_15_31_2),
		.in_wire_3_3(vertical_tile_14_31_to_tile_15_31_3),
		.out_wire_1_0(vertical_tile_15_31_to_tile_16_31_0),
		.out_wire_1_1(vertical_tile_15_31_to_tile_16_31_1),
		.out_wire_1_2(vertical_tile_15_31_to_tile_16_31_2),
		.out_wire_1_3(vertical_tile_15_31_to_tile_16_31_3),
		.in_wire_1_0(vertical_tile_16_31_to_tile_15_31_0),
		.in_wire_1_1(vertical_tile_16_31_to_tile_15_31_1),
		.in_wire_1_2(vertical_tile_16_31_to_tile_15_31_2),
		.in_wire_1_3(vertical_tile_16_31_to_tile_15_31_3),
		.out_wire_2_0(horizontal_tile_15_31_to_tile_15_30_0),
		.out_wire_2_1(horizontal_tile_15_31_to_tile_15_30_1),
		.out_wire_2_2(horizontal_tile_15_31_to_tile_15_30_2),
		.out_wire_2_3(horizontal_tile_15_31_to_tile_15_30_3),
		.in_wire_2_0(horizontal_tile_15_30_to_tile_15_31_0),
		.in_wire_2_1(horizontal_tile_15_30_to_tile_15_31_1),
		.in_wire_2_2(horizontal_tile_15_30_to_tile_15_31_2),
		.in_wire_2_3(horizontal_tile_15_30_to_tile_15_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(512)
	);

	pe_tile_left pe_tile_16_0(
		.out_wire_3_0(vertical_tile_16_0_to_tile_15_0_0),
		.out_wire_3_1(vertical_tile_16_0_to_tile_15_0_1),
		.out_wire_3_2(vertical_tile_16_0_to_tile_15_0_2),
		.out_wire_3_3(vertical_tile_16_0_to_tile_15_0_3),
		.in_wire_3_0(vertical_tile_15_0_to_tile_16_0_0),
		.in_wire_3_1(vertical_tile_15_0_to_tile_16_0_1),
		.in_wire_3_2(vertical_tile_15_0_to_tile_16_0_2),
		.in_wire_3_3(vertical_tile_15_0_to_tile_16_0_3),
		.out_wire_1_0(vertical_tile_16_0_to_tile_17_0_0),
		.out_wire_1_1(vertical_tile_16_0_to_tile_17_0_1),
		.out_wire_1_2(vertical_tile_16_0_to_tile_17_0_2),
		.out_wire_1_3(vertical_tile_16_0_to_tile_17_0_3),
		.in_wire_1_0(vertical_tile_17_0_to_tile_16_0_0),
		.in_wire_1_1(vertical_tile_17_0_to_tile_16_0_1),
		.in_wire_1_2(vertical_tile_17_0_to_tile_16_0_2),
		.in_wire_1_3(vertical_tile_17_0_to_tile_16_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_16_0_to_tile_16_1_0),
		.out_wire_0_1(horizontal_tile_16_0_to_tile_16_1_1),
		.out_wire_0_2(horizontal_tile_16_0_to_tile_16_1_2),
		.out_wire_0_3(horizontal_tile_16_0_to_tile_16_1_3),
		.in_wire_0_0(horizontal_tile_16_1_to_tile_16_0_0),
		.in_wire_0_1(horizontal_tile_16_1_to_tile_16_0_1),
		.in_wire_0_2(horizontal_tile_16_1_to_tile_16_0_2),
		.in_wire_0_3(horizontal_tile_16_1_to_tile_16_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(513)
	);

	pe_tile pe_tile_16_1(
		.out_wire_3_0(vertical_tile_16_1_to_tile_15_1_0),
		.out_wire_3_1(vertical_tile_16_1_to_tile_15_1_1),
		.out_wire_3_2(vertical_tile_16_1_to_tile_15_1_2),
		.out_wire_3_3(vertical_tile_16_1_to_tile_15_1_3),
		.in_wire_3_0(vertical_tile_15_1_to_tile_16_1_0),
		.in_wire_3_1(vertical_tile_15_1_to_tile_16_1_1),
		.in_wire_3_2(vertical_tile_15_1_to_tile_16_1_2),
		.in_wire_3_3(vertical_tile_15_1_to_tile_16_1_3),
		.out_wire_1_0(vertical_tile_16_1_to_tile_17_1_0),
		.out_wire_1_1(vertical_tile_16_1_to_tile_17_1_1),
		.out_wire_1_2(vertical_tile_16_1_to_tile_17_1_2),
		.out_wire_1_3(vertical_tile_16_1_to_tile_17_1_3),
		.in_wire_1_0(vertical_tile_17_1_to_tile_16_1_0),
		.in_wire_1_1(vertical_tile_17_1_to_tile_16_1_1),
		.in_wire_1_2(vertical_tile_17_1_to_tile_16_1_2),
		.in_wire_1_3(vertical_tile_17_1_to_tile_16_1_3),
		.out_wire_2_0(horizontal_tile_16_1_to_tile_16_0_0),
		.out_wire_2_1(horizontal_tile_16_1_to_tile_16_0_1),
		.out_wire_2_2(horizontal_tile_16_1_to_tile_16_0_2),
		.out_wire_2_3(horizontal_tile_16_1_to_tile_16_0_3),
		.in_wire_2_0(horizontal_tile_16_0_to_tile_16_1_0),
		.in_wire_2_1(horizontal_tile_16_0_to_tile_16_1_1),
		.in_wire_2_2(horizontal_tile_16_0_to_tile_16_1_2),
		.in_wire_2_3(horizontal_tile_16_0_to_tile_16_1_3),
		.out_wire_0_0(horizontal_tile_16_1_to_tile_16_2_0),
		.out_wire_0_1(horizontal_tile_16_1_to_tile_16_2_1),
		.out_wire_0_2(horizontal_tile_16_1_to_tile_16_2_2),
		.out_wire_0_3(horizontal_tile_16_1_to_tile_16_2_3),
		.in_wire_0_0(horizontal_tile_16_2_to_tile_16_1_0),
		.in_wire_0_1(horizontal_tile_16_2_to_tile_16_1_1),
		.in_wire_0_2(horizontal_tile_16_2_to_tile_16_1_2),
		.in_wire_0_3(horizontal_tile_16_2_to_tile_16_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(514)
	);

	pe_tile pe_tile_16_2(
		.out_wire_3_0(vertical_tile_16_2_to_tile_15_2_0),
		.out_wire_3_1(vertical_tile_16_2_to_tile_15_2_1),
		.out_wire_3_2(vertical_tile_16_2_to_tile_15_2_2),
		.out_wire_3_3(vertical_tile_16_2_to_tile_15_2_3),
		.in_wire_3_0(vertical_tile_15_2_to_tile_16_2_0),
		.in_wire_3_1(vertical_tile_15_2_to_tile_16_2_1),
		.in_wire_3_2(vertical_tile_15_2_to_tile_16_2_2),
		.in_wire_3_3(vertical_tile_15_2_to_tile_16_2_3),
		.out_wire_1_0(vertical_tile_16_2_to_tile_17_2_0),
		.out_wire_1_1(vertical_tile_16_2_to_tile_17_2_1),
		.out_wire_1_2(vertical_tile_16_2_to_tile_17_2_2),
		.out_wire_1_3(vertical_tile_16_2_to_tile_17_2_3),
		.in_wire_1_0(vertical_tile_17_2_to_tile_16_2_0),
		.in_wire_1_1(vertical_tile_17_2_to_tile_16_2_1),
		.in_wire_1_2(vertical_tile_17_2_to_tile_16_2_2),
		.in_wire_1_3(vertical_tile_17_2_to_tile_16_2_3),
		.out_wire_2_0(horizontal_tile_16_2_to_tile_16_1_0),
		.out_wire_2_1(horizontal_tile_16_2_to_tile_16_1_1),
		.out_wire_2_2(horizontal_tile_16_2_to_tile_16_1_2),
		.out_wire_2_3(horizontal_tile_16_2_to_tile_16_1_3),
		.in_wire_2_0(horizontal_tile_16_1_to_tile_16_2_0),
		.in_wire_2_1(horizontal_tile_16_1_to_tile_16_2_1),
		.in_wire_2_2(horizontal_tile_16_1_to_tile_16_2_2),
		.in_wire_2_3(horizontal_tile_16_1_to_tile_16_2_3),
		.out_wire_0_0(horizontal_tile_16_2_to_tile_16_3_0),
		.out_wire_0_1(horizontal_tile_16_2_to_tile_16_3_1),
		.out_wire_0_2(horizontal_tile_16_2_to_tile_16_3_2),
		.out_wire_0_3(horizontal_tile_16_2_to_tile_16_3_3),
		.in_wire_0_0(horizontal_tile_16_3_to_tile_16_2_0),
		.in_wire_0_1(horizontal_tile_16_3_to_tile_16_2_1),
		.in_wire_0_2(horizontal_tile_16_3_to_tile_16_2_2),
		.in_wire_0_3(horizontal_tile_16_3_to_tile_16_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(515)
	);

	pe_tile pe_tile_16_3(
		.out_wire_3_0(vertical_tile_16_3_to_tile_15_3_0),
		.out_wire_3_1(vertical_tile_16_3_to_tile_15_3_1),
		.out_wire_3_2(vertical_tile_16_3_to_tile_15_3_2),
		.out_wire_3_3(vertical_tile_16_3_to_tile_15_3_3),
		.in_wire_3_0(vertical_tile_15_3_to_tile_16_3_0),
		.in_wire_3_1(vertical_tile_15_3_to_tile_16_3_1),
		.in_wire_3_2(vertical_tile_15_3_to_tile_16_3_2),
		.in_wire_3_3(vertical_tile_15_3_to_tile_16_3_3),
		.out_wire_1_0(vertical_tile_16_3_to_tile_17_3_0),
		.out_wire_1_1(vertical_tile_16_3_to_tile_17_3_1),
		.out_wire_1_2(vertical_tile_16_3_to_tile_17_3_2),
		.out_wire_1_3(vertical_tile_16_3_to_tile_17_3_3),
		.in_wire_1_0(vertical_tile_17_3_to_tile_16_3_0),
		.in_wire_1_1(vertical_tile_17_3_to_tile_16_3_1),
		.in_wire_1_2(vertical_tile_17_3_to_tile_16_3_2),
		.in_wire_1_3(vertical_tile_17_3_to_tile_16_3_3),
		.out_wire_2_0(horizontal_tile_16_3_to_tile_16_2_0),
		.out_wire_2_1(horizontal_tile_16_3_to_tile_16_2_1),
		.out_wire_2_2(horizontal_tile_16_3_to_tile_16_2_2),
		.out_wire_2_3(horizontal_tile_16_3_to_tile_16_2_3),
		.in_wire_2_0(horizontal_tile_16_2_to_tile_16_3_0),
		.in_wire_2_1(horizontal_tile_16_2_to_tile_16_3_1),
		.in_wire_2_2(horizontal_tile_16_2_to_tile_16_3_2),
		.in_wire_2_3(horizontal_tile_16_2_to_tile_16_3_3),
		.out_wire_0_0(horizontal_tile_16_3_to_tile_16_4_0),
		.out_wire_0_1(horizontal_tile_16_3_to_tile_16_4_1),
		.out_wire_0_2(horizontal_tile_16_3_to_tile_16_4_2),
		.out_wire_0_3(horizontal_tile_16_3_to_tile_16_4_3),
		.in_wire_0_0(horizontal_tile_16_4_to_tile_16_3_0),
		.in_wire_0_1(horizontal_tile_16_4_to_tile_16_3_1),
		.in_wire_0_2(horizontal_tile_16_4_to_tile_16_3_2),
		.in_wire_0_3(horizontal_tile_16_4_to_tile_16_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(516)
	);

	pe_tile pe_tile_16_4(
		.out_wire_3_0(vertical_tile_16_4_to_tile_15_4_0),
		.out_wire_3_1(vertical_tile_16_4_to_tile_15_4_1),
		.out_wire_3_2(vertical_tile_16_4_to_tile_15_4_2),
		.out_wire_3_3(vertical_tile_16_4_to_tile_15_4_3),
		.in_wire_3_0(vertical_tile_15_4_to_tile_16_4_0),
		.in_wire_3_1(vertical_tile_15_4_to_tile_16_4_1),
		.in_wire_3_2(vertical_tile_15_4_to_tile_16_4_2),
		.in_wire_3_3(vertical_tile_15_4_to_tile_16_4_3),
		.out_wire_1_0(vertical_tile_16_4_to_tile_17_4_0),
		.out_wire_1_1(vertical_tile_16_4_to_tile_17_4_1),
		.out_wire_1_2(vertical_tile_16_4_to_tile_17_4_2),
		.out_wire_1_3(vertical_tile_16_4_to_tile_17_4_3),
		.in_wire_1_0(vertical_tile_17_4_to_tile_16_4_0),
		.in_wire_1_1(vertical_tile_17_4_to_tile_16_4_1),
		.in_wire_1_2(vertical_tile_17_4_to_tile_16_4_2),
		.in_wire_1_3(vertical_tile_17_4_to_tile_16_4_3),
		.out_wire_2_0(horizontal_tile_16_4_to_tile_16_3_0),
		.out_wire_2_1(horizontal_tile_16_4_to_tile_16_3_1),
		.out_wire_2_2(horizontal_tile_16_4_to_tile_16_3_2),
		.out_wire_2_3(horizontal_tile_16_4_to_tile_16_3_3),
		.in_wire_2_0(horizontal_tile_16_3_to_tile_16_4_0),
		.in_wire_2_1(horizontal_tile_16_3_to_tile_16_4_1),
		.in_wire_2_2(horizontal_tile_16_3_to_tile_16_4_2),
		.in_wire_2_3(horizontal_tile_16_3_to_tile_16_4_3),
		.out_wire_0_0(horizontal_tile_16_4_to_tile_16_5_0),
		.out_wire_0_1(horizontal_tile_16_4_to_tile_16_5_1),
		.out_wire_0_2(horizontal_tile_16_4_to_tile_16_5_2),
		.out_wire_0_3(horizontal_tile_16_4_to_tile_16_5_3),
		.in_wire_0_0(horizontal_tile_16_5_to_tile_16_4_0),
		.in_wire_0_1(horizontal_tile_16_5_to_tile_16_4_1),
		.in_wire_0_2(horizontal_tile_16_5_to_tile_16_4_2),
		.in_wire_0_3(horizontal_tile_16_5_to_tile_16_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(517)
	);

	pe_tile pe_tile_16_5(
		.out_wire_3_0(vertical_tile_16_5_to_tile_15_5_0),
		.out_wire_3_1(vertical_tile_16_5_to_tile_15_5_1),
		.out_wire_3_2(vertical_tile_16_5_to_tile_15_5_2),
		.out_wire_3_3(vertical_tile_16_5_to_tile_15_5_3),
		.in_wire_3_0(vertical_tile_15_5_to_tile_16_5_0),
		.in_wire_3_1(vertical_tile_15_5_to_tile_16_5_1),
		.in_wire_3_2(vertical_tile_15_5_to_tile_16_5_2),
		.in_wire_3_3(vertical_tile_15_5_to_tile_16_5_3),
		.out_wire_1_0(vertical_tile_16_5_to_tile_17_5_0),
		.out_wire_1_1(vertical_tile_16_5_to_tile_17_5_1),
		.out_wire_1_2(vertical_tile_16_5_to_tile_17_5_2),
		.out_wire_1_3(vertical_tile_16_5_to_tile_17_5_3),
		.in_wire_1_0(vertical_tile_17_5_to_tile_16_5_0),
		.in_wire_1_1(vertical_tile_17_5_to_tile_16_5_1),
		.in_wire_1_2(vertical_tile_17_5_to_tile_16_5_2),
		.in_wire_1_3(vertical_tile_17_5_to_tile_16_5_3),
		.out_wire_2_0(horizontal_tile_16_5_to_tile_16_4_0),
		.out_wire_2_1(horizontal_tile_16_5_to_tile_16_4_1),
		.out_wire_2_2(horizontal_tile_16_5_to_tile_16_4_2),
		.out_wire_2_3(horizontal_tile_16_5_to_tile_16_4_3),
		.in_wire_2_0(horizontal_tile_16_4_to_tile_16_5_0),
		.in_wire_2_1(horizontal_tile_16_4_to_tile_16_5_1),
		.in_wire_2_2(horizontal_tile_16_4_to_tile_16_5_2),
		.in_wire_2_3(horizontal_tile_16_4_to_tile_16_5_3),
		.out_wire_0_0(horizontal_tile_16_5_to_tile_16_6_0),
		.out_wire_0_1(horizontal_tile_16_5_to_tile_16_6_1),
		.out_wire_0_2(horizontal_tile_16_5_to_tile_16_6_2),
		.out_wire_0_3(horizontal_tile_16_5_to_tile_16_6_3),
		.in_wire_0_0(horizontal_tile_16_6_to_tile_16_5_0),
		.in_wire_0_1(horizontal_tile_16_6_to_tile_16_5_1),
		.in_wire_0_2(horizontal_tile_16_6_to_tile_16_5_2),
		.in_wire_0_3(horizontal_tile_16_6_to_tile_16_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(518)
	);

	pe_tile pe_tile_16_6(
		.out_wire_3_0(vertical_tile_16_6_to_tile_15_6_0),
		.out_wire_3_1(vertical_tile_16_6_to_tile_15_6_1),
		.out_wire_3_2(vertical_tile_16_6_to_tile_15_6_2),
		.out_wire_3_3(vertical_tile_16_6_to_tile_15_6_3),
		.in_wire_3_0(vertical_tile_15_6_to_tile_16_6_0),
		.in_wire_3_1(vertical_tile_15_6_to_tile_16_6_1),
		.in_wire_3_2(vertical_tile_15_6_to_tile_16_6_2),
		.in_wire_3_3(vertical_tile_15_6_to_tile_16_6_3),
		.out_wire_1_0(vertical_tile_16_6_to_tile_17_6_0),
		.out_wire_1_1(vertical_tile_16_6_to_tile_17_6_1),
		.out_wire_1_2(vertical_tile_16_6_to_tile_17_6_2),
		.out_wire_1_3(vertical_tile_16_6_to_tile_17_6_3),
		.in_wire_1_0(vertical_tile_17_6_to_tile_16_6_0),
		.in_wire_1_1(vertical_tile_17_6_to_tile_16_6_1),
		.in_wire_1_2(vertical_tile_17_6_to_tile_16_6_2),
		.in_wire_1_3(vertical_tile_17_6_to_tile_16_6_3),
		.out_wire_2_0(horizontal_tile_16_6_to_tile_16_5_0),
		.out_wire_2_1(horizontal_tile_16_6_to_tile_16_5_1),
		.out_wire_2_2(horizontal_tile_16_6_to_tile_16_5_2),
		.out_wire_2_3(horizontal_tile_16_6_to_tile_16_5_3),
		.in_wire_2_0(horizontal_tile_16_5_to_tile_16_6_0),
		.in_wire_2_1(horizontal_tile_16_5_to_tile_16_6_1),
		.in_wire_2_2(horizontal_tile_16_5_to_tile_16_6_2),
		.in_wire_2_3(horizontal_tile_16_5_to_tile_16_6_3),
		.out_wire_0_0(horizontal_tile_16_6_to_tile_16_7_0),
		.out_wire_0_1(horizontal_tile_16_6_to_tile_16_7_1),
		.out_wire_0_2(horizontal_tile_16_6_to_tile_16_7_2),
		.out_wire_0_3(horizontal_tile_16_6_to_tile_16_7_3),
		.in_wire_0_0(horizontal_tile_16_7_to_tile_16_6_0),
		.in_wire_0_1(horizontal_tile_16_7_to_tile_16_6_1),
		.in_wire_0_2(horizontal_tile_16_7_to_tile_16_6_2),
		.in_wire_0_3(horizontal_tile_16_7_to_tile_16_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(519)
	);

	pe_tile pe_tile_16_7(
		.out_wire_3_0(vertical_tile_16_7_to_tile_15_7_0),
		.out_wire_3_1(vertical_tile_16_7_to_tile_15_7_1),
		.out_wire_3_2(vertical_tile_16_7_to_tile_15_7_2),
		.out_wire_3_3(vertical_tile_16_7_to_tile_15_7_3),
		.in_wire_3_0(vertical_tile_15_7_to_tile_16_7_0),
		.in_wire_3_1(vertical_tile_15_7_to_tile_16_7_1),
		.in_wire_3_2(vertical_tile_15_7_to_tile_16_7_2),
		.in_wire_3_3(vertical_tile_15_7_to_tile_16_7_3),
		.out_wire_1_0(vertical_tile_16_7_to_tile_17_7_0),
		.out_wire_1_1(vertical_tile_16_7_to_tile_17_7_1),
		.out_wire_1_2(vertical_tile_16_7_to_tile_17_7_2),
		.out_wire_1_3(vertical_tile_16_7_to_tile_17_7_3),
		.in_wire_1_0(vertical_tile_17_7_to_tile_16_7_0),
		.in_wire_1_1(vertical_tile_17_7_to_tile_16_7_1),
		.in_wire_1_2(vertical_tile_17_7_to_tile_16_7_2),
		.in_wire_1_3(vertical_tile_17_7_to_tile_16_7_3),
		.out_wire_2_0(horizontal_tile_16_7_to_tile_16_6_0),
		.out_wire_2_1(horizontal_tile_16_7_to_tile_16_6_1),
		.out_wire_2_2(horizontal_tile_16_7_to_tile_16_6_2),
		.out_wire_2_3(horizontal_tile_16_7_to_tile_16_6_3),
		.in_wire_2_0(horizontal_tile_16_6_to_tile_16_7_0),
		.in_wire_2_1(horizontal_tile_16_6_to_tile_16_7_1),
		.in_wire_2_2(horizontal_tile_16_6_to_tile_16_7_2),
		.in_wire_2_3(horizontal_tile_16_6_to_tile_16_7_3),
		.out_wire_0_0(horizontal_tile_16_7_to_tile_16_8_0),
		.out_wire_0_1(horizontal_tile_16_7_to_tile_16_8_1),
		.out_wire_0_2(horizontal_tile_16_7_to_tile_16_8_2),
		.out_wire_0_3(horizontal_tile_16_7_to_tile_16_8_3),
		.in_wire_0_0(horizontal_tile_16_8_to_tile_16_7_0),
		.in_wire_0_1(horizontal_tile_16_8_to_tile_16_7_1),
		.in_wire_0_2(horizontal_tile_16_8_to_tile_16_7_2),
		.in_wire_0_3(horizontal_tile_16_8_to_tile_16_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(520)
	);

	pe_tile pe_tile_16_8(
		.out_wire_3_0(vertical_tile_16_8_to_tile_15_8_0),
		.out_wire_3_1(vertical_tile_16_8_to_tile_15_8_1),
		.out_wire_3_2(vertical_tile_16_8_to_tile_15_8_2),
		.out_wire_3_3(vertical_tile_16_8_to_tile_15_8_3),
		.in_wire_3_0(vertical_tile_15_8_to_tile_16_8_0),
		.in_wire_3_1(vertical_tile_15_8_to_tile_16_8_1),
		.in_wire_3_2(vertical_tile_15_8_to_tile_16_8_2),
		.in_wire_3_3(vertical_tile_15_8_to_tile_16_8_3),
		.out_wire_1_0(vertical_tile_16_8_to_tile_17_8_0),
		.out_wire_1_1(vertical_tile_16_8_to_tile_17_8_1),
		.out_wire_1_2(vertical_tile_16_8_to_tile_17_8_2),
		.out_wire_1_3(vertical_tile_16_8_to_tile_17_8_3),
		.in_wire_1_0(vertical_tile_17_8_to_tile_16_8_0),
		.in_wire_1_1(vertical_tile_17_8_to_tile_16_8_1),
		.in_wire_1_2(vertical_tile_17_8_to_tile_16_8_2),
		.in_wire_1_3(vertical_tile_17_8_to_tile_16_8_3),
		.out_wire_2_0(horizontal_tile_16_8_to_tile_16_7_0),
		.out_wire_2_1(horizontal_tile_16_8_to_tile_16_7_1),
		.out_wire_2_2(horizontal_tile_16_8_to_tile_16_7_2),
		.out_wire_2_3(horizontal_tile_16_8_to_tile_16_7_3),
		.in_wire_2_0(horizontal_tile_16_7_to_tile_16_8_0),
		.in_wire_2_1(horizontal_tile_16_7_to_tile_16_8_1),
		.in_wire_2_2(horizontal_tile_16_7_to_tile_16_8_2),
		.in_wire_2_3(horizontal_tile_16_7_to_tile_16_8_3),
		.out_wire_0_0(horizontal_tile_16_8_to_tile_16_9_0),
		.out_wire_0_1(horizontal_tile_16_8_to_tile_16_9_1),
		.out_wire_0_2(horizontal_tile_16_8_to_tile_16_9_2),
		.out_wire_0_3(horizontal_tile_16_8_to_tile_16_9_3),
		.in_wire_0_0(horizontal_tile_16_9_to_tile_16_8_0),
		.in_wire_0_1(horizontal_tile_16_9_to_tile_16_8_1),
		.in_wire_0_2(horizontal_tile_16_9_to_tile_16_8_2),
		.in_wire_0_3(horizontal_tile_16_9_to_tile_16_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(521)
	);

	pe_tile pe_tile_16_9(
		.out_wire_3_0(vertical_tile_16_9_to_tile_15_9_0),
		.out_wire_3_1(vertical_tile_16_9_to_tile_15_9_1),
		.out_wire_3_2(vertical_tile_16_9_to_tile_15_9_2),
		.out_wire_3_3(vertical_tile_16_9_to_tile_15_9_3),
		.in_wire_3_0(vertical_tile_15_9_to_tile_16_9_0),
		.in_wire_3_1(vertical_tile_15_9_to_tile_16_9_1),
		.in_wire_3_2(vertical_tile_15_9_to_tile_16_9_2),
		.in_wire_3_3(vertical_tile_15_9_to_tile_16_9_3),
		.out_wire_1_0(vertical_tile_16_9_to_tile_17_9_0),
		.out_wire_1_1(vertical_tile_16_9_to_tile_17_9_1),
		.out_wire_1_2(vertical_tile_16_9_to_tile_17_9_2),
		.out_wire_1_3(vertical_tile_16_9_to_tile_17_9_3),
		.in_wire_1_0(vertical_tile_17_9_to_tile_16_9_0),
		.in_wire_1_1(vertical_tile_17_9_to_tile_16_9_1),
		.in_wire_1_2(vertical_tile_17_9_to_tile_16_9_2),
		.in_wire_1_3(vertical_tile_17_9_to_tile_16_9_3),
		.out_wire_2_0(horizontal_tile_16_9_to_tile_16_8_0),
		.out_wire_2_1(horizontal_tile_16_9_to_tile_16_8_1),
		.out_wire_2_2(horizontal_tile_16_9_to_tile_16_8_2),
		.out_wire_2_3(horizontal_tile_16_9_to_tile_16_8_3),
		.in_wire_2_0(horizontal_tile_16_8_to_tile_16_9_0),
		.in_wire_2_1(horizontal_tile_16_8_to_tile_16_9_1),
		.in_wire_2_2(horizontal_tile_16_8_to_tile_16_9_2),
		.in_wire_2_3(horizontal_tile_16_8_to_tile_16_9_3),
		.out_wire_0_0(horizontal_tile_16_9_to_tile_16_10_0),
		.out_wire_0_1(horizontal_tile_16_9_to_tile_16_10_1),
		.out_wire_0_2(horizontal_tile_16_9_to_tile_16_10_2),
		.out_wire_0_3(horizontal_tile_16_9_to_tile_16_10_3),
		.in_wire_0_0(horizontal_tile_16_10_to_tile_16_9_0),
		.in_wire_0_1(horizontal_tile_16_10_to_tile_16_9_1),
		.in_wire_0_2(horizontal_tile_16_10_to_tile_16_9_2),
		.in_wire_0_3(horizontal_tile_16_10_to_tile_16_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(522)
	);

	pe_tile pe_tile_16_10(
		.out_wire_3_0(vertical_tile_16_10_to_tile_15_10_0),
		.out_wire_3_1(vertical_tile_16_10_to_tile_15_10_1),
		.out_wire_3_2(vertical_tile_16_10_to_tile_15_10_2),
		.out_wire_3_3(vertical_tile_16_10_to_tile_15_10_3),
		.in_wire_3_0(vertical_tile_15_10_to_tile_16_10_0),
		.in_wire_3_1(vertical_tile_15_10_to_tile_16_10_1),
		.in_wire_3_2(vertical_tile_15_10_to_tile_16_10_2),
		.in_wire_3_3(vertical_tile_15_10_to_tile_16_10_3),
		.out_wire_1_0(vertical_tile_16_10_to_tile_17_10_0),
		.out_wire_1_1(vertical_tile_16_10_to_tile_17_10_1),
		.out_wire_1_2(vertical_tile_16_10_to_tile_17_10_2),
		.out_wire_1_3(vertical_tile_16_10_to_tile_17_10_3),
		.in_wire_1_0(vertical_tile_17_10_to_tile_16_10_0),
		.in_wire_1_1(vertical_tile_17_10_to_tile_16_10_1),
		.in_wire_1_2(vertical_tile_17_10_to_tile_16_10_2),
		.in_wire_1_3(vertical_tile_17_10_to_tile_16_10_3),
		.out_wire_2_0(horizontal_tile_16_10_to_tile_16_9_0),
		.out_wire_2_1(horizontal_tile_16_10_to_tile_16_9_1),
		.out_wire_2_2(horizontal_tile_16_10_to_tile_16_9_2),
		.out_wire_2_3(horizontal_tile_16_10_to_tile_16_9_3),
		.in_wire_2_0(horizontal_tile_16_9_to_tile_16_10_0),
		.in_wire_2_1(horizontal_tile_16_9_to_tile_16_10_1),
		.in_wire_2_2(horizontal_tile_16_9_to_tile_16_10_2),
		.in_wire_2_3(horizontal_tile_16_9_to_tile_16_10_3),
		.out_wire_0_0(horizontal_tile_16_10_to_tile_16_11_0),
		.out_wire_0_1(horizontal_tile_16_10_to_tile_16_11_1),
		.out_wire_0_2(horizontal_tile_16_10_to_tile_16_11_2),
		.out_wire_0_3(horizontal_tile_16_10_to_tile_16_11_3),
		.in_wire_0_0(horizontal_tile_16_11_to_tile_16_10_0),
		.in_wire_0_1(horizontal_tile_16_11_to_tile_16_10_1),
		.in_wire_0_2(horizontal_tile_16_11_to_tile_16_10_2),
		.in_wire_0_3(horizontal_tile_16_11_to_tile_16_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(523)
	);

	pe_tile pe_tile_16_11(
		.out_wire_3_0(vertical_tile_16_11_to_tile_15_11_0),
		.out_wire_3_1(vertical_tile_16_11_to_tile_15_11_1),
		.out_wire_3_2(vertical_tile_16_11_to_tile_15_11_2),
		.out_wire_3_3(vertical_tile_16_11_to_tile_15_11_3),
		.in_wire_3_0(vertical_tile_15_11_to_tile_16_11_0),
		.in_wire_3_1(vertical_tile_15_11_to_tile_16_11_1),
		.in_wire_3_2(vertical_tile_15_11_to_tile_16_11_2),
		.in_wire_3_3(vertical_tile_15_11_to_tile_16_11_3),
		.out_wire_1_0(vertical_tile_16_11_to_tile_17_11_0),
		.out_wire_1_1(vertical_tile_16_11_to_tile_17_11_1),
		.out_wire_1_2(vertical_tile_16_11_to_tile_17_11_2),
		.out_wire_1_3(vertical_tile_16_11_to_tile_17_11_3),
		.in_wire_1_0(vertical_tile_17_11_to_tile_16_11_0),
		.in_wire_1_1(vertical_tile_17_11_to_tile_16_11_1),
		.in_wire_1_2(vertical_tile_17_11_to_tile_16_11_2),
		.in_wire_1_3(vertical_tile_17_11_to_tile_16_11_3),
		.out_wire_2_0(horizontal_tile_16_11_to_tile_16_10_0),
		.out_wire_2_1(horizontal_tile_16_11_to_tile_16_10_1),
		.out_wire_2_2(horizontal_tile_16_11_to_tile_16_10_2),
		.out_wire_2_3(horizontal_tile_16_11_to_tile_16_10_3),
		.in_wire_2_0(horizontal_tile_16_10_to_tile_16_11_0),
		.in_wire_2_1(horizontal_tile_16_10_to_tile_16_11_1),
		.in_wire_2_2(horizontal_tile_16_10_to_tile_16_11_2),
		.in_wire_2_3(horizontal_tile_16_10_to_tile_16_11_3),
		.out_wire_0_0(horizontal_tile_16_11_to_tile_16_12_0),
		.out_wire_0_1(horizontal_tile_16_11_to_tile_16_12_1),
		.out_wire_0_2(horizontal_tile_16_11_to_tile_16_12_2),
		.out_wire_0_3(horizontal_tile_16_11_to_tile_16_12_3),
		.in_wire_0_0(horizontal_tile_16_12_to_tile_16_11_0),
		.in_wire_0_1(horizontal_tile_16_12_to_tile_16_11_1),
		.in_wire_0_2(horizontal_tile_16_12_to_tile_16_11_2),
		.in_wire_0_3(horizontal_tile_16_12_to_tile_16_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(524)
	);

	pe_tile pe_tile_16_12(
		.out_wire_3_0(vertical_tile_16_12_to_tile_15_12_0),
		.out_wire_3_1(vertical_tile_16_12_to_tile_15_12_1),
		.out_wire_3_2(vertical_tile_16_12_to_tile_15_12_2),
		.out_wire_3_3(vertical_tile_16_12_to_tile_15_12_3),
		.in_wire_3_0(vertical_tile_15_12_to_tile_16_12_0),
		.in_wire_3_1(vertical_tile_15_12_to_tile_16_12_1),
		.in_wire_3_2(vertical_tile_15_12_to_tile_16_12_2),
		.in_wire_3_3(vertical_tile_15_12_to_tile_16_12_3),
		.out_wire_1_0(vertical_tile_16_12_to_tile_17_12_0),
		.out_wire_1_1(vertical_tile_16_12_to_tile_17_12_1),
		.out_wire_1_2(vertical_tile_16_12_to_tile_17_12_2),
		.out_wire_1_3(vertical_tile_16_12_to_tile_17_12_3),
		.in_wire_1_0(vertical_tile_17_12_to_tile_16_12_0),
		.in_wire_1_1(vertical_tile_17_12_to_tile_16_12_1),
		.in_wire_1_2(vertical_tile_17_12_to_tile_16_12_2),
		.in_wire_1_3(vertical_tile_17_12_to_tile_16_12_3),
		.out_wire_2_0(horizontal_tile_16_12_to_tile_16_11_0),
		.out_wire_2_1(horizontal_tile_16_12_to_tile_16_11_1),
		.out_wire_2_2(horizontal_tile_16_12_to_tile_16_11_2),
		.out_wire_2_3(horizontal_tile_16_12_to_tile_16_11_3),
		.in_wire_2_0(horizontal_tile_16_11_to_tile_16_12_0),
		.in_wire_2_1(horizontal_tile_16_11_to_tile_16_12_1),
		.in_wire_2_2(horizontal_tile_16_11_to_tile_16_12_2),
		.in_wire_2_3(horizontal_tile_16_11_to_tile_16_12_3),
		.out_wire_0_0(horizontal_tile_16_12_to_tile_16_13_0),
		.out_wire_0_1(horizontal_tile_16_12_to_tile_16_13_1),
		.out_wire_0_2(horizontal_tile_16_12_to_tile_16_13_2),
		.out_wire_0_3(horizontal_tile_16_12_to_tile_16_13_3),
		.in_wire_0_0(horizontal_tile_16_13_to_tile_16_12_0),
		.in_wire_0_1(horizontal_tile_16_13_to_tile_16_12_1),
		.in_wire_0_2(horizontal_tile_16_13_to_tile_16_12_2),
		.in_wire_0_3(horizontal_tile_16_13_to_tile_16_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(525)
	);

	pe_tile pe_tile_16_13(
		.out_wire_3_0(vertical_tile_16_13_to_tile_15_13_0),
		.out_wire_3_1(vertical_tile_16_13_to_tile_15_13_1),
		.out_wire_3_2(vertical_tile_16_13_to_tile_15_13_2),
		.out_wire_3_3(vertical_tile_16_13_to_tile_15_13_3),
		.in_wire_3_0(vertical_tile_15_13_to_tile_16_13_0),
		.in_wire_3_1(vertical_tile_15_13_to_tile_16_13_1),
		.in_wire_3_2(vertical_tile_15_13_to_tile_16_13_2),
		.in_wire_3_3(vertical_tile_15_13_to_tile_16_13_3),
		.out_wire_1_0(vertical_tile_16_13_to_tile_17_13_0),
		.out_wire_1_1(vertical_tile_16_13_to_tile_17_13_1),
		.out_wire_1_2(vertical_tile_16_13_to_tile_17_13_2),
		.out_wire_1_3(vertical_tile_16_13_to_tile_17_13_3),
		.in_wire_1_0(vertical_tile_17_13_to_tile_16_13_0),
		.in_wire_1_1(vertical_tile_17_13_to_tile_16_13_1),
		.in_wire_1_2(vertical_tile_17_13_to_tile_16_13_2),
		.in_wire_1_3(vertical_tile_17_13_to_tile_16_13_3),
		.out_wire_2_0(horizontal_tile_16_13_to_tile_16_12_0),
		.out_wire_2_1(horizontal_tile_16_13_to_tile_16_12_1),
		.out_wire_2_2(horizontal_tile_16_13_to_tile_16_12_2),
		.out_wire_2_3(horizontal_tile_16_13_to_tile_16_12_3),
		.in_wire_2_0(horizontal_tile_16_12_to_tile_16_13_0),
		.in_wire_2_1(horizontal_tile_16_12_to_tile_16_13_1),
		.in_wire_2_2(horizontal_tile_16_12_to_tile_16_13_2),
		.in_wire_2_3(horizontal_tile_16_12_to_tile_16_13_3),
		.out_wire_0_0(horizontal_tile_16_13_to_tile_16_14_0),
		.out_wire_0_1(horizontal_tile_16_13_to_tile_16_14_1),
		.out_wire_0_2(horizontal_tile_16_13_to_tile_16_14_2),
		.out_wire_0_3(horizontal_tile_16_13_to_tile_16_14_3),
		.in_wire_0_0(horizontal_tile_16_14_to_tile_16_13_0),
		.in_wire_0_1(horizontal_tile_16_14_to_tile_16_13_1),
		.in_wire_0_2(horizontal_tile_16_14_to_tile_16_13_2),
		.in_wire_0_3(horizontal_tile_16_14_to_tile_16_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(526)
	);

	pe_tile pe_tile_16_14(
		.out_wire_3_0(vertical_tile_16_14_to_tile_15_14_0),
		.out_wire_3_1(vertical_tile_16_14_to_tile_15_14_1),
		.out_wire_3_2(vertical_tile_16_14_to_tile_15_14_2),
		.out_wire_3_3(vertical_tile_16_14_to_tile_15_14_3),
		.in_wire_3_0(vertical_tile_15_14_to_tile_16_14_0),
		.in_wire_3_1(vertical_tile_15_14_to_tile_16_14_1),
		.in_wire_3_2(vertical_tile_15_14_to_tile_16_14_2),
		.in_wire_3_3(vertical_tile_15_14_to_tile_16_14_3),
		.out_wire_1_0(vertical_tile_16_14_to_tile_17_14_0),
		.out_wire_1_1(vertical_tile_16_14_to_tile_17_14_1),
		.out_wire_1_2(vertical_tile_16_14_to_tile_17_14_2),
		.out_wire_1_3(vertical_tile_16_14_to_tile_17_14_3),
		.in_wire_1_0(vertical_tile_17_14_to_tile_16_14_0),
		.in_wire_1_1(vertical_tile_17_14_to_tile_16_14_1),
		.in_wire_1_2(vertical_tile_17_14_to_tile_16_14_2),
		.in_wire_1_3(vertical_tile_17_14_to_tile_16_14_3),
		.out_wire_2_0(horizontal_tile_16_14_to_tile_16_13_0),
		.out_wire_2_1(horizontal_tile_16_14_to_tile_16_13_1),
		.out_wire_2_2(horizontal_tile_16_14_to_tile_16_13_2),
		.out_wire_2_3(horizontal_tile_16_14_to_tile_16_13_3),
		.in_wire_2_0(horizontal_tile_16_13_to_tile_16_14_0),
		.in_wire_2_1(horizontal_tile_16_13_to_tile_16_14_1),
		.in_wire_2_2(horizontal_tile_16_13_to_tile_16_14_2),
		.in_wire_2_3(horizontal_tile_16_13_to_tile_16_14_3),
		.out_wire_0_0(horizontal_tile_16_14_to_tile_16_15_0),
		.out_wire_0_1(horizontal_tile_16_14_to_tile_16_15_1),
		.out_wire_0_2(horizontal_tile_16_14_to_tile_16_15_2),
		.out_wire_0_3(horizontal_tile_16_14_to_tile_16_15_3),
		.in_wire_0_0(horizontal_tile_16_15_to_tile_16_14_0),
		.in_wire_0_1(horizontal_tile_16_15_to_tile_16_14_1),
		.in_wire_0_2(horizontal_tile_16_15_to_tile_16_14_2),
		.in_wire_0_3(horizontal_tile_16_15_to_tile_16_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(527)
	);

	pe_tile pe_tile_16_15(
		.out_wire_3_0(vertical_tile_16_15_to_tile_15_15_0),
		.out_wire_3_1(vertical_tile_16_15_to_tile_15_15_1),
		.out_wire_3_2(vertical_tile_16_15_to_tile_15_15_2),
		.out_wire_3_3(vertical_tile_16_15_to_tile_15_15_3),
		.in_wire_3_0(vertical_tile_15_15_to_tile_16_15_0),
		.in_wire_3_1(vertical_tile_15_15_to_tile_16_15_1),
		.in_wire_3_2(vertical_tile_15_15_to_tile_16_15_2),
		.in_wire_3_3(vertical_tile_15_15_to_tile_16_15_3),
		.out_wire_1_0(vertical_tile_16_15_to_tile_17_15_0),
		.out_wire_1_1(vertical_tile_16_15_to_tile_17_15_1),
		.out_wire_1_2(vertical_tile_16_15_to_tile_17_15_2),
		.out_wire_1_3(vertical_tile_16_15_to_tile_17_15_3),
		.in_wire_1_0(vertical_tile_17_15_to_tile_16_15_0),
		.in_wire_1_1(vertical_tile_17_15_to_tile_16_15_1),
		.in_wire_1_2(vertical_tile_17_15_to_tile_16_15_2),
		.in_wire_1_3(vertical_tile_17_15_to_tile_16_15_3),
		.out_wire_2_0(horizontal_tile_16_15_to_tile_16_14_0),
		.out_wire_2_1(horizontal_tile_16_15_to_tile_16_14_1),
		.out_wire_2_2(horizontal_tile_16_15_to_tile_16_14_2),
		.out_wire_2_3(horizontal_tile_16_15_to_tile_16_14_3),
		.in_wire_2_0(horizontal_tile_16_14_to_tile_16_15_0),
		.in_wire_2_1(horizontal_tile_16_14_to_tile_16_15_1),
		.in_wire_2_2(horizontal_tile_16_14_to_tile_16_15_2),
		.in_wire_2_3(horizontal_tile_16_14_to_tile_16_15_3),
		.out_wire_0_0(horizontal_tile_16_15_to_tile_16_16_0),
		.out_wire_0_1(horizontal_tile_16_15_to_tile_16_16_1),
		.out_wire_0_2(horizontal_tile_16_15_to_tile_16_16_2),
		.out_wire_0_3(horizontal_tile_16_15_to_tile_16_16_3),
		.in_wire_0_0(horizontal_tile_16_16_to_tile_16_15_0),
		.in_wire_0_1(horizontal_tile_16_16_to_tile_16_15_1),
		.in_wire_0_2(horizontal_tile_16_16_to_tile_16_15_2),
		.in_wire_0_3(horizontal_tile_16_16_to_tile_16_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(528)
	);

	pe_tile pe_tile_16_16(
		.out_wire_3_0(vertical_tile_16_16_to_tile_15_16_0),
		.out_wire_3_1(vertical_tile_16_16_to_tile_15_16_1),
		.out_wire_3_2(vertical_tile_16_16_to_tile_15_16_2),
		.out_wire_3_3(vertical_tile_16_16_to_tile_15_16_3),
		.in_wire_3_0(vertical_tile_15_16_to_tile_16_16_0),
		.in_wire_3_1(vertical_tile_15_16_to_tile_16_16_1),
		.in_wire_3_2(vertical_tile_15_16_to_tile_16_16_2),
		.in_wire_3_3(vertical_tile_15_16_to_tile_16_16_3),
		.out_wire_1_0(vertical_tile_16_16_to_tile_17_16_0),
		.out_wire_1_1(vertical_tile_16_16_to_tile_17_16_1),
		.out_wire_1_2(vertical_tile_16_16_to_tile_17_16_2),
		.out_wire_1_3(vertical_tile_16_16_to_tile_17_16_3),
		.in_wire_1_0(vertical_tile_17_16_to_tile_16_16_0),
		.in_wire_1_1(vertical_tile_17_16_to_tile_16_16_1),
		.in_wire_1_2(vertical_tile_17_16_to_tile_16_16_2),
		.in_wire_1_3(vertical_tile_17_16_to_tile_16_16_3),
		.out_wire_2_0(horizontal_tile_16_16_to_tile_16_15_0),
		.out_wire_2_1(horizontal_tile_16_16_to_tile_16_15_1),
		.out_wire_2_2(horizontal_tile_16_16_to_tile_16_15_2),
		.out_wire_2_3(horizontal_tile_16_16_to_tile_16_15_3),
		.in_wire_2_0(horizontal_tile_16_15_to_tile_16_16_0),
		.in_wire_2_1(horizontal_tile_16_15_to_tile_16_16_1),
		.in_wire_2_2(horizontal_tile_16_15_to_tile_16_16_2),
		.in_wire_2_3(horizontal_tile_16_15_to_tile_16_16_3),
		.out_wire_0_0(horizontal_tile_16_16_to_tile_16_17_0),
		.out_wire_0_1(horizontal_tile_16_16_to_tile_16_17_1),
		.out_wire_0_2(horizontal_tile_16_16_to_tile_16_17_2),
		.out_wire_0_3(horizontal_tile_16_16_to_tile_16_17_3),
		.in_wire_0_0(horizontal_tile_16_17_to_tile_16_16_0),
		.in_wire_0_1(horizontal_tile_16_17_to_tile_16_16_1),
		.in_wire_0_2(horizontal_tile_16_17_to_tile_16_16_2),
		.in_wire_0_3(horizontal_tile_16_17_to_tile_16_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(529)
	);

	pe_tile pe_tile_16_17(
		.out_wire_3_0(vertical_tile_16_17_to_tile_15_17_0),
		.out_wire_3_1(vertical_tile_16_17_to_tile_15_17_1),
		.out_wire_3_2(vertical_tile_16_17_to_tile_15_17_2),
		.out_wire_3_3(vertical_tile_16_17_to_tile_15_17_3),
		.in_wire_3_0(vertical_tile_15_17_to_tile_16_17_0),
		.in_wire_3_1(vertical_tile_15_17_to_tile_16_17_1),
		.in_wire_3_2(vertical_tile_15_17_to_tile_16_17_2),
		.in_wire_3_3(vertical_tile_15_17_to_tile_16_17_3),
		.out_wire_1_0(vertical_tile_16_17_to_tile_17_17_0),
		.out_wire_1_1(vertical_tile_16_17_to_tile_17_17_1),
		.out_wire_1_2(vertical_tile_16_17_to_tile_17_17_2),
		.out_wire_1_3(vertical_tile_16_17_to_tile_17_17_3),
		.in_wire_1_0(vertical_tile_17_17_to_tile_16_17_0),
		.in_wire_1_1(vertical_tile_17_17_to_tile_16_17_1),
		.in_wire_1_2(vertical_tile_17_17_to_tile_16_17_2),
		.in_wire_1_3(vertical_tile_17_17_to_tile_16_17_3),
		.out_wire_2_0(horizontal_tile_16_17_to_tile_16_16_0),
		.out_wire_2_1(horizontal_tile_16_17_to_tile_16_16_1),
		.out_wire_2_2(horizontal_tile_16_17_to_tile_16_16_2),
		.out_wire_2_3(horizontal_tile_16_17_to_tile_16_16_3),
		.in_wire_2_0(horizontal_tile_16_16_to_tile_16_17_0),
		.in_wire_2_1(horizontal_tile_16_16_to_tile_16_17_1),
		.in_wire_2_2(horizontal_tile_16_16_to_tile_16_17_2),
		.in_wire_2_3(horizontal_tile_16_16_to_tile_16_17_3),
		.out_wire_0_0(horizontal_tile_16_17_to_tile_16_18_0),
		.out_wire_0_1(horizontal_tile_16_17_to_tile_16_18_1),
		.out_wire_0_2(horizontal_tile_16_17_to_tile_16_18_2),
		.out_wire_0_3(horizontal_tile_16_17_to_tile_16_18_3),
		.in_wire_0_0(horizontal_tile_16_18_to_tile_16_17_0),
		.in_wire_0_1(horizontal_tile_16_18_to_tile_16_17_1),
		.in_wire_0_2(horizontal_tile_16_18_to_tile_16_17_2),
		.in_wire_0_3(horizontal_tile_16_18_to_tile_16_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(530)
	);

	pe_tile pe_tile_16_18(
		.out_wire_3_0(vertical_tile_16_18_to_tile_15_18_0),
		.out_wire_3_1(vertical_tile_16_18_to_tile_15_18_1),
		.out_wire_3_2(vertical_tile_16_18_to_tile_15_18_2),
		.out_wire_3_3(vertical_tile_16_18_to_tile_15_18_3),
		.in_wire_3_0(vertical_tile_15_18_to_tile_16_18_0),
		.in_wire_3_1(vertical_tile_15_18_to_tile_16_18_1),
		.in_wire_3_2(vertical_tile_15_18_to_tile_16_18_2),
		.in_wire_3_3(vertical_tile_15_18_to_tile_16_18_3),
		.out_wire_1_0(vertical_tile_16_18_to_tile_17_18_0),
		.out_wire_1_1(vertical_tile_16_18_to_tile_17_18_1),
		.out_wire_1_2(vertical_tile_16_18_to_tile_17_18_2),
		.out_wire_1_3(vertical_tile_16_18_to_tile_17_18_3),
		.in_wire_1_0(vertical_tile_17_18_to_tile_16_18_0),
		.in_wire_1_1(vertical_tile_17_18_to_tile_16_18_1),
		.in_wire_1_2(vertical_tile_17_18_to_tile_16_18_2),
		.in_wire_1_3(vertical_tile_17_18_to_tile_16_18_3),
		.out_wire_2_0(horizontal_tile_16_18_to_tile_16_17_0),
		.out_wire_2_1(horizontal_tile_16_18_to_tile_16_17_1),
		.out_wire_2_2(horizontal_tile_16_18_to_tile_16_17_2),
		.out_wire_2_3(horizontal_tile_16_18_to_tile_16_17_3),
		.in_wire_2_0(horizontal_tile_16_17_to_tile_16_18_0),
		.in_wire_2_1(horizontal_tile_16_17_to_tile_16_18_1),
		.in_wire_2_2(horizontal_tile_16_17_to_tile_16_18_2),
		.in_wire_2_3(horizontal_tile_16_17_to_tile_16_18_3),
		.out_wire_0_0(horizontal_tile_16_18_to_tile_16_19_0),
		.out_wire_0_1(horizontal_tile_16_18_to_tile_16_19_1),
		.out_wire_0_2(horizontal_tile_16_18_to_tile_16_19_2),
		.out_wire_0_3(horizontal_tile_16_18_to_tile_16_19_3),
		.in_wire_0_0(horizontal_tile_16_19_to_tile_16_18_0),
		.in_wire_0_1(horizontal_tile_16_19_to_tile_16_18_1),
		.in_wire_0_2(horizontal_tile_16_19_to_tile_16_18_2),
		.in_wire_0_3(horizontal_tile_16_19_to_tile_16_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(531)
	);

	pe_tile pe_tile_16_19(
		.out_wire_3_0(vertical_tile_16_19_to_tile_15_19_0),
		.out_wire_3_1(vertical_tile_16_19_to_tile_15_19_1),
		.out_wire_3_2(vertical_tile_16_19_to_tile_15_19_2),
		.out_wire_3_3(vertical_tile_16_19_to_tile_15_19_3),
		.in_wire_3_0(vertical_tile_15_19_to_tile_16_19_0),
		.in_wire_3_1(vertical_tile_15_19_to_tile_16_19_1),
		.in_wire_3_2(vertical_tile_15_19_to_tile_16_19_2),
		.in_wire_3_3(vertical_tile_15_19_to_tile_16_19_3),
		.out_wire_1_0(vertical_tile_16_19_to_tile_17_19_0),
		.out_wire_1_1(vertical_tile_16_19_to_tile_17_19_1),
		.out_wire_1_2(vertical_tile_16_19_to_tile_17_19_2),
		.out_wire_1_3(vertical_tile_16_19_to_tile_17_19_3),
		.in_wire_1_0(vertical_tile_17_19_to_tile_16_19_0),
		.in_wire_1_1(vertical_tile_17_19_to_tile_16_19_1),
		.in_wire_1_2(vertical_tile_17_19_to_tile_16_19_2),
		.in_wire_1_3(vertical_tile_17_19_to_tile_16_19_3),
		.out_wire_2_0(horizontal_tile_16_19_to_tile_16_18_0),
		.out_wire_2_1(horizontal_tile_16_19_to_tile_16_18_1),
		.out_wire_2_2(horizontal_tile_16_19_to_tile_16_18_2),
		.out_wire_2_3(horizontal_tile_16_19_to_tile_16_18_3),
		.in_wire_2_0(horizontal_tile_16_18_to_tile_16_19_0),
		.in_wire_2_1(horizontal_tile_16_18_to_tile_16_19_1),
		.in_wire_2_2(horizontal_tile_16_18_to_tile_16_19_2),
		.in_wire_2_3(horizontal_tile_16_18_to_tile_16_19_3),
		.out_wire_0_0(horizontal_tile_16_19_to_tile_16_20_0),
		.out_wire_0_1(horizontal_tile_16_19_to_tile_16_20_1),
		.out_wire_0_2(horizontal_tile_16_19_to_tile_16_20_2),
		.out_wire_0_3(horizontal_tile_16_19_to_tile_16_20_3),
		.in_wire_0_0(horizontal_tile_16_20_to_tile_16_19_0),
		.in_wire_0_1(horizontal_tile_16_20_to_tile_16_19_1),
		.in_wire_0_2(horizontal_tile_16_20_to_tile_16_19_2),
		.in_wire_0_3(horizontal_tile_16_20_to_tile_16_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(532)
	);

	pe_tile pe_tile_16_20(
		.out_wire_3_0(vertical_tile_16_20_to_tile_15_20_0),
		.out_wire_3_1(vertical_tile_16_20_to_tile_15_20_1),
		.out_wire_3_2(vertical_tile_16_20_to_tile_15_20_2),
		.out_wire_3_3(vertical_tile_16_20_to_tile_15_20_3),
		.in_wire_3_0(vertical_tile_15_20_to_tile_16_20_0),
		.in_wire_3_1(vertical_tile_15_20_to_tile_16_20_1),
		.in_wire_3_2(vertical_tile_15_20_to_tile_16_20_2),
		.in_wire_3_3(vertical_tile_15_20_to_tile_16_20_3),
		.out_wire_1_0(vertical_tile_16_20_to_tile_17_20_0),
		.out_wire_1_1(vertical_tile_16_20_to_tile_17_20_1),
		.out_wire_1_2(vertical_tile_16_20_to_tile_17_20_2),
		.out_wire_1_3(vertical_tile_16_20_to_tile_17_20_3),
		.in_wire_1_0(vertical_tile_17_20_to_tile_16_20_0),
		.in_wire_1_1(vertical_tile_17_20_to_tile_16_20_1),
		.in_wire_1_2(vertical_tile_17_20_to_tile_16_20_2),
		.in_wire_1_3(vertical_tile_17_20_to_tile_16_20_3),
		.out_wire_2_0(horizontal_tile_16_20_to_tile_16_19_0),
		.out_wire_2_1(horizontal_tile_16_20_to_tile_16_19_1),
		.out_wire_2_2(horizontal_tile_16_20_to_tile_16_19_2),
		.out_wire_2_3(horizontal_tile_16_20_to_tile_16_19_3),
		.in_wire_2_0(horizontal_tile_16_19_to_tile_16_20_0),
		.in_wire_2_1(horizontal_tile_16_19_to_tile_16_20_1),
		.in_wire_2_2(horizontal_tile_16_19_to_tile_16_20_2),
		.in_wire_2_3(horizontal_tile_16_19_to_tile_16_20_3),
		.out_wire_0_0(horizontal_tile_16_20_to_tile_16_21_0),
		.out_wire_0_1(horizontal_tile_16_20_to_tile_16_21_1),
		.out_wire_0_2(horizontal_tile_16_20_to_tile_16_21_2),
		.out_wire_0_3(horizontal_tile_16_20_to_tile_16_21_3),
		.in_wire_0_0(horizontal_tile_16_21_to_tile_16_20_0),
		.in_wire_0_1(horizontal_tile_16_21_to_tile_16_20_1),
		.in_wire_0_2(horizontal_tile_16_21_to_tile_16_20_2),
		.in_wire_0_3(horizontal_tile_16_21_to_tile_16_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(533)
	);

	pe_tile pe_tile_16_21(
		.out_wire_3_0(vertical_tile_16_21_to_tile_15_21_0),
		.out_wire_3_1(vertical_tile_16_21_to_tile_15_21_1),
		.out_wire_3_2(vertical_tile_16_21_to_tile_15_21_2),
		.out_wire_3_3(vertical_tile_16_21_to_tile_15_21_3),
		.in_wire_3_0(vertical_tile_15_21_to_tile_16_21_0),
		.in_wire_3_1(vertical_tile_15_21_to_tile_16_21_1),
		.in_wire_3_2(vertical_tile_15_21_to_tile_16_21_2),
		.in_wire_3_3(vertical_tile_15_21_to_tile_16_21_3),
		.out_wire_1_0(vertical_tile_16_21_to_tile_17_21_0),
		.out_wire_1_1(vertical_tile_16_21_to_tile_17_21_1),
		.out_wire_1_2(vertical_tile_16_21_to_tile_17_21_2),
		.out_wire_1_3(vertical_tile_16_21_to_tile_17_21_3),
		.in_wire_1_0(vertical_tile_17_21_to_tile_16_21_0),
		.in_wire_1_1(vertical_tile_17_21_to_tile_16_21_1),
		.in_wire_1_2(vertical_tile_17_21_to_tile_16_21_2),
		.in_wire_1_3(vertical_tile_17_21_to_tile_16_21_3),
		.out_wire_2_0(horizontal_tile_16_21_to_tile_16_20_0),
		.out_wire_2_1(horizontal_tile_16_21_to_tile_16_20_1),
		.out_wire_2_2(horizontal_tile_16_21_to_tile_16_20_2),
		.out_wire_2_3(horizontal_tile_16_21_to_tile_16_20_3),
		.in_wire_2_0(horizontal_tile_16_20_to_tile_16_21_0),
		.in_wire_2_1(horizontal_tile_16_20_to_tile_16_21_1),
		.in_wire_2_2(horizontal_tile_16_20_to_tile_16_21_2),
		.in_wire_2_3(horizontal_tile_16_20_to_tile_16_21_3),
		.out_wire_0_0(horizontal_tile_16_21_to_tile_16_22_0),
		.out_wire_0_1(horizontal_tile_16_21_to_tile_16_22_1),
		.out_wire_0_2(horizontal_tile_16_21_to_tile_16_22_2),
		.out_wire_0_3(horizontal_tile_16_21_to_tile_16_22_3),
		.in_wire_0_0(horizontal_tile_16_22_to_tile_16_21_0),
		.in_wire_0_1(horizontal_tile_16_22_to_tile_16_21_1),
		.in_wire_0_2(horizontal_tile_16_22_to_tile_16_21_2),
		.in_wire_0_3(horizontal_tile_16_22_to_tile_16_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(534)
	);

	pe_tile pe_tile_16_22(
		.out_wire_3_0(vertical_tile_16_22_to_tile_15_22_0),
		.out_wire_3_1(vertical_tile_16_22_to_tile_15_22_1),
		.out_wire_3_2(vertical_tile_16_22_to_tile_15_22_2),
		.out_wire_3_3(vertical_tile_16_22_to_tile_15_22_3),
		.in_wire_3_0(vertical_tile_15_22_to_tile_16_22_0),
		.in_wire_3_1(vertical_tile_15_22_to_tile_16_22_1),
		.in_wire_3_2(vertical_tile_15_22_to_tile_16_22_2),
		.in_wire_3_3(vertical_tile_15_22_to_tile_16_22_3),
		.out_wire_1_0(vertical_tile_16_22_to_tile_17_22_0),
		.out_wire_1_1(vertical_tile_16_22_to_tile_17_22_1),
		.out_wire_1_2(vertical_tile_16_22_to_tile_17_22_2),
		.out_wire_1_3(vertical_tile_16_22_to_tile_17_22_3),
		.in_wire_1_0(vertical_tile_17_22_to_tile_16_22_0),
		.in_wire_1_1(vertical_tile_17_22_to_tile_16_22_1),
		.in_wire_1_2(vertical_tile_17_22_to_tile_16_22_2),
		.in_wire_1_3(vertical_tile_17_22_to_tile_16_22_3),
		.out_wire_2_0(horizontal_tile_16_22_to_tile_16_21_0),
		.out_wire_2_1(horizontal_tile_16_22_to_tile_16_21_1),
		.out_wire_2_2(horizontal_tile_16_22_to_tile_16_21_2),
		.out_wire_2_3(horizontal_tile_16_22_to_tile_16_21_3),
		.in_wire_2_0(horizontal_tile_16_21_to_tile_16_22_0),
		.in_wire_2_1(horizontal_tile_16_21_to_tile_16_22_1),
		.in_wire_2_2(horizontal_tile_16_21_to_tile_16_22_2),
		.in_wire_2_3(horizontal_tile_16_21_to_tile_16_22_3),
		.out_wire_0_0(horizontal_tile_16_22_to_tile_16_23_0),
		.out_wire_0_1(horizontal_tile_16_22_to_tile_16_23_1),
		.out_wire_0_2(horizontal_tile_16_22_to_tile_16_23_2),
		.out_wire_0_3(horizontal_tile_16_22_to_tile_16_23_3),
		.in_wire_0_0(horizontal_tile_16_23_to_tile_16_22_0),
		.in_wire_0_1(horizontal_tile_16_23_to_tile_16_22_1),
		.in_wire_0_2(horizontal_tile_16_23_to_tile_16_22_2),
		.in_wire_0_3(horizontal_tile_16_23_to_tile_16_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(535)
	);

	pe_tile pe_tile_16_23(
		.out_wire_3_0(vertical_tile_16_23_to_tile_15_23_0),
		.out_wire_3_1(vertical_tile_16_23_to_tile_15_23_1),
		.out_wire_3_2(vertical_tile_16_23_to_tile_15_23_2),
		.out_wire_3_3(vertical_tile_16_23_to_tile_15_23_3),
		.in_wire_3_0(vertical_tile_15_23_to_tile_16_23_0),
		.in_wire_3_1(vertical_tile_15_23_to_tile_16_23_1),
		.in_wire_3_2(vertical_tile_15_23_to_tile_16_23_2),
		.in_wire_3_3(vertical_tile_15_23_to_tile_16_23_3),
		.out_wire_1_0(vertical_tile_16_23_to_tile_17_23_0),
		.out_wire_1_1(vertical_tile_16_23_to_tile_17_23_1),
		.out_wire_1_2(vertical_tile_16_23_to_tile_17_23_2),
		.out_wire_1_3(vertical_tile_16_23_to_tile_17_23_3),
		.in_wire_1_0(vertical_tile_17_23_to_tile_16_23_0),
		.in_wire_1_1(vertical_tile_17_23_to_tile_16_23_1),
		.in_wire_1_2(vertical_tile_17_23_to_tile_16_23_2),
		.in_wire_1_3(vertical_tile_17_23_to_tile_16_23_3),
		.out_wire_2_0(horizontal_tile_16_23_to_tile_16_22_0),
		.out_wire_2_1(horizontal_tile_16_23_to_tile_16_22_1),
		.out_wire_2_2(horizontal_tile_16_23_to_tile_16_22_2),
		.out_wire_2_3(horizontal_tile_16_23_to_tile_16_22_3),
		.in_wire_2_0(horizontal_tile_16_22_to_tile_16_23_0),
		.in_wire_2_1(horizontal_tile_16_22_to_tile_16_23_1),
		.in_wire_2_2(horizontal_tile_16_22_to_tile_16_23_2),
		.in_wire_2_3(horizontal_tile_16_22_to_tile_16_23_3),
		.out_wire_0_0(horizontal_tile_16_23_to_tile_16_24_0),
		.out_wire_0_1(horizontal_tile_16_23_to_tile_16_24_1),
		.out_wire_0_2(horizontal_tile_16_23_to_tile_16_24_2),
		.out_wire_0_3(horizontal_tile_16_23_to_tile_16_24_3),
		.in_wire_0_0(horizontal_tile_16_24_to_tile_16_23_0),
		.in_wire_0_1(horizontal_tile_16_24_to_tile_16_23_1),
		.in_wire_0_2(horizontal_tile_16_24_to_tile_16_23_2),
		.in_wire_0_3(horizontal_tile_16_24_to_tile_16_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(536)
	);

	pe_tile pe_tile_16_24(
		.out_wire_3_0(vertical_tile_16_24_to_tile_15_24_0),
		.out_wire_3_1(vertical_tile_16_24_to_tile_15_24_1),
		.out_wire_3_2(vertical_tile_16_24_to_tile_15_24_2),
		.out_wire_3_3(vertical_tile_16_24_to_tile_15_24_3),
		.in_wire_3_0(vertical_tile_15_24_to_tile_16_24_0),
		.in_wire_3_1(vertical_tile_15_24_to_tile_16_24_1),
		.in_wire_3_2(vertical_tile_15_24_to_tile_16_24_2),
		.in_wire_3_3(vertical_tile_15_24_to_tile_16_24_3),
		.out_wire_1_0(vertical_tile_16_24_to_tile_17_24_0),
		.out_wire_1_1(vertical_tile_16_24_to_tile_17_24_1),
		.out_wire_1_2(vertical_tile_16_24_to_tile_17_24_2),
		.out_wire_1_3(vertical_tile_16_24_to_tile_17_24_3),
		.in_wire_1_0(vertical_tile_17_24_to_tile_16_24_0),
		.in_wire_1_1(vertical_tile_17_24_to_tile_16_24_1),
		.in_wire_1_2(vertical_tile_17_24_to_tile_16_24_2),
		.in_wire_1_3(vertical_tile_17_24_to_tile_16_24_3),
		.out_wire_2_0(horizontal_tile_16_24_to_tile_16_23_0),
		.out_wire_2_1(horizontal_tile_16_24_to_tile_16_23_1),
		.out_wire_2_2(horizontal_tile_16_24_to_tile_16_23_2),
		.out_wire_2_3(horizontal_tile_16_24_to_tile_16_23_3),
		.in_wire_2_0(horizontal_tile_16_23_to_tile_16_24_0),
		.in_wire_2_1(horizontal_tile_16_23_to_tile_16_24_1),
		.in_wire_2_2(horizontal_tile_16_23_to_tile_16_24_2),
		.in_wire_2_3(horizontal_tile_16_23_to_tile_16_24_3),
		.out_wire_0_0(horizontal_tile_16_24_to_tile_16_25_0),
		.out_wire_0_1(horizontal_tile_16_24_to_tile_16_25_1),
		.out_wire_0_2(horizontal_tile_16_24_to_tile_16_25_2),
		.out_wire_0_3(horizontal_tile_16_24_to_tile_16_25_3),
		.in_wire_0_0(horizontal_tile_16_25_to_tile_16_24_0),
		.in_wire_0_1(horizontal_tile_16_25_to_tile_16_24_1),
		.in_wire_0_2(horizontal_tile_16_25_to_tile_16_24_2),
		.in_wire_0_3(horizontal_tile_16_25_to_tile_16_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(537)
	);

	pe_tile pe_tile_16_25(
		.out_wire_3_0(vertical_tile_16_25_to_tile_15_25_0),
		.out_wire_3_1(vertical_tile_16_25_to_tile_15_25_1),
		.out_wire_3_2(vertical_tile_16_25_to_tile_15_25_2),
		.out_wire_3_3(vertical_tile_16_25_to_tile_15_25_3),
		.in_wire_3_0(vertical_tile_15_25_to_tile_16_25_0),
		.in_wire_3_1(vertical_tile_15_25_to_tile_16_25_1),
		.in_wire_3_2(vertical_tile_15_25_to_tile_16_25_2),
		.in_wire_3_3(vertical_tile_15_25_to_tile_16_25_3),
		.out_wire_1_0(vertical_tile_16_25_to_tile_17_25_0),
		.out_wire_1_1(vertical_tile_16_25_to_tile_17_25_1),
		.out_wire_1_2(vertical_tile_16_25_to_tile_17_25_2),
		.out_wire_1_3(vertical_tile_16_25_to_tile_17_25_3),
		.in_wire_1_0(vertical_tile_17_25_to_tile_16_25_0),
		.in_wire_1_1(vertical_tile_17_25_to_tile_16_25_1),
		.in_wire_1_2(vertical_tile_17_25_to_tile_16_25_2),
		.in_wire_1_3(vertical_tile_17_25_to_tile_16_25_3),
		.out_wire_2_0(horizontal_tile_16_25_to_tile_16_24_0),
		.out_wire_2_1(horizontal_tile_16_25_to_tile_16_24_1),
		.out_wire_2_2(horizontal_tile_16_25_to_tile_16_24_2),
		.out_wire_2_3(horizontal_tile_16_25_to_tile_16_24_3),
		.in_wire_2_0(horizontal_tile_16_24_to_tile_16_25_0),
		.in_wire_2_1(horizontal_tile_16_24_to_tile_16_25_1),
		.in_wire_2_2(horizontal_tile_16_24_to_tile_16_25_2),
		.in_wire_2_3(horizontal_tile_16_24_to_tile_16_25_3),
		.out_wire_0_0(horizontal_tile_16_25_to_tile_16_26_0),
		.out_wire_0_1(horizontal_tile_16_25_to_tile_16_26_1),
		.out_wire_0_2(horizontal_tile_16_25_to_tile_16_26_2),
		.out_wire_0_3(horizontal_tile_16_25_to_tile_16_26_3),
		.in_wire_0_0(horizontal_tile_16_26_to_tile_16_25_0),
		.in_wire_0_1(horizontal_tile_16_26_to_tile_16_25_1),
		.in_wire_0_2(horizontal_tile_16_26_to_tile_16_25_2),
		.in_wire_0_3(horizontal_tile_16_26_to_tile_16_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(538)
	);

	pe_tile pe_tile_16_26(
		.out_wire_3_0(vertical_tile_16_26_to_tile_15_26_0),
		.out_wire_3_1(vertical_tile_16_26_to_tile_15_26_1),
		.out_wire_3_2(vertical_tile_16_26_to_tile_15_26_2),
		.out_wire_3_3(vertical_tile_16_26_to_tile_15_26_3),
		.in_wire_3_0(vertical_tile_15_26_to_tile_16_26_0),
		.in_wire_3_1(vertical_tile_15_26_to_tile_16_26_1),
		.in_wire_3_2(vertical_tile_15_26_to_tile_16_26_2),
		.in_wire_3_3(vertical_tile_15_26_to_tile_16_26_3),
		.out_wire_1_0(vertical_tile_16_26_to_tile_17_26_0),
		.out_wire_1_1(vertical_tile_16_26_to_tile_17_26_1),
		.out_wire_1_2(vertical_tile_16_26_to_tile_17_26_2),
		.out_wire_1_3(vertical_tile_16_26_to_tile_17_26_3),
		.in_wire_1_0(vertical_tile_17_26_to_tile_16_26_0),
		.in_wire_1_1(vertical_tile_17_26_to_tile_16_26_1),
		.in_wire_1_2(vertical_tile_17_26_to_tile_16_26_2),
		.in_wire_1_3(vertical_tile_17_26_to_tile_16_26_3),
		.out_wire_2_0(horizontal_tile_16_26_to_tile_16_25_0),
		.out_wire_2_1(horizontal_tile_16_26_to_tile_16_25_1),
		.out_wire_2_2(horizontal_tile_16_26_to_tile_16_25_2),
		.out_wire_2_3(horizontal_tile_16_26_to_tile_16_25_3),
		.in_wire_2_0(horizontal_tile_16_25_to_tile_16_26_0),
		.in_wire_2_1(horizontal_tile_16_25_to_tile_16_26_1),
		.in_wire_2_2(horizontal_tile_16_25_to_tile_16_26_2),
		.in_wire_2_3(horizontal_tile_16_25_to_tile_16_26_3),
		.out_wire_0_0(horizontal_tile_16_26_to_tile_16_27_0),
		.out_wire_0_1(horizontal_tile_16_26_to_tile_16_27_1),
		.out_wire_0_2(horizontal_tile_16_26_to_tile_16_27_2),
		.out_wire_0_3(horizontal_tile_16_26_to_tile_16_27_3),
		.in_wire_0_0(horizontal_tile_16_27_to_tile_16_26_0),
		.in_wire_0_1(horizontal_tile_16_27_to_tile_16_26_1),
		.in_wire_0_2(horizontal_tile_16_27_to_tile_16_26_2),
		.in_wire_0_3(horizontal_tile_16_27_to_tile_16_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(539)
	);

	pe_tile pe_tile_16_27(
		.out_wire_3_0(vertical_tile_16_27_to_tile_15_27_0),
		.out_wire_3_1(vertical_tile_16_27_to_tile_15_27_1),
		.out_wire_3_2(vertical_tile_16_27_to_tile_15_27_2),
		.out_wire_3_3(vertical_tile_16_27_to_tile_15_27_3),
		.in_wire_3_0(vertical_tile_15_27_to_tile_16_27_0),
		.in_wire_3_1(vertical_tile_15_27_to_tile_16_27_1),
		.in_wire_3_2(vertical_tile_15_27_to_tile_16_27_2),
		.in_wire_3_3(vertical_tile_15_27_to_tile_16_27_3),
		.out_wire_1_0(vertical_tile_16_27_to_tile_17_27_0),
		.out_wire_1_1(vertical_tile_16_27_to_tile_17_27_1),
		.out_wire_1_2(vertical_tile_16_27_to_tile_17_27_2),
		.out_wire_1_3(vertical_tile_16_27_to_tile_17_27_3),
		.in_wire_1_0(vertical_tile_17_27_to_tile_16_27_0),
		.in_wire_1_1(vertical_tile_17_27_to_tile_16_27_1),
		.in_wire_1_2(vertical_tile_17_27_to_tile_16_27_2),
		.in_wire_1_3(vertical_tile_17_27_to_tile_16_27_3),
		.out_wire_2_0(horizontal_tile_16_27_to_tile_16_26_0),
		.out_wire_2_1(horizontal_tile_16_27_to_tile_16_26_1),
		.out_wire_2_2(horizontal_tile_16_27_to_tile_16_26_2),
		.out_wire_2_3(horizontal_tile_16_27_to_tile_16_26_3),
		.in_wire_2_0(horizontal_tile_16_26_to_tile_16_27_0),
		.in_wire_2_1(horizontal_tile_16_26_to_tile_16_27_1),
		.in_wire_2_2(horizontal_tile_16_26_to_tile_16_27_2),
		.in_wire_2_3(horizontal_tile_16_26_to_tile_16_27_3),
		.out_wire_0_0(horizontal_tile_16_27_to_tile_16_28_0),
		.out_wire_0_1(horizontal_tile_16_27_to_tile_16_28_1),
		.out_wire_0_2(horizontal_tile_16_27_to_tile_16_28_2),
		.out_wire_0_3(horizontal_tile_16_27_to_tile_16_28_3),
		.in_wire_0_0(horizontal_tile_16_28_to_tile_16_27_0),
		.in_wire_0_1(horizontal_tile_16_28_to_tile_16_27_1),
		.in_wire_0_2(horizontal_tile_16_28_to_tile_16_27_2),
		.in_wire_0_3(horizontal_tile_16_28_to_tile_16_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(540)
	);

	pe_tile pe_tile_16_28(
		.out_wire_3_0(vertical_tile_16_28_to_tile_15_28_0),
		.out_wire_3_1(vertical_tile_16_28_to_tile_15_28_1),
		.out_wire_3_2(vertical_tile_16_28_to_tile_15_28_2),
		.out_wire_3_3(vertical_tile_16_28_to_tile_15_28_3),
		.in_wire_3_0(vertical_tile_15_28_to_tile_16_28_0),
		.in_wire_3_1(vertical_tile_15_28_to_tile_16_28_1),
		.in_wire_3_2(vertical_tile_15_28_to_tile_16_28_2),
		.in_wire_3_3(vertical_tile_15_28_to_tile_16_28_3),
		.out_wire_1_0(vertical_tile_16_28_to_tile_17_28_0),
		.out_wire_1_1(vertical_tile_16_28_to_tile_17_28_1),
		.out_wire_1_2(vertical_tile_16_28_to_tile_17_28_2),
		.out_wire_1_3(vertical_tile_16_28_to_tile_17_28_3),
		.in_wire_1_0(vertical_tile_17_28_to_tile_16_28_0),
		.in_wire_1_1(vertical_tile_17_28_to_tile_16_28_1),
		.in_wire_1_2(vertical_tile_17_28_to_tile_16_28_2),
		.in_wire_1_3(vertical_tile_17_28_to_tile_16_28_3),
		.out_wire_2_0(horizontal_tile_16_28_to_tile_16_27_0),
		.out_wire_2_1(horizontal_tile_16_28_to_tile_16_27_1),
		.out_wire_2_2(horizontal_tile_16_28_to_tile_16_27_2),
		.out_wire_2_3(horizontal_tile_16_28_to_tile_16_27_3),
		.in_wire_2_0(horizontal_tile_16_27_to_tile_16_28_0),
		.in_wire_2_1(horizontal_tile_16_27_to_tile_16_28_1),
		.in_wire_2_2(horizontal_tile_16_27_to_tile_16_28_2),
		.in_wire_2_3(horizontal_tile_16_27_to_tile_16_28_3),
		.out_wire_0_0(horizontal_tile_16_28_to_tile_16_29_0),
		.out_wire_0_1(horizontal_tile_16_28_to_tile_16_29_1),
		.out_wire_0_2(horizontal_tile_16_28_to_tile_16_29_2),
		.out_wire_0_3(horizontal_tile_16_28_to_tile_16_29_3),
		.in_wire_0_0(horizontal_tile_16_29_to_tile_16_28_0),
		.in_wire_0_1(horizontal_tile_16_29_to_tile_16_28_1),
		.in_wire_0_2(horizontal_tile_16_29_to_tile_16_28_2),
		.in_wire_0_3(horizontal_tile_16_29_to_tile_16_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(541)
	);

	pe_tile pe_tile_16_29(
		.out_wire_3_0(vertical_tile_16_29_to_tile_15_29_0),
		.out_wire_3_1(vertical_tile_16_29_to_tile_15_29_1),
		.out_wire_3_2(vertical_tile_16_29_to_tile_15_29_2),
		.out_wire_3_3(vertical_tile_16_29_to_tile_15_29_3),
		.in_wire_3_0(vertical_tile_15_29_to_tile_16_29_0),
		.in_wire_3_1(vertical_tile_15_29_to_tile_16_29_1),
		.in_wire_3_2(vertical_tile_15_29_to_tile_16_29_2),
		.in_wire_3_3(vertical_tile_15_29_to_tile_16_29_3),
		.out_wire_1_0(vertical_tile_16_29_to_tile_17_29_0),
		.out_wire_1_1(vertical_tile_16_29_to_tile_17_29_1),
		.out_wire_1_2(vertical_tile_16_29_to_tile_17_29_2),
		.out_wire_1_3(vertical_tile_16_29_to_tile_17_29_3),
		.in_wire_1_0(vertical_tile_17_29_to_tile_16_29_0),
		.in_wire_1_1(vertical_tile_17_29_to_tile_16_29_1),
		.in_wire_1_2(vertical_tile_17_29_to_tile_16_29_2),
		.in_wire_1_3(vertical_tile_17_29_to_tile_16_29_3),
		.out_wire_2_0(horizontal_tile_16_29_to_tile_16_28_0),
		.out_wire_2_1(horizontal_tile_16_29_to_tile_16_28_1),
		.out_wire_2_2(horizontal_tile_16_29_to_tile_16_28_2),
		.out_wire_2_3(horizontal_tile_16_29_to_tile_16_28_3),
		.in_wire_2_0(horizontal_tile_16_28_to_tile_16_29_0),
		.in_wire_2_1(horizontal_tile_16_28_to_tile_16_29_1),
		.in_wire_2_2(horizontal_tile_16_28_to_tile_16_29_2),
		.in_wire_2_3(horizontal_tile_16_28_to_tile_16_29_3),
		.out_wire_0_0(horizontal_tile_16_29_to_tile_16_30_0),
		.out_wire_0_1(horizontal_tile_16_29_to_tile_16_30_1),
		.out_wire_0_2(horizontal_tile_16_29_to_tile_16_30_2),
		.out_wire_0_3(horizontal_tile_16_29_to_tile_16_30_3),
		.in_wire_0_0(horizontal_tile_16_30_to_tile_16_29_0),
		.in_wire_0_1(horizontal_tile_16_30_to_tile_16_29_1),
		.in_wire_0_2(horizontal_tile_16_30_to_tile_16_29_2),
		.in_wire_0_3(horizontal_tile_16_30_to_tile_16_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(542)
	);

	pe_tile pe_tile_16_30(
		.out_wire_3_0(vertical_tile_16_30_to_tile_15_30_0),
		.out_wire_3_1(vertical_tile_16_30_to_tile_15_30_1),
		.out_wire_3_2(vertical_tile_16_30_to_tile_15_30_2),
		.out_wire_3_3(vertical_tile_16_30_to_tile_15_30_3),
		.in_wire_3_0(vertical_tile_15_30_to_tile_16_30_0),
		.in_wire_3_1(vertical_tile_15_30_to_tile_16_30_1),
		.in_wire_3_2(vertical_tile_15_30_to_tile_16_30_2),
		.in_wire_3_3(vertical_tile_15_30_to_tile_16_30_3),
		.out_wire_1_0(vertical_tile_16_30_to_tile_17_30_0),
		.out_wire_1_1(vertical_tile_16_30_to_tile_17_30_1),
		.out_wire_1_2(vertical_tile_16_30_to_tile_17_30_2),
		.out_wire_1_3(vertical_tile_16_30_to_tile_17_30_3),
		.in_wire_1_0(vertical_tile_17_30_to_tile_16_30_0),
		.in_wire_1_1(vertical_tile_17_30_to_tile_16_30_1),
		.in_wire_1_2(vertical_tile_17_30_to_tile_16_30_2),
		.in_wire_1_3(vertical_tile_17_30_to_tile_16_30_3),
		.out_wire_2_0(horizontal_tile_16_30_to_tile_16_29_0),
		.out_wire_2_1(horizontal_tile_16_30_to_tile_16_29_1),
		.out_wire_2_2(horizontal_tile_16_30_to_tile_16_29_2),
		.out_wire_2_3(horizontal_tile_16_30_to_tile_16_29_3),
		.in_wire_2_0(horizontal_tile_16_29_to_tile_16_30_0),
		.in_wire_2_1(horizontal_tile_16_29_to_tile_16_30_1),
		.in_wire_2_2(horizontal_tile_16_29_to_tile_16_30_2),
		.in_wire_2_3(horizontal_tile_16_29_to_tile_16_30_3),
		.out_wire_0_0(horizontal_tile_16_30_to_tile_16_31_0),
		.out_wire_0_1(horizontal_tile_16_30_to_tile_16_31_1),
		.out_wire_0_2(horizontal_tile_16_30_to_tile_16_31_2),
		.out_wire_0_3(horizontal_tile_16_30_to_tile_16_31_3),
		.in_wire_0_0(horizontal_tile_16_31_to_tile_16_30_0),
		.in_wire_0_1(horizontal_tile_16_31_to_tile_16_30_1),
		.in_wire_0_2(horizontal_tile_16_31_to_tile_16_30_2),
		.in_wire_0_3(horizontal_tile_16_31_to_tile_16_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(543)
	);

	pe_tile_right pe_tile_16_31(
		.out_wire_3_0(vertical_tile_16_31_to_tile_15_31_0),
		.out_wire_3_1(vertical_tile_16_31_to_tile_15_31_1),
		.out_wire_3_2(vertical_tile_16_31_to_tile_15_31_2),
		.out_wire_3_3(vertical_tile_16_31_to_tile_15_31_3),
		.in_wire_3_0(vertical_tile_15_31_to_tile_16_31_0),
		.in_wire_3_1(vertical_tile_15_31_to_tile_16_31_1),
		.in_wire_3_2(vertical_tile_15_31_to_tile_16_31_2),
		.in_wire_3_3(vertical_tile_15_31_to_tile_16_31_3),
		.out_wire_1_0(vertical_tile_16_31_to_tile_17_31_0),
		.out_wire_1_1(vertical_tile_16_31_to_tile_17_31_1),
		.out_wire_1_2(vertical_tile_16_31_to_tile_17_31_2),
		.out_wire_1_3(vertical_tile_16_31_to_tile_17_31_3),
		.in_wire_1_0(vertical_tile_17_31_to_tile_16_31_0),
		.in_wire_1_1(vertical_tile_17_31_to_tile_16_31_1),
		.in_wire_1_2(vertical_tile_17_31_to_tile_16_31_2),
		.in_wire_1_3(vertical_tile_17_31_to_tile_16_31_3),
		.out_wire_2_0(horizontal_tile_16_31_to_tile_16_30_0),
		.out_wire_2_1(horizontal_tile_16_31_to_tile_16_30_1),
		.out_wire_2_2(horizontal_tile_16_31_to_tile_16_30_2),
		.out_wire_2_3(horizontal_tile_16_31_to_tile_16_30_3),
		.in_wire_2_0(horizontal_tile_16_30_to_tile_16_31_0),
		.in_wire_2_1(horizontal_tile_16_30_to_tile_16_31_1),
		.in_wire_2_2(horizontal_tile_16_30_to_tile_16_31_2),
		.in_wire_2_3(horizontal_tile_16_30_to_tile_16_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(544)
	);

	pe_tile_left pe_tile_17_0(
		.out_wire_3_0(vertical_tile_17_0_to_tile_16_0_0),
		.out_wire_3_1(vertical_tile_17_0_to_tile_16_0_1),
		.out_wire_3_2(vertical_tile_17_0_to_tile_16_0_2),
		.out_wire_3_3(vertical_tile_17_0_to_tile_16_0_3),
		.in_wire_3_0(vertical_tile_16_0_to_tile_17_0_0),
		.in_wire_3_1(vertical_tile_16_0_to_tile_17_0_1),
		.in_wire_3_2(vertical_tile_16_0_to_tile_17_0_2),
		.in_wire_3_3(vertical_tile_16_0_to_tile_17_0_3),
		.out_wire_1_0(vertical_tile_17_0_to_tile_18_0_0),
		.out_wire_1_1(vertical_tile_17_0_to_tile_18_0_1),
		.out_wire_1_2(vertical_tile_17_0_to_tile_18_0_2),
		.out_wire_1_3(vertical_tile_17_0_to_tile_18_0_3),
		.in_wire_1_0(vertical_tile_18_0_to_tile_17_0_0),
		.in_wire_1_1(vertical_tile_18_0_to_tile_17_0_1),
		.in_wire_1_2(vertical_tile_18_0_to_tile_17_0_2),
		.in_wire_1_3(vertical_tile_18_0_to_tile_17_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_17_0_to_tile_17_1_0),
		.out_wire_0_1(horizontal_tile_17_0_to_tile_17_1_1),
		.out_wire_0_2(horizontal_tile_17_0_to_tile_17_1_2),
		.out_wire_0_3(horizontal_tile_17_0_to_tile_17_1_3),
		.in_wire_0_0(horizontal_tile_17_1_to_tile_17_0_0),
		.in_wire_0_1(horizontal_tile_17_1_to_tile_17_0_1),
		.in_wire_0_2(horizontal_tile_17_1_to_tile_17_0_2),
		.in_wire_0_3(horizontal_tile_17_1_to_tile_17_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(545)
	);

	pe_tile pe_tile_17_1(
		.out_wire_3_0(vertical_tile_17_1_to_tile_16_1_0),
		.out_wire_3_1(vertical_tile_17_1_to_tile_16_1_1),
		.out_wire_3_2(vertical_tile_17_1_to_tile_16_1_2),
		.out_wire_3_3(vertical_tile_17_1_to_tile_16_1_3),
		.in_wire_3_0(vertical_tile_16_1_to_tile_17_1_0),
		.in_wire_3_1(vertical_tile_16_1_to_tile_17_1_1),
		.in_wire_3_2(vertical_tile_16_1_to_tile_17_1_2),
		.in_wire_3_3(vertical_tile_16_1_to_tile_17_1_3),
		.out_wire_1_0(vertical_tile_17_1_to_tile_18_1_0),
		.out_wire_1_1(vertical_tile_17_1_to_tile_18_1_1),
		.out_wire_1_2(vertical_tile_17_1_to_tile_18_1_2),
		.out_wire_1_3(vertical_tile_17_1_to_tile_18_1_3),
		.in_wire_1_0(vertical_tile_18_1_to_tile_17_1_0),
		.in_wire_1_1(vertical_tile_18_1_to_tile_17_1_1),
		.in_wire_1_2(vertical_tile_18_1_to_tile_17_1_2),
		.in_wire_1_3(vertical_tile_18_1_to_tile_17_1_3),
		.out_wire_2_0(horizontal_tile_17_1_to_tile_17_0_0),
		.out_wire_2_1(horizontal_tile_17_1_to_tile_17_0_1),
		.out_wire_2_2(horizontal_tile_17_1_to_tile_17_0_2),
		.out_wire_2_3(horizontal_tile_17_1_to_tile_17_0_3),
		.in_wire_2_0(horizontal_tile_17_0_to_tile_17_1_0),
		.in_wire_2_1(horizontal_tile_17_0_to_tile_17_1_1),
		.in_wire_2_2(horizontal_tile_17_0_to_tile_17_1_2),
		.in_wire_2_3(horizontal_tile_17_0_to_tile_17_1_3),
		.out_wire_0_0(horizontal_tile_17_1_to_tile_17_2_0),
		.out_wire_0_1(horizontal_tile_17_1_to_tile_17_2_1),
		.out_wire_0_2(horizontal_tile_17_1_to_tile_17_2_2),
		.out_wire_0_3(horizontal_tile_17_1_to_tile_17_2_3),
		.in_wire_0_0(horizontal_tile_17_2_to_tile_17_1_0),
		.in_wire_0_1(horizontal_tile_17_2_to_tile_17_1_1),
		.in_wire_0_2(horizontal_tile_17_2_to_tile_17_1_2),
		.in_wire_0_3(horizontal_tile_17_2_to_tile_17_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(546)
	);

	pe_tile pe_tile_17_2(
		.out_wire_3_0(vertical_tile_17_2_to_tile_16_2_0),
		.out_wire_3_1(vertical_tile_17_2_to_tile_16_2_1),
		.out_wire_3_2(vertical_tile_17_2_to_tile_16_2_2),
		.out_wire_3_3(vertical_tile_17_2_to_tile_16_2_3),
		.in_wire_3_0(vertical_tile_16_2_to_tile_17_2_0),
		.in_wire_3_1(vertical_tile_16_2_to_tile_17_2_1),
		.in_wire_3_2(vertical_tile_16_2_to_tile_17_2_2),
		.in_wire_3_3(vertical_tile_16_2_to_tile_17_2_3),
		.out_wire_1_0(vertical_tile_17_2_to_tile_18_2_0),
		.out_wire_1_1(vertical_tile_17_2_to_tile_18_2_1),
		.out_wire_1_2(vertical_tile_17_2_to_tile_18_2_2),
		.out_wire_1_3(vertical_tile_17_2_to_tile_18_2_3),
		.in_wire_1_0(vertical_tile_18_2_to_tile_17_2_0),
		.in_wire_1_1(vertical_tile_18_2_to_tile_17_2_1),
		.in_wire_1_2(vertical_tile_18_2_to_tile_17_2_2),
		.in_wire_1_3(vertical_tile_18_2_to_tile_17_2_3),
		.out_wire_2_0(horizontal_tile_17_2_to_tile_17_1_0),
		.out_wire_2_1(horizontal_tile_17_2_to_tile_17_1_1),
		.out_wire_2_2(horizontal_tile_17_2_to_tile_17_1_2),
		.out_wire_2_3(horizontal_tile_17_2_to_tile_17_1_3),
		.in_wire_2_0(horizontal_tile_17_1_to_tile_17_2_0),
		.in_wire_2_1(horizontal_tile_17_1_to_tile_17_2_1),
		.in_wire_2_2(horizontal_tile_17_1_to_tile_17_2_2),
		.in_wire_2_3(horizontal_tile_17_1_to_tile_17_2_3),
		.out_wire_0_0(horizontal_tile_17_2_to_tile_17_3_0),
		.out_wire_0_1(horizontal_tile_17_2_to_tile_17_3_1),
		.out_wire_0_2(horizontal_tile_17_2_to_tile_17_3_2),
		.out_wire_0_3(horizontal_tile_17_2_to_tile_17_3_3),
		.in_wire_0_0(horizontal_tile_17_3_to_tile_17_2_0),
		.in_wire_0_1(horizontal_tile_17_3_to_tile_17_2_1),
		.in_wire_0_2(horizontal_tile_17_3_to_tile_17_2_2),
		.in_wire_0_3(horizontal_tile_17_3_to_tile_17_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(547)
	);

	pe_tile pe_tile_17_3(
		.out_wire_3_0(vertical_tile_17_3_to_tile_16_3_0),
		.out_wire_3_1(vertical_tile_17_3_to_tile_16_3_1),
		.out_wire_3_2(vertical_tile_17_3_to_tile_16_3_2),
		.out_wire_3_3(vertical_tile_17_3_to_tile_16_3_3),
		.in_wire_3_0(vertical_tile_16_3_to_tile_17_3_0),
		.in_wire_3_1(vertical_tile_16_3_to_tile_17_3_1),
		.in_wire_3_2(vertical_tile_16_3_to_tile_17_3_2),
		.in_wire_3_3(vertical_tile_16_3_to_tile_17_3_3),
		.out_wire_1_0(vertical_tile_17_3_to_tile_18_3_0),
		.out_wire_1_1(vertical_tile_17_3_to_tile_18_3_1),
		.out_wire_1_2(vertical_tile_17_3_to_tile_18_3_2),
		.out_wire_1_3(vertical_tile_17_3_to_tile_18_3_3),
		.in_wire_1_0(vertical_tile_18_3_to_tile_17_3_0),
		.in_wire_1_1(vertical_tile_18_3_to_tile_17_3_1),
		.in_wire_1_2(vertical_tile_18_3_to_tile_17_3_2),
		.in_wire_1_3(vertical_tile_18_3_to_tile_17_3_3),
		.out_wire_2_0(horizontal_tile_17_3_to_tile_17_2_0),
		.out_wire_2_1(horizontal_tile_17_3_to_tile_17_2_1),
		.out_wire_2_2(horizontal_tile_17_3_to_tile_17_2_2),
		.out_wire_2_3(horizontal_tile_17_3_to_tile_17_2_3),
		.in_wire_2_0(horizontal_tile_17_2_to_tile_17_3_0),
		.in_wire_2_1(horizontal_tile_17_2_to_tile_17_3_1),
		.in_wire_2_2(horizontal_tile_17_2_to_tile_17_3_2),
		.in_wire_2_3(horizontal_tile_17_2_to_tile_17_3_3),
		.out_wire_0_0(horizontal_tile_17_3_to_tile_17_4_0),
		.out_wire_0_1(horizontal_tile_17_3_to_tile_17_4_1),
		.out_wire_0_2(horizontal_tile_17_3_to_tile_17_4_2),
		.out_wire_0_3(horizontal_tile_17_3_to_tile_17_4_3),
		.in_wire_0_0(horizontal_tile_17_4_to_tile_17_3_0),
		.in_wire_0_1(horizontal_tile_17_4_to_tile_17_3_1),
		.in_wire_0_2(horizontal_tile_17_4_to_tile_17_3_2),
		.in_wire_0_3(horizontal_tile_17_4_to_tile_17_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(548)
	);

	pe_tile pe_tile_17_4(
		.out_wire_3_0(vertical_tile_17_4_to_tile_16_4_0),
		.out_wire_3_1(vertical_tile_17_4_to_tile_16_4_1),
		.out_wire_3_2(vertical_tile_17_4_to_tile_16_4_2),
		.out_wire_3_3(vertical_tile_17_4_to_tile_16_4_3),
		.in_wire_3_0(vertical_tile_16_4_to_tile_17_4_0),
		.in_wire_3_1(vertical_tile_16_4_to_tile_17_4_1),
		.in_wire_3_2(vertical_tile_16_4_to_tile_17_4_2),
		.in_wire_3_3(vertical_tile_16_4_to_tile_17_4_3),
		.out_wire_1_0(vertical_tile_17_4_to_tile_18_4_0),
		.out_wire_1_1(vertical_tile_17_4_to_tile_18_4_1),
		.out_wire_1_2(vertical_tile_17_4_to_tile_18_4_2),
		.out_wire_1_3(vertical_tile_17_4_to_tile_18_4_3),
		.in_wire_1_0(vertical_tile_18_4_to_tile_17_4_0),
		.in_wire_1_1(vertical_tile_18_4_to_tile_17_4_1),
		.in_wire_1_2(vertical_tile_18_4_to_tile_17_4_2),
		.in_wire_1_3(vertical_tile_18_4_to_tile_17_4_3),
		.out_wire_2_0(horizontal_tile_17_4_to_tile_17_3_0),
		.out_wire_2_1(horizontal_tile_17_4_to_tile_17_3_1),
		.out_wire_2_2(horizontal_tile_17_4_to_tile_17_3_2),
		.out_wire_2_3(horizontal_tile_17_4_to_tile_17_3_3),
		.in_wire_2_0(horizontal_tile_17_3_to_tile_17_4_0),
		.in_wire_2_1(horizontal_tile_17_3_to_tile_17_4_1),
		.in_wire_2_2(horizontal_tile_17_3_to_tile_17_4_2),
		.in_wire_2_3(horizontal_tile_17_3_to_tile_17_4_3),
		.out_wire_0_0(horizontal_tile_17_4_to_tile_17_5_0),
		.out_wire_0_1(horizontal_tile_17_4_to_tile_17_5_1),
		.out_wire_0_2(horizontal_tile_17_4_to_tile_17_5_2),
		.out_wire_0_3(horizontal_tile_17_4_to_tile_17_5_3),
		.in_wire_0_0(horizontal_tile_17_5_to_tile_17_4_0),
		.in_wire_0_1(horizontal_tile_17_5_to_tile_17_4_1),
		.in_wire_0_2(horizontal_tile_17_5_to_tile_17_4_2),
		.in_wire_0_3(horizontal_tile_17_5_to_tile_17_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(549)
	);

	pe_tile pe_tile_17_5(
		.out_wire_3_0(vertical_tile_17_5_to_tile_16_5_0),
		.out_wire_3_1(vertical_tile_17_5_to_tile_16_5_1),
		.out_wire_3_2(vertical_tile_17_5_to_tile_16_5_2),
		.out_wire_3_3(vertical_tile_17_5_to_tile_16_5_3),
		.in_wire_3_0(vertical_tile_16_5_to_tile_17_5_0),
		.in_wire_3_1(vertical_tile_16_5_to_tile_17_5_1),
		.in_wire_3_2(vertical_tile_16_5_to_tile_17_5_2),
		.in_wire_3_3(vertical_tile_16_5_to_tile_17_5_3),
		.out_wire_1_0(vertical_tile_17_5_to_tile_18_5_0),
		.out_wire_1_1(vertical_tile_17_5_to_tile_18_5_1),
		.out_wire_1_2(vertical_tile_17_5_to_tile_18_5_2),
		.out_wire_1_3(vertical_tile_17_5_to_tile_18_5_3),
		.in_wire_1_0(vertical_tile_18_5_to_tile_17_5_0),
		.in_wire_1_1(vertical_tile_18_5_to_tile_17_5_1),
		.in_wire_1_2(vertical_tile_18_5_to_tile_17_5_2),
		.in_wire_1_3(vertical_tile_18_5_to_tile_17_5_3),
		.out_wire_2_0(horizontal_tile_17_5_to_tile_17_4_0),
		.out_wire_2_1(horizontal_tile_17_5_to_tile_17_4_1),
		.out_wire_2_2(horizontal_tile_17_5_to_tile_17_4_2),
		.out_wire_2_3(horizontal_tile_17_5_to_tile_17_4_3),
		.in_wire_2_0(horizontal_tile_17_4_to_tile_17_5_0),
		.in_wire_2_1(horizontal_tile_17_4_to_tile_17_5_1),
		.in_wire_2_2(horizontal_tile_17_4_to_tile_17_5_2),
		.in_wire_2_3(horizontal_tile_17_4_to_tile_17_5_3),
		.out_wire_0_0(horizontal_tile_17_5_to_tile_17_6_0),
		.out_wire_0_1(horizontal_tile_17_5_to_tile_17_6_1),
		.out_wire_0_2(horizontal_tile_17_5_to_tile_17_6_2),
		.out_wire_0_3(horizontal_tile_17_5_to_tile_17_6_3),
		.in_wire_0_0(horizontal_tile_17_6_to_tile_17_5_0),
		.in_wire_0_1(horizontal_tile_17_6_to_tile_17_5_1),
		.in_wire_0_2(horizontal_tile_17_6_to_tile_17_5_2),
		.in_wire_0_3(horizontal_tile_17_6_to_tile_17_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(550)
	);

	pe_tile pe_tile_17_6(
		.out_wire_3_0(vertical_tile_17_6_to_tile_16_6_0),
		.out_wire_3_1(vertical_tile_17_6_to_tile_16_6_1),
		.out_wire_3_2(vertical_tile_17_6_to_tile_16_6_2),
		.out_wire_3_3(vertical_tile_17_6_to_tile_16_6_3),
		.in_wire_3_0(vertical_tile_16_6_to_tile_17_6_0),
		.in_wire_3_1(vertical_tile_16_6_to_tile_17_6_1),
		.in_wire_3_2(vertical_tile_16_6_to_tile_17_6_2),
		.in_wire_3_3(vertical_tile_16_6_to_tile_17_6_3),
		.out_wire_1_0(vertical_tile_17_6_to_tile_18_6_0),
		.out_wire_1_1(vertical_tile_17_6_to_tile_18_6_1),
		.out_wire_1_2(vertical_tile_17_6_to_tile_18_6_2),
		.out_wire_1_3(vertical_tile_17_6_to_tile_18_6_3),
		.in_wire_1_0(vertical_tile_18_6_to_tile_17_6_0),
		.in_wire_1_1(vertical_tile_18_6_to_tile_17_6_1),
		.in_wire_1_2(vertical_tile_18_6_to_tile_17_6_2),
		.in_wire_1_3(vertical_tile_18_6_to_tile_17_6_3),
		.out_wire_2_0(horizontal_tile_17_6_to_tile_17_5_0),
		.out_wire_2_1(horizontal_tile_17_6_to_tile_17_5_1),
		.out_wire_2_2(horizontal_tile_17_6_to_tile_17_5_2),
		.out_wire_2_3(horizontal_tile_17_6_to_tile_17_5_3),
		.in_wire_2_0(horizontal_tile_17_5_to_tile_17_6_0),
		.in_wire_2_1(horizontal_tile_17_5_to_tile_17_6_1),
		.in_wire_2_2(horizontal_tile_17_5_to_tile_17_6_2),
		.in_wire_2_3(horizontal_tile_17_5_to_tile_17_6_3),
		.out_wire_0_0(horizontal_tile_17_6_to_tile_17_7_0),
		.out_wire_0_1(horizontal_tile_17_6_to_tile_17_7_1),
		.out_wire_0_2(horizontal_tile_17_6_to_tile_17_7_2),
		.out_wire_0_3(horizontal_tile_17_6_to_tile_17_7_3),
		.in_wire_0_0(horizontal_tile_17_7_to_tile_17_6_0),
		.in_wire_0_1(horizontal_tile_17_7_to_tile_17_6_1),
		.in_wire_0_2(horizontal_tile_17_7_to_tile_17_6_2),
		.in_wire_0_3(horizontal_tile_17_7_to_tile_17_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(551)
	);

	pe_tile pe_tile_17_7(
		.out_wire_3_0(vertical_tile_17_7_to_tile_16_7_0),
		.out_wire_3_1(vertical_tile_17_7_to_tile_16_7_1),
		.out_wire_3_2(vertical_tile_17_7_to_tile_16_7_2),
		.out_wire_3_3(vertical_tile_17_7_to_tile_16_7_3),
		.in_wire_3_0(vertical_tile_16_7_to_tile_17_7_0),
		.in_wire_3_1(vertical_tile_16_7_to_tile_17_7_1),
		.in_wire_3_2(vertical_tile_16_7_to_tile_17_7_2),
		.in_wire_3_3(vertical_tile_16_7_to_tile_17_7_3),
		.out_wire_1_0(vertical_tile_17_7_to_tile_18_7_0),
		.out_wire_1_1(vertical_tile_17_7_to_tile_18_7_1),
		.out_wire_1_2(vertical_tile_17_7_to_tile_18_7_2),
		.out_wire_1_3(vertical_tile_17_7_to_tile_18_7_3),
		.in_wire_1_0(vertical_tile_18_7_to_tile_17_7_0),
		.in_wire_1_1(vertical_tile_18_7_to_tile_17_7_1),
		.in_wire_1_2(vertical_tile_18_7_to_tile_17_7_2),
		.in_wire_1_3(vertical_tile_18_7_to_tile_17_7_3),
		.out_wire_2_0(horizontal_tile_17_7_to_tile_17_6_0),
		.out_wire_2_1(horizontal_tile_17_7_to_tile_17_6_1),
		.out_wire_2_2(horizontal_tile_17_7_to_tile_17_6_2),
		.out_wire_2_3(horizontal_tile_17_7_to_tile_17_6_3),
		.in_wire_2_0(horizontal_tile_17_6_to_tile_17_7_0),
		.in_wire_2_1(horizontal_tile_17_6_to_tile_17_7_1),
		.in_wire_2_2(horizontal_tile_17_6_to_tile_17_7_2),
		.in_wire_2_3(horizontal_tile_17_6_to_tile_17_7_3),
		.out_wire_0_0(horizontal_tile_17_7_to_tile_17_8_0),
		.out_wire_0_1(horizontal_tile_17_7_to_tile_17_8_1),
		.out_wire_0_2(horizontal_tile_17_7_to_tile_17_8_2),
		.out_wire_0_3(horizontal_tile_17_7_to_tile_17_8_3),
		.in_wire_0_0(horizontal_tile_17_8_to_tile_17_7_0),
		.in_wire_0_1(horizontal_tile_17_8_to_tile_17_7_1),
		.in_wire_0_2(horizontal_tile_17_8_to_tile_17_7_2),
		.in_wire_0_3(horizontal_tile_17_8_to_tile_17_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(552)
	);

	pe_tile pe_tile_17_8(
		.out_wire_3_0(vertical_tile_17_8_to_tile_16_8_0),
		.out_wire_3_1(vertical_tile_17_8_to_tile_16_8_1),
		.out_wire_3_2(vertical_tile_17_8_to_tile_16_8_2),
		.out_wire_3_3(vertical_tile_17_8_to_tile_16_8_3),
		.in_wire_3_0(vertical_tile_16_8_to_tile_17_8_0),
		.in_wire_3_1(vertical_tile_16_8_to_tile_17_8_1),
		.in_wire_3_2(vertical_tile_16_8_to_tile_17_8_2),
		.in_wire_3_3(vertical_tile_16_8_to_tile_17_8_3),
		.out_wire_1_0(vertical_tile_17_8_to_tile_18_8_0),
		.out_wire_1_1(vertical_tile_17_8_to_tile_18_8_1),
		.out_wire_1_2(vertical_tile_17_8_to_tile_18_8_2),
		.out_wire_1_3(vertical_tile_17_8_to_tile_18_8_3),
		.in_wire_1_0(vertical_tile_18_8_to_tile_17_8_0),
		.in_wire_1_1(vertical_tile_18_8_to_tile_17_8_1),
		.in_wire_1_2(vertical_tile_18_8_to_tile_17_8_2),
		.in_wire_1_3(vertical_tile_18_8_to_tile_17_8_3),
		.out_wire_2_0(horizontal_tile_17_8_to_tile_17_7_0),
		.out_wire_2_1(horizontal_tile_17_8_to_tile_17_7_1),
		.out_wire_2_2(horizontal_tile_17_8_to_tile_17_7_2),
		.out_wire_2_3(horizontal_tile_17_8_to_tile_17_7_3),
		.in_wire_2_0(horizontal_tile_17_7_to_tile_17_8_0),
		.in_wire_2_1(horizontal_tile_17_7_to_tile_17_8_1),
		.in_wire_2_2(horizontal_tile_17_7_to_tile_17_8_2),
		.in_wire_2_3(horizontal_tile_17_7_to_tile_17_8_3),
		.out_wire_0_0(horizontal_tile_17_8_to_tile_17_9_0),
		.out_wire_0_1(horizontal_tile_17_8_to_tile_17_9_1),
		.out_wire_0_2(horizontal_tile_17_8_to_tile_17_9_2),
		.out_wire_0_3(horizontal_tile_17_8_to_tile_17_9_3),
		.in_wire_0_0(horizontal_tile_17_9_to_tile_17_8_0),
		.in_wire_0_1(horizontal_tile_17_9_to_tile_17_8_1),
		.in_wire_0_2(horizontal_tile_17_9_to_tile_17_8_2),
		.in_wire_0_3(horizontal_tile_17_9_to_tile_17_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(553)
	);

	pe_tile pe_tile_17_9(
		.out_wire_3_0(vertical_tile_17_9_to_tile_16_9_0),
		.out_wire_3_1(vertical_tile_17_9_to_tile_16_9_1),
		.out_wire_3_2(vertical_tile_17_9_to_tile_16_9_2),
		.out_wire_3_3(vertical_tile_17_9_to_tile_16_9_3),
		.in_wire_3_0(vertical_tile_16_9_to_tile_17_9_0),
		.in_wire_3_1(vertical_tile_16_9_to_tile_17_9_1),
		.in_wire_3_2(vertical_tile_16_9_to_tile_17_9_2),
		.in_wire_3_3(vertical_tile_16_9_to_tile_17_9_3),
		.out_wire_1_0(vertical_tile_17_9_to_tile_18_9_0),
		.out_wire_1_1(vertical_tile_17_9_to_tile_18_9_1),
		.out_wire_1_2(vertical_tile_17_9_to_tile_18_9_2),
		.out_wire_1_3(vertical_tile_17_9_to_tile_18_9_3),
		.in_wire_1_0(vertical_tile_18_9_to_tile_17_9_0),
		.in_wire_1_1(vertical_tile_18_9_to_tile_17_9_1),
		.in_wire_1_2(vertical_tile_18_9_to_tile_17_9_2),
		.in_wire_1_3(vertical_tile_18_9_to_tile_17_9_3),
		.out_wire_2_0(horizontal_tile_17_9_to_tile_17_8_0),
		.out_wire_2_1(horizontal_tile_17_9_to_tile_17_8_1),
		.out_wire_2_2(horizontal_tile_17_9_to_tile_17_8_2),
		.out_wire_2_3(horizontal_tile_17_9_to_tile_17_8_3),
		.in_wire_2_0(horizontal_tile_17_8_to_tile_17_9_0),
		.in_wire_2_1(horizontal_tile_17_8_to_tile_17_9_1),
		.in_wire_2_2(horizontal_tile_17_8_to_tile_17_9_2),
		.in_wire_2_3(horizontal_tile_17_8_to_tile_17_9_3),
		.out_wire_0_0(horizontal_tile_17_9_to_tile_17_10_0),
		.out_wire_0_1(horizontal_tile_17_9_to_tile_17_10_1),
		.out_wire_0_2(horizontal_tile_17_9_to_tile_17_10_2),
		.out_wire_0_3(horizontal_tile_17_9_to_tile_17_10_3),
		.in_wire_0_0(horizontal_tile_17_10_to_tile_17_9_0),
		.in_wire_0_1(horizontal_tile_17_10_to_tile_17_9_1),
		.in_wire_0_2(horizontal_tile_17_10_to_tile_17_9_2),
		.in_wire_0_3(horizontal_tile_17_10_to_tile_17_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(554)
	);

	pe_tile pe_tile_17_10(
		.out_wire_3_0(vertical_tile_17_10_to_tile_16_10_0),
		.out_wire_3_1(vertical_tile_17_10_to_tile_16_10_1),
		.out_wire_3_2(vertical_tile_17_10_to_tile_16_10_2),
		.out_wire_3_3(vertical_tile_17_10_to_tile_16_10_3),
		.in_wire_3_0(vertical_tile_16_10_to_tile_17_10_0),
		.in_wire_3_1(vertical_tile_16_10_to_tile_17_10_1),
		.in_wire_3_2(vertical_tile_16_10_to_tile_17_10_2),
		.in_wire_3_3(vertical_tile_16_10_to_tile_17_10_3),
		.out_wire_1_0(vertical_tile_17_10_to_tile_18_10_0),
		.out_wire_1_1(vertical_tile_17_10_to_tile_18_10_1),
		.out_wire_1_2(vertical_tile_17_10_to_tile_18_10_2),
		.out_wire_1_3(vertical_tile_17_10_to_tile_18_10_3),
		.in_wire_1_0(vertical_tile_18_10_to_tile_17_10_0),
		.in_wire_1_1(vertical_tile_18_10_to_tile_17_10_1),
		.in_wire_1_2(vertical_tile_18_10_to_tile_17_10_2),
		.in_wire_1_3(vertical_tile_18_10_to_tile_17_10_3),
		.out_wire_2_0(horizontal_tile_17_10_to_tile_17_9_0),
		.out_wire_2_1(horizontal_tile_17_10_to_tile_17_9_1),
		.out_wire_2_2(horizontal_tile_17_10_to_tile_17_9_2),
		.out_wire_2_3(horizontal_tile_17_10_to_tile_17_9_3),
		.in_wire_2_0(horizontal_tile_17_9_to_tile_17_10_0),
		.in_wire_2_1(horizontal_tile_17_9_to_tile_17_10_1),
		.in_wire_2_2(horizontal_tile_17_9_to_tile_17_10_2),
		.in_wire_2_3(horizontal_tile_17_9_to_tile_17_10_3),
		.out_wire_0_0(horizontal_tile_17_10_to_tile_17_11_0),
		.out_wire_0_1(horizontal_tile_17_10_to_tile_17_11_1),
		.out_wire_0_2(horizontal_tile_17_10_to_tile_17_11_2),
		.out_wire_0_3(horizontal_tile_17_10_to_tile_17_11_3),
		.in_wire_0_0(horizontal_tile_17_11_to_tile_17_10_0),
		.in_wire_0_1(horizontal_tile_17_11_to_tile_17_10_1),
		.in_wire_0_2(horizontal_tile_17_11_to_tile_17_10_2),
		.in_wire_0_3(horizontal_tile_17_11_to_tile_17_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(555)
	);

	pe_tile pe_tile_17_11(
		.out_wire_3_0(vertical_tile_17_11_to_tile_16_11_0),
		.out_wire_3_1(vertical_tile_17_11_to_tile_16_11_1),
		.out_wire_3_2(vertical_tile_17_11_to_tile_16_11_2),
		.out_wire_3_3(vertical_tile_17_11_to_tile_16_11_3),
		.in_wire_3_0(vertical_tile_16_11_to_tile_17_11_0),
		.in_wire_3_1(vertical_tile_16_11_to_tile_17_11_1),
		.in_wire_3_2(vertical_tile_16_11_to_tile_17_11_2),
		.in_wire_3_3(vertical_tile_16_11_to_tile_17_11_3),
		.out_wire_1_0(vertical_tile_17_11_to_tile_18_11_0),
		.out_wire_1_1(vertical_tile_17_11_to_tile_18_11_1),
		.out_wire_1_2(vertical_tile_17_11_to_tile_18_11_2),
		.out_wire_1_3(vertical_tile_17_11_to_tile_18_11_3),
		.in_wire_1_0(vertical_tile_18_11_to_tile_17_11_0),
		.in_wire_1_1(vertical_tile_18_11_to_tile_17_11_1),
		.in_wire_1_2(vertical_tile_18_11_to_tile_17_11_2),
		.in_wire_1_3(vertical_tile_18_11_to_tile_17_11_3),
		.out_wire_2_0(horizontal_tile_17_11_to_tile_17_10_0),
		.out_wire_2_1(horizontal_tile_17_11_to_tile_17_10_1),
		.out_wire_2_2(horizontal_tile_17_11_to_tile_17_10_2),
		.out_wire_2_3(horizontal_tile_17_11_to_tile_17_10_3),
		.in_wire_2_0(horizontal_tile_17_10_to_tile_17_11_0),
		.in_wire_2_1(horizontal_tile_17_10_to_tile_17_11_1),
		.in_wire_2_2(horizontal_tile_17_10_to_tile_17_11_2),
		.in_wire_2_3(horizontal_tile_17_10_to_tile_17_11_3),
		.out_wire_0_0(horizontal_tile_17_11_to_tile_17_12_0),
		.out_wire_0_1(horizontal_tile_17_11_to_tile_17_12_1),
		.out_wire_0_2(horizontal_tile_17_11_to_tile_17_12_2),
		.out_wire_0_3(horizontal_tile_17_11_to_tile_17_12_3),
		.in_wire_0_0(horizontal_tile_17_12_to_tile_17_11_0),
		.in_wire_0_1(horizontal_tile_17_12_to_tile_17_11_1),
		.in_wire_0_2(horizontal_tile_17_12_to_tile_17_11_2),
		.in_wire_0_3(horizontal_tile_17_12_to_tile_17_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(556)
	);

	pe_tile pe_tile_17_12(
		.out_wire_3_0(vertical_tile_17_12_to_tile_16_12_0),
		.out_wire_3_1(vertical_tile_17_12_to_tile_16_12_1),
		.out_wire_3_2(vertical_tile_17_12_to_tile_16_12_2),
		.out_wire_3_3(vertical_tile_17_12_to_tile_16_12_3),
		.in_wire_3_0(vertical_tile_16_12_to_tile_17_12_0),
		.in_wire_3_1(vertical_tile_16_12_to_tile_17_12_1),
		.in_wire_3_2(vertical_tile_16_12_to_tile_17_12_2),
		.in_wire_3_3(vertical_tile_16_12_to_tile_17_12_3),
		.out_wire_1_0(vertical_tile_17_12_to_tile_18_12_0),
		.out_wire_1_1(vertical_tile_17_12_to_tile_18_12_1),
		.out_wire_1_2(vertical_tile_17_12_to_tile_18_12_2),
		.out_wire_1_3(vertical_tile_17_12_to_tile_18_12_3),
		.in_wire_1_0(vertical_tile_18_12_to_tile_17_12_0),
		.in_wire_1_1(vertical_tile_18_12_to_tile_17_12_1),
		.in_wire_1_2(vertical_tile_18_12_to_tile_17_12_2),
		.in_wire_1_3(vertical_tile_18_12_to_tile_17_12_3),
		.out_wire_2_0(horizontal_tile_17_12_to_tile_17_11_0),
		.out_wire_2_1(horizontal_tile_17_12_to_tile_17_11_1),
		.out_wire_2_2(horizontal_tile_17_12_to_tile_17_11_2),
		.out_wire_2_3(horizontal_tile_17_12_to_tile_17_11_3),
		.in_wire_2_0(horizontal_tile_17_11_to_tile_17_12_0),
		.in_wire_2_1(horizontal_tile_17_11_to_tile_17_12_1),
		.in_wire_2_2(horizontal_tile_17_11_to_tile_17_12_2),
		.in_wire_2_3(horizontal_tile_17_11_to_tile_17_12_3),
		.out_wire_0_0(horizontal_tile_17_12_to_tile_17_13_0),
		.out_wire_0_1(horizontal_tile_17_12_to_tile_17_13_1),
		.out_wire_0_2(horizontal_tile_17_12_to_tile_17_13_2),
		.out_wire_0_3(horizontal_tile_17_12_to_tile_17_13_3),
		.in_wire_0_0(horizontal_tile_17_13_to_tile_17_12_0),
		.in_wire_0_1(horizontal_tile_17_13_to_tile_17_12_1),
		.in_wire_0_2(horizontal_tile_17_13_to_tile_17_12_2),
		.in_wire_0_3(horizontal_tile_17_13_to_tile_17_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(557)
	);

	pe_tile pe_tile_17_13(
		.out_wire_3_0(vertical_tile_17_13_to_tile_16_13_0),
		.out_wire_3_1(vertical_tile_17_13_to_tile_16_13_1),
		.out_wire_3_2(vertical_tile_17_13_to_tile_16_13_2),
		.out_wire_3_3(vertical_tile_17_13_to_tile_16_13_3),
		.in_wire_3_0(vertical_tile_16_13_to_tile_17_13_0),
		.in_wire_3_1(vertical_tile_16_13_to_tile_17_13_1),
		.in_wire_3_2(vertical_tile_16_13_to_tile_17_13_2),
		.in_wire_3_3(vertical_tile_16_13_to_tile_17_13_3),
		.out_wire_1_0(vertical_tile_17_13_to_tile_18_13_0),
		.out_wire_1_1(vertical_tile_17_13_to_tile_18_13_1),
		.out_wire_1_2(vertical_tile_17_13_to_tile_18_13_2),
		.out_wire_1_3(vertical_tile_17_13_to_tile_18_13_3),
		.in_wire_1_0(vertical_tile_18_13_to_tile_17_13_0),
		.in_wire_1_1(vertical_tile_18_13_to_tile_17_13_1),
		.in_wire_1_2(vertical_tile_18_13_to_tile_17_13_2),
		.in_wire_1_3(vertical_tile_18_13_to_tile_17_13_3),
		.out_wire_2_0(horizontal_tile_17_13_to_tile_17_12_0),
		.out_wire_2_1(horizontal_tile_17_13_to_tile_17_12_1),
		.out_wire_2_2(horizontal_tile_17_13_to_tile_17_12_2),
		.out_wire_2_3(horizontal_tile_17_13_to_tile_17_12_3),
		.in_wire_2_0(horizontal_tile_17_12_to_tile_17_13_0),
		.in_wire_2_1(horizontal_tile_17_12_to_tile_17_13_1),
		.in_wire_2_2(horizontal_tile_17_12_to_tile_17_13_2),
		.in_wire_2_3(horizontal_tile_17_12_to_tile_17_13_3),
		.out_wire_0_0(horizontal_tile_17_13_to_tile_17_14_0),
		.out_wire_0_1(horizontal_tile_17_13_to_tile_17_14_1),
		.out_wire_0_2(horizontal_tile_17_13_to_tile_17_14_2),
		.out_wire_0_3(horizontal_tile_17_13_to_tile_17_14_3),
		.in_wire_0_0(horizontal_tile_17_14_to_tile_17_13_0),
		.in_wire_0_1(horizontal_tile_17_14_to_tile_17_13_1),
		.in_wire_0_2(horizontal_tile_17_14_to_tile_17_13_2),
		.in_wire_0_3(horizontal_tile_17_14_to_tile_17_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(558)
	);

	pe_tile pe_tile_17_14(
		.out_wire_3_0(vertical_tile_17_14_to_tile_16_14_0),
		.out_wire_3_1(vertical_tile_17_14_to_tile_16_14_1),
		.out_wire_3_2(vertical_tile_17_14_to_tile_16_14_2),
		.out_wire_3_3(vertical_tile_17_14_to_tile_16_14_3),
		.in_wire_3_0(vertical_tile_16_14_to_tile_17_14_0),
		.in_wire_3_1(vertical_tile_16_14_to_tile_17_14_1),
		.in_wire_3_2(vertical_tile_16_14_to_tile_17_14_2),
		.in_wire_3_3(vertical_tile_16_14_to_tile_17_14_3),
		.out_wire_1_0(vertical_tile_17_14_to_tile_18_14_0),
		.out_wire_1_1(vertical_tile_17_14_to_tile_18_14_1),
		.out_wire_1_2(vertical_tile_17_14_to_tile_18_14_2),
		.out_wire_1_3(vertical_tile_17_14_to_tile_18_14_3),
		.in_wire_1_0(vertical_tile_18_14_to_tile_17_14_0),
		.in_wire_1_1(vertical_tile_18_14_to_tile_17_14_1),
		.in_wire_1_2(vertical_tile_18_14_to_tile_17_14_2),
		.in_wire_1_3(vertical_tile_18_14_to_tile_17_14_3),
		.out_wire_2_0(horizontal_tile_17_14_to_tile_17_13_0),
		.out_wire_2_1(horizontal_tile_17_14_to_tile_17_13_1),
		.out_wire_2_2(horizontal_tile_17_14_to_tile_17_13_2),
		.out_wire_2_3(horizontal_tile_17_14_to_tile_17_13_3),
		.in_wire_2_0(horizontal_tile_17_13_to_tile_17_14_0),
		.in_wire_2_1(horizontal_tile_17_13_to_tile_17_14_1),
		.in_wire_2_2(horizontal_tile_17_13_to_tile_17_14_2),
		.in_wire_2_3(horizontal_tile_17_13_to_tile_17_14_3),
		.out_wire_0_0(horizontal_tile_17_14_to_tile_17_15_0),
		.out_wire_0_1(horizontal_tile_17_14_to_tile_17_15_1),
		.out_wire_0_2(horizontal_tile_17_14_to_tile_17_15_2),
		.out_wire_0_3(horizontal_tile_17_14_to_tile_17_15_3),
		.in_wire_0_0(horizontal_tile_17_15_to_tile_17_14_0),
		.in_wire_0_1(horizontal_tile_17_15_to_tile_17_14_1),
		.in_wire_0_2(horizontal_tile_17_15_to_tile_17_14_2),
		.in_wire_0_3(horizontal_tile_17_15_to_tile_17_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(559)
	);

	pe_tile pe_tile_17_15(
		.out_wire_3_0(vertical_tile_17_15_to_tile_16_15_0),
		.out_wire_3_1(vertical_tile_17_15_to_tile_16_15_1),
		.out_wire_3_2(vertical_tile_17_15_to_tile_16_15_2),
		.out_wire_3_3(vertical_tile_17_15_to_tile_16_15_3),
		.in_wire_3_0(vertical_tile_16_15_to_tile_17_15_0),
		.in_wire_3_1(vertical_tile_16_15_to_tile_17_15_1),
		.in_wire_3_2(vertical_tile_16_15_to_tile_17_15_2),
		.in_wire_3_3(vertical_tile_16_15_to_tile_17_15_3),
		.out_wire_1_0(vertical_tile_17_15_to_tile_18_15_0),
		.out_wire_1_1(vertical_tile_17_15_to_tile_18_15_1),
		.out_wire_1_2(vertical_tile_17_15_to_tile_18_15_2),
		.out_wire_1_3(vertical_tile_17_15_to_tile_18_15_3),
		.in_wire_1_0(vertical_tile_18_15_to_tile_17_15_0),
		.in_wire_1_1(vertical_tile_18_15_to_tile_17_15_1),
		.in_wire_1_2(vertical_tile_18_15_to_tile_17_15_2),
		.in_wire_1_3(vertical_tile_18_15_to_tile_17_15_3),
		.out_wire_2_0(horizontal_tile_17_15_to_tile_17_14_0),
		.out_wire_2_1(horizontal_tile_17_15_to_tile_17_14_1),
		.out_wire_2_2(horizontal_tile_17_15_to_tile_17_14_2),
		.out_wire_2_3(horizontal_tile_17_15_to_tile_17_14_3),
		.in_wire_2_0(horizontal_tile_17_14_to_tile_17_15_0),
		.in_wire_2_1(horizontal_tile_17_14_to_tile_17_15_1),
		.in_wire_2_2(horizontal_tile_17_14_to_tile_17_15_2),
		.in_wire_2_3(horizontal_tile_17_14_to_tile_17_15_3),
		.out_wire_0_0(horizontal_tile_17_15_to_tile_17_16_0),
		.out_wire_0_1(horizontal_tile_17_15_to_tile_17_16_1),
		.out_wire_0_2(horizontal_tile_17_15_to_tile_17_16_2),
		.out_wire_0_3(horizontal_tile_17_15_to_tile_17_16_3),
		.in_wire_0_0(horizontal_tile_17_16_to_tile_17_15_0),
		.in_wire_0_1(horizontal_tile_17_16_to_tile_17_15_1),
		.in_wire_0_2(horizontal_tile_17_16_to_tile_17_15_2),
		.in_wire_0_3(horizontal_tile_17_16_to_tile_17_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(560)
	);

	pe_tile pe_tile_17_16(
		.out_wire_3_0(vertical_tile_17_16_to_tile_16_16_0),
		.out_wire_3_1(vertical_tile_17_16_to_tile_16_16_1),
		.out_wire_3_2(vertical_tile_17_16_to_tile_16_16_2),
		.out_wire_3_3(vertical_tile_17_16_to_tile_16_16_3),
		.in_wire_3_0(vertical_tile_16_16_to_tile_17_16_0),
		.in_wire_3_1(vertical_tile_16_16_to_tile_17_16_1),
		.in_wire_3_2(vertical_tile_16_16_to_tile_17_16_2),
		.in_wire_3_3(vertical_tile_16_16_to_tile_17_16_3),
		.out_wire_1_0(vertical_tile_17_16_to_tile_18_16_0),
		.out_wire_1_1(vertical_tile_17_16_to_tile_18_16_1),
		.out_wire_1_2(vertical_tile_17_16_to_tile_18_16_2),
		.out_wire_1_3(vertical_tile_17_16_to_tile_18_16_3),
		.in_wire_1_0(vertical_tile_18_16_to_tile_17_16_0),
		.in_wire_1_1(vertical_tile_18_16_to_tile_17_16_1),
		.in_wire_1_2(vertical_tile_18_16_to_tile_17_16_2),
		.in_wire_1_3(vertical_tile_18_16_to_tile_17_16_3),
		.out_wire_2_0(horizontal_tile_17_16_to_tile_17_15_0),
		.out_wire_2_1(horizontal_tile_17_16_to_tile_17_15_1),
		.out_wire_2_2(horizontal_tile_17_16_to_tile_17_15_2),
		.out_wire_2_3(horizontal_tile_17_16_to_tile_17_15_3),
		.in_wire_2_0(horizontal_tile_17_15_to_tile_17_16_0),
		.in_wire_2_1(horizontal_tile_17_15_to_tile_17_16_1),
		.in_wire_2_2(horizontal_tile_17_15_to_tile_17_16_2),
		.in_wire_2_3(horizontal_tile_17_15_to_tile_17_16_3),
		.out_wire_0_0(horizontal_tile_17_16_to_tile_17_17_0),
		.out_wire_0_1(horizontal_tile_17_16_to_tile_17_17_1),
		.out_wire_0_2(horizontal_tile_17_16_to_tile_17_17_2),
		.out_wire_0_3(horizontal_tile_17_16_to_tile_17_17_3),
		.in_wire_0_0(horizontal_tile_17_17_to_tile_17_16_0),
		.in_wire_0_1(horizontal_tile_17_17_to_tile_17_16_1),
		.in_wire_0_2(horizontal_tile_17_17_to_tile_17_16_2),
		.in_wire_0_3(horizontal_tile_17_17_to_tile_17_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(561)
	);

	pe_tile pe_tile_17_17(
		.out_wire_3_0(vertical_tile_17_17_to_tile_16_17_0),
		.out_wire_3_1(vertical_tile_17_17_to_tile_16_17_1),
		.out_wire_3_2(vertical_tile_17_17_to_tile_16_17_2),
		.out_wire_3_3(vertical_tile_17_17_to_tile_16_17_3),
		.in_wire_3_0(vertical_tile_16_17_to_tile_17_17_0),
		.in_wire_3_1(vertical_tile_16_17_to_tile_17_17_1),
		.in_wire_3_2(vertical_tile_16_17_to_tile_17_17_2),
		.in_wire_3_3(vertical_tile_16_17_to_tile_17_17_3),
		.out_wire_1_0(vertical_tile_17_17_to_tile_18_17_0),
		.out_wire_1_1(vertical_tile_17_17_to_tile_18_17_1),
		.out_wire_1_2(vertical_tile_17_17_to_tile_18_17_2),
		.out_wire_1_3(vertical_tile_17_17_to_tile_18_17_3),
		.in_wire_1_0(vertical_tile_18_17_to_tile_17_17_0),
		.in_wire_1_1(vertical_tile_18_17_to_tile_17_17_1),
		.in_wire_1_2(vertical_tile_18_17_to_tile_17_17_2),
		.in_wire_1_3(vertical_tile_18_17_to_tile_17_17_3),
		.out_wire_2_0(horizontal_tile_17_17_to_tile_17_16_0),
		.out_wire_2_1(horizontal_tile_17_17_to_tile_17_16_1),
		.out_wire_2_2(horizontal_tile_17_17_to_tile_17_16_2),
		.out_wire_2_3(horizontal_tile_17_17_to_tile_17_16_3),
		.in_wire_2_0(horizontal_tile_17_16_to_tile_17_17_0),
		.in_wire_2_1(horizontal_tile_17_16_to_tile_17_17_1),
		.in_wire_2_2(horizontal_tile_17_16_to_tile_17_17_2),
		.in_wire_2_3(horizontal_tile_17_16_to_tile_17_17_3),
		.out_wire_0_0(horizontal_tile_17_17_to_tile_17_18_0),
		.out_wire_0_1(horizontal_tile_17_17_to_tile_17_18_1),
		.out_wire_0_2(horizontal_tile_17_17_to_tile_17_18_2),
		.out_wire_0_3(horizontal_tile_17_17_to_tile_17_18_3),
		.in_wire_0_0(horizontal_tile_17_18_to_tile_17_17_0),
		.in_wire_0_1(horizontal_tile_17_18_to_tile_17_17_1),
		.in_wire_0_2(horizontal_tile_17_18_to_tile_17_17_2),
		.in_wire_0_3(horizontal_tile_17_18_to_tile_17_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(562)
	);

	pe_tile pe_tile_17_18(
		.out_wire_3_0(vertical_tile_17_18_to_tile_16_18_0),
		.out_wire_3_1(vertical_tile_17_18_to_tile_16_18_1),
		.out_wire_3_2(vertical_tile_17_18_to_tile_16_18_2),
		.out_wire_3_3(vertical_tile_17_18_to_tile_16_18_3),
		.in_wire_3_0(vertical_tile_16_18_to_tile_17_18_0),
		.in_wire_3_1(vertical_tile_16_18_to_tile_17_18_1),
		.in_wire_3_2(vertical_tile_16_18_to_tile_17_18_2),
		.in_wire_3_3(vertical_tile_16_18_to_tile_17_18_3),
		.out_wire_1_0(vertical_tile_17_18_to_tile_18_18_0),
		.out_wire_1_1(vertical_tile_17_18_to_tile_18_18_1),
		.out_wire_1_2(vertical_tile_17_18_to_tile_18_18_2),
		.out_wire_1_3(vertical_tile_17_18_to_tile_18_18_3),
		.in_wire_1_0(vertical_tile_18_18_to_tile_17_18_0),
		.in_wire_1_1(vertical_tile_18_18_to_tile_17_18_1),
		.in_wire_1_2(vertical_tile_18_18_to_tile_17_18_2),
		.in_wire_1_3(vertical_tile_18_18_to_tile_17_18_3),
		.out_wire_2_0(horizontal_tile_17_18_to_tile_17_17_0),
		.out_wire_2_1(horizontal_tile_17_18_to_tile_17_17_1),
		.out_wire_2_2(horizontal_tile_17_18_to_tile_17_17_2),
		.out_wire_2_3(horizontal_tile_17_18_to_tile_17_17_3),
		.in_wire_2_0(horizontal_tile_17_17_to_tile_17_18_0),
		.in_wire_2_1(horizontal_tile_17_17_to_tile_17_18_1),
		.in_wire_2_2(horizontal_tile_17_17_to_tile_17_18_2),
		.in_wire_2_3(horizontal_tile_17_17_to_tile_17_18_3),
		.out_wire_0_0(horizontal_tile_17_18_to_tile_17_19_0),
		.out_wire_0_1(horizontal_tile_17_18_to_tile_17_19_1),
		.out_wire_0_2(horizontal_tile_17_18_to_tile_17_19_2),
		.out_wire_0_3(horizontal_tile_17_18_to_tile_17_19_3),
		.in_wire_0_0(horizontal_tile_17_19_to_tile_17_18_0),
		.in_wire_0_1(horizontal_tile_17_19_to_tile_17_18_1),
		.in_wire_0_2(horizontal_tile_17_19_to_tile_17_18_2),
		.in_wire_0_3(horizontal_tile_17_19_to_tile_17_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(563)
	);

	pe_tile pe_tile_17_19(
		.out_wire_3_0(vertical_tile_17_19_to_tile_16_19_0),
		.out_wire_3_1(vertical_tile_17_19_to_tile_16_19_1),
		.out_wire_3_2(vertical_tile_17_19_to_tile_16_19_2),
		.out_wire_3_3(vertical_tile_17_19_to_tile_16_19_3),
		.in_wire_3_0(vertical_tile_16_19_to_tile_17_19_0),
		.in_wire_3_1(vertical_tile_16_19_to_tile_17_19_1),
		.in_wire_3_2(vertical_tile_16_19_to_tile_17_19_2),
		.in_wire_3_3(vertical_tile_16_19_to_tile_17_19_3),
		.out_wire_1_0(vertical_tile_17_19_to_tile_18_19_0),
		.out_wire_1_1(vertical_tile_17_19_to_tile_18_19_1),
		.out_wire_1_2(vertical_tile_17_19_to_tile_18_19_2),
		.out_wire_1_3(vertical_tile_17_19_to_tile_18_19_3),
		.in_wire_1_0(vertical_tile_18_19_to_tile_17_19_0),
		.in_wire_1_1(vertical_tile_18_19_to_tile_17_19_1),
		.in_wire_1_2(vertical_tile_18_19_to_tile_17_19_2),
		.in_wire_1_3(vertical_tile_18_19_to_tile_17_19_3),
		.out_wire_2_0(horizontal_tile_17_19_to_tile_17_18_0),
		.out_wire_2_1(horizontal_tile_17_19_to_tile_17_18_1),
		.out_wire_2_2(horizontal_tile_17_19_to_tile_17_18_2),
		.out_wire_2_3(horizontal_tile_17_19_to_tile_17_18_3),
		.in_wire_2_0(horizontal_tile_17_18_to_tile_17_19_0),
		.in_wire_2_1(horizontal_tile_17_18_to_tile_17_19_1),
		.in_wire_2_2(horizontal_tile_17_18_to_tile_17_19_2),
		.in_wire_2_3(horizontal_tile_17_18_to_tile_17_19_3),
		.out_wire_0_0(horizontal_tile_17_19_to_tile_17_20_0),
		.out_wire_0_1(horizontal_tile_17_19_to_tile_17_20_1),
		.out_wire_0_2(horizontal_tile_17_19_to_tile_17_20_2),
		.out_wire_0_3(horizontal_tile_17_19_to_tile_17_20_3),
		.in_wire_0_0(horizontal_tile_17_20_to_tile_17_19_0),
		.in_wire_0_1(horizontal_tile_17_20_to_tile_17_19_1),
		.in_wire_0_2(horizontal_tile_17_20_to_tile_17_19_2),
		.in_wire_0_3(horizontal_tile_17_20_to_tile_17_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(564)
	);

	pe_tile pe_tile_17_20(
		.out_wire_3_0(vertical_tile_17_20_to_tile_16_20_0),
		.out_wire_3_1(vertical_tile_17_20_to_tile_16_20_1),
		.out_wire_3_2(vertical_tile_17_20_to_tile_16_20_2),
		.out_wire_3_3(vertical_tile_17_20_to_tile_16_20_3),
		.in_wire_3_0(vertical_tile_16_20_to_tile_17_20_0),
		.in_wire_3_1(vertical_tile_16_20_to_tile_17_20_1),
		.in_wire_3_2(vertical_tile_16_20_to_tile_17_20_2),
		.in_wire_3_3(vertical_tile_16_20_to_tile_17_20_3),
		.out_wire_1_0(vertical_tile_17_20_to_tile_18_20_0),
		.out_wire_1_1(vertical_tile_17_20_to_tile_18_20_1),
		.out_wire_1_2(vertical_tile_17_20_to_tile_18_20_2),
		.out_wire_1_3(vertical_tile_17_20_to_tile_18_20_3),
		.in_wire_1_0(vertical_tile_18_20_to_tile_17_20_0),
		.in_wire_1_1(vertical_tile_18_20_to_tile_17_20_1),
		.in_wire_1_2(vertical_tile_18_20_to_tile_17_20_2),
		.in_wire_1_3(vertical_tile_18_20_to_tile_17_20_3),
		.out_wire_2_0(horizontal_tile_17_20_to_tile_17_19_0),
		.out_wire_2_1(horizontal_tile_17_20_to_tile_17_19_1),
		.out_wire_2_2(horizontal_tile_17_20_to_tile_17_19_2),
		.out_wire_2_3(horizontal_tile_17_20_to_tile_17_19_3),
		.in_wire_2_0(horizontal_tile_17_19_to_tile_17_20_0),
		.in_wire_2_1(horizontal_tile_17_19_to_tile_17_20_1),
		.in_wire_2_2(horizontal_tile_17_19_to_tile_17_20_2),
		.in_wire_2_3(horizontal_tile_17_19_to_tile_17_20_3),
		.out_wire_0_0(horizontal_tile_17_20_to_tile_17_21_0),
		.out_wire_0_1(horizontal_tile_17_20_to_tile_17_21_1),
		.out_wire_0_2(horizontal_tile_17_20_to_tile_17_21_2),
		.out_wire_0_3(horizontal_tile_17_20_to_tile_17_21_3),
		.in_wire_0_0(horizontal_tile_17_21_to_tile_17_20_0),
		.in_wire_0_1(horizontal_tile_17_21_to_tile_17_20_1),
		.in_wire_0_2(horizontal_tile_17_21_to_tile_17_20_2),
		.in_wire_0_3(horizontal_tile_17_21_to_tile_17_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(565)
	);

	pe_tile pe_tile_17_21(
		.out_wire_3_0(vertical_tile_17_21_to_tile_16_21_0),
		.out_wire_3_1(vertical_tile_17_21_to_tile_16_21_1),
		.out_wire_3_2(vertical_tile_17_21_to_tile_16_21_2),
		.out_wire_3_3(vertical_tile_17_21_to_tile_16_21_3),
		.in_wire_3_0(vertical_tile_16_21_to_tile_17_21_0),
		.in_wire_3_1(vertical_tile_16_21_to_tile_17_21_1),
		.in_wire_3_2(vertical_tile_16_21_to_tile_17_21_2),
		.in_wire_3_3(vertical_tile_16_21_to_tile_17_21_3),
		.out_wire_1_0(vertical_tile_17_21_to_tile_18_21_0),
		.out_wire_1_1(vertical_tile_17_21_to_tile_18_21_1),
		.out_wire_1_2(vertical_tile_17_21_to_tile_18_21_2),
		.out_wire_1_3(vertical_tile_17_21_to_tile_18_21_3),
		.in_wire_1_0(vertical_tile_18_21_to_tile_17_21_0),
		.in_wire_1_1(vertical_tile_18_21_to_tile_17_21_1),
		.in_wire_1_2(vertical_tile_18_21_to_tile_17_21_2),
		.in_wire_1_3(vertical_tile_18_21_to_tile_17_21_3),
		.out_wire_2_0(horizontal_tile_17_21_to_tile_17_20_0),
		.out_wire_2_1(horizontal_tile_17_21_to_tile_17_20_1),
		.out_wire_2_2(horizontal_tile_17_21_to_tile_17_20_2),
		.out_wire_2_3(horizontal_tile_17_21_to_tile_17_20_3),
		.in_wire_2_0(horizontal_tile_17_20_to_tile_17_21_0),
		.in_wire_2_1(horizontal_tile_17_20_to_tile_17_21_1),
		.in_wire_2_2(horizontal_tile_17_20_to_tile_17_21_2),
		.in_wire_2_3(horizontal_tile_17_20_to_tile_17_21_3),
		.out_wire_0_0(horizontal_tile_17_21_to_tile_17_22_0),
		.out_wire_0_1(horizontal_tile_17_21_to_tile_17_22_1),
		.out_wire_0_2(horizontal_tile_17_21_to_tile_17_22_2),
		.out_wire_0_3(horizontal_tile_17_21_to_tile_17_22_3),
		.in_wire_0_0(horizontal_tile_17_22_to_tile_17_21_0),
		.in_wire_0_1(horizontal_tile_17_22_to_tile_17_21_1),
		.in_wire_0_2(horizontal_tile_17_22_to_tile_17_21_2),
		.in_wire_0_3(horizontal_tile_17_22_to_tile_17_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(566)
	);

	pe_tile pe_tile_17_22(
		.out_wire_3_0(vertical_tile_17_22_to_tile_16_22_0),
		.out_wire_3_1(vertical_tile_17_22_to_tile_16_22_1),
		.out_wire_3_2(vertical_tile_17_22_to_tile_16_22_2),
		.out_wire_3_3(vertical_tile_17_22_to_tile_16_22_3),
		.in_wire_3_0(vertical_tile_16_22_to_tile_17_22_0),
		.in_wire_3_1(vertical_tile_16_22_to_tile_17_22_1),
		.in_wire_3_2(vertical_tile_16_22_to_tile_17_22_2),
		.in_wire_3_3(vertical_tile_16_22_to_tile_17_22_3),
		.out_wire_1_0(vertical_tile_17_22_to_tile_18_22_0),
		.out_wire_1_1(vertical_tile_17_22_to_tile_18_22_1),
		.out_wire_1_2(vertical_tile_17_22_to_tile_18_22_2),
		.out_wire_1_3(vertical_tile_17_22_to_tile_18_22_3),
		.in_wire_1_0(vertical_tile_18_22_to_tile_17_22_0),
		.in_wire_1_1(vertical_tile_18_22_to_tile_17_22_1),
		.in_wire_1_2(vertical_tile_18_22_to_tile_17_22_2),
		.in_wire_1_3(vertical_tile_18_22_to_tile_17_22_3),
		.out_wire_2_0(horizontal_tile_17_22_to_tile_17_21_0),
		.out_wire_2_1(horizontal_tile_17_22_to_tile_17_21_1),
		.out_wire_2_2(horizontal_tile_17_22_to_tile_17_21_2),
		.out_wire_2_3(horizontal_tile_17_22_to_tile_17_21_3),
		.in_wire_2_0(horizontal_tile_17_21_to_tile_17_22_0),
		.in_wire_2_1(horizontal_tile_17_21_to_tile_17_22_1),
		.in_wire_2_2(horizontal_tile_17_21_to_tile_17_22_2),
		.in_wire_2_3(horizontal_tile_17_21_to_tile_17_22_3),
		.out_wire_0_0(horizontal_tile_17_22_to_tile_17_23_0),
		.out_wire_0_1(horizontal_tile_17_22_to_tile_17_23_1),
		.out_wire_0_2(horizontal_tile_17_22_to_tile_17_23_2),
		.out_wire_0_3(horizontal_tile_17_22_to_tile_17_23_3),
		.in_wire_0_0(horizontal_tile_17_23_to_tile_17_22_0),
		.in_wire_0_1(horizontal_tile_17_23_to_tile_17_22_1),
		.in_wire_0_2(horizontal_tile_17_23_to_tile_17_22_2),
		.in_wire_0_3(horizontal_tile_17_23_to_tile_17_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(567)
	);

	pe_tile pe_tile_17_23(
		.out_wire_3_0(vertical_tile_17_23_to_tile_16_23_0),
		.out_wire_3_1(vertical_tile_17_23_to_tile_16_23_1),
		.out_wire_3_2(vertical_tile_17_23_to_tile_16_23_2),
		.out_wire_3_3(vertical_tile_17_23_to_tile_16_23_3),
		.in_wire_3_0(vertical_tile_16_23_to_tile_17_23_0),
		.in_wire_3_1(vertical_tile_16_23_to_tile_17_23_1),
		.in_wire_3_2(vertical_tile_16_23_to_tile_17_23_2),
		.in_wire_3_3(vertical_tile_16_23_to_tile_17_23_3),
		.out_wire_1_0(vertical_tile_17_23_to_tile_18_23_0),
		.out_wire_1_1(vertical_tile_17_23_to_tile_18_23_1),
		.out_wire_1_2(vertical_tile_17_23_to_tile_18_23_2),
		.out_wire_1_3(vertical_tile_17_23_to_tile_18_23_3),
		.in_wire_1_0(vertical_tile_18_23_to_tile_17_23_0),
		.in_wire_1_1(vertical_tile_18_23_to_tile_17_23_1),
		.in_wire_1_2(vertical_tile_18_23_to_tile_17_23_2),
		.in_wire_1_3(vertical_tile_18_23_to_tile_17_23_3),
		.out_wire_2_0(horizontal_tile_17_23_to_tile_17_22_0),
		.out_wire_2_1(horizontal_tile_17_23_to_tile_17_22_1),
		.out_wire_2_2(horizontal_tile_17_23_to_tile_17_22_2),
		.out_wire_2_3(horizontal_tile_17_23_to_tile_17_22_3),
		.in_wire_2_0(horizontal_tile_17_22_to_tile_17_23_0),
		.in_wire_2_1(horizontal_tile_17_22_to_tile_17_23_1),
		.in_wire_2_2(horizontal_tile_17_22_to_tile_17_23_2),
		.in_wire_2_3(horizontal_tile_17_22_to_tile_17_23_3),
		.out_wire_0_0(horizontal_tile_17_23_to_tile_17_24_0),
		.out_wire_0_1(horizontal_tile_17_23_to_tile_17_24_1),
		.out_wire_0_2(horizontal_tile_17_23_to_tile_17_24_2),
		.out_wire_0_3(horizontal_tile_17_23_to_tile_17_24_3),
		.in_wire_0_0(horizontal_tile_17_24_to_tile_17_23_0),
		.in_wire_0_1(horizontal_tile_17_24_to_tile_17_23_1),
		.in_wire_0_2(horizontal_tile_17_24_to_tile_17_23_2),
		.in_wire_0_3(horizontal_tile_17_24_to_tile_17_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(568)
	);

	pe_tile pe_tile_17_24(
		.out_wire_3_0(vertical_tile_17_24_to_tile_16_24_0),
		.out_wire_3_1(vertical_tile_17_24_to_tile_16_24_1),
		.out_wire_3_2(vertical_tile_17_24_to_tile_16_24_2),
		.out_wire_3_3(vertical_tile_17_24_to_tile_16_24_3),
		.in_wire_3_0(vertical_tile_16_24_to_tile_17_24_0),
		.in_wire_3_1(vertical_tile_16_24_to_tile_17_24_1),
		.in_wire_3_2(vertical_tile_16_24_to_tile_17_24_2),
		.in_wire_3_3(vertical_tile_16_24_to_tile_17_24_3),
		.out_wire_1_0(vertical_tile_17_24_to_tile_18_24_0),
		.out_wire_1_1(vertical_tile_17_24_to_tile_18_24_1),
		.out_wire_1_2(vertical_tile_17_24_to_tile_18_24_2),
		.out_wire_1_3(vertical_tile_17_24_to_tile_18_24_3),
		.in_wire_1_0(vertical_tile_18_24_to_tile_17_24_0),
		.in_wire_1_1(vertical_tile_18_24_to_tile_17_24_1),
		.in_wire_1_2(vertical_tile_18_24_to_tile_17_24_2),
		.in_wire_1_3(vertical_tile_18_24_to_tile_17_24_3),
		.out_wire_2_0(horizontal_tile_17_24_to_tile_17_23_0),
		.out_wire_2_1(horizontal_tile_17_24_to_tile_17_23_1),
		.out_wire_2_2(horizontal_tile_17_24_to_tile_17_23_2),
		.out_wire_2_3(horizontal_tile_17_24_to_tile_17_23_3),
		.in_wire_2_0(horizontal_tile_17_23_to_tile_17_24_0),
		.in_wire_2_1(horizontal_tile_17_23_to_tile_17_24_1),
		.in_wire_2_2(horizontal_tile_17_23_to_tile_17_24_2),
		.in_wire_2_3(horizontal_tile_17_23_to_tile_17_24_3),
		.out_wire_0_0(horizontal_tile_17_24_to_tile_17_25_0),
		.out_wire_0_1(horizontal_tile_17_24_to_tile_17_25_1),
		.out_wire_0_2(horizontal_tile_17_24_to_tile_17_25_2),
		.out_wire_0_3(horizontal_tile_17_24_to_tile_17_25_3),
		.in_wire_0_0(horizontal_tile_17_25_to_tile_17_24_0),
		.in_wire_0_1(horizontal_tile_17_25_to_tile_17_24_1),
		.in_wire_0_2(horizontal_tile_17_25_to_tile_17_24_2),
		.in_wire_0_3(horizontal_tile_17_25_to_tile_17_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(569)
	);

	pe_tile pe_tile_17_25(
		.out_wire_3_0(vertical_tile_17_25_to_tile_16_25_0),
		.out_wire_3_1(vertical_tile_17_25_to_tile_16_25_1),
		.out_wire_3_2(vertical_tile_17_25_to_tile_16_25_2),
		.out_wire_3_3(vertical_tile_17_25_to_tile_16_25_3),
		.in_wire_3_0(vertical_tile_16_25_to_tile_17_25_0),
		.in_wire_3_1(vertical_tile_16_25_to_tile_17_25_1),
		.in_wire_3_2(vertical_tile_16_25_to_tile_17_25_2),
		.in_wire_3_3(vertical_tile_16_25_to_tile_17_25_3),
		.out_wire_1_0(vertical_tile_17_25_to_tile_18_25_0),
		.out_wire_1_1(vertical_tile_17_25_to_tile_18_25_1),
		.out_wire_1_2(vertical_tile_17_25_to_tile_18_25_2),
		.out_wire_1_3(vertical_tile_17_25_to_tile_18_25_3),
		.in_wire_1_0(vertical_tile_18_25_to_tile_17_25_0),
		.in_wire_1_1(vertical_tile_18_25_to_tile_17_25_1),
		.in_wire_1_2(vertical_tile_18_25_to_tile_17_25_2),
		.in_wire_1_3(vertical_tile_18_25_to_tile_17_25_3),
		.out_wire_2_0(horizontal_tile_17_25_to_tile_17_24_0),
		.out_wire_2_1(horizontal_tile_17_25_to_tile_17_24_1),
		.out_wire_2_2(horizontal_tile_17_25_to_tile_17_24_2),
		.out_wire_2_3(horizontal_tile_17_25_to_tile_17_24_3),
		.in_wire_2_0(horizontal_tile_17_24_to_tile_17_25_0),
		.in_wire_2_1(horizontal_tile_17_24_to_tile_17_25_1),
		.in_wire_2_2(horizontal_tile_17_24_to_tile_17_25_2),
		.in_wire_2_3(horizontal_tile_17_24_to_tile_17_25_3),
		.out_wire_0_0(horizontal_tile_17_25_to_tile_17_26_0),
		.out_wire_0_1(horizontal_tile_17_25_to_tile_17_26_1),
		.out_wire_0_2(horizontal_tile_17_25_to_tile_17_26_2),
		.out_wire_0_3(horizontal_tile_17_25_to_tile_17_26_3),
		.in_wire_0_0(horizontal_tile_17_26_to_tile_17_25_0),
		.in_wire_0_1(horizontal_tile_17_26_to_tile_17_25_1),
		.in_wire_0_2(horizontal_tile_17_26_to_tile_17_25_2),
		.in_wire_0_3(horizontal_tile_17_26_to_tile_17_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(570)
	);

	pe_tile pe_tile_17_26(
		.out_wire_3_0(vertical_tile_17_26_to_tile_16_26_0),
		.out_wire_3_1(vertical_tile_17_26_to_tile_16_26_1),
		.out_wire_3_2(vertical_tile_17_26_to_tile_16_26_2),
		.out_wire_3_3(vertical_tile_17_26_to_tile_16_26_3),
		.in_wire_3_0(vertical_tile_16_26_to_tile_17_26_0),
		.in_wire_3_1(vertical_tile_16_26_to_tile_17_26_1),
		.in_wire_3_2(vertical_tile_16_26_to_tile_17_26_2),
		.in_wire_3_3(vertical_tile_16_26_to_tile_17_26_3),
		.out_wire_1_0(vertical_tile_17_26_to_tile_18_26_0),
		.out_wire_1_1(vertical_tile_17_26_to_tile_18_26_1),
		.out_wire_1_2(vertical_tile_17_26_to_tile_18_26_2),
		.out_wire_1_3(vertical_tile_17_26_to_tile_18_26_3),
		.in_wire_1_0(vertical_tile_18_26_to_tile_17_26_0),
		.in_wire_1_1(vertical_tile_18_26_to_tile_17_26_1),
		.in_wire_1_2(vertical_tile_18_26_to_tile_17_26_2),
		.in_wire_1_3(vertical_tile_18_26_to_tile_17_26_3),
		.out_wire_2_0(horizontal_tile_17_26_to_tile_17_25_0),
		.out_wire_2_1(horizontal_tile_17_26_to_tile_17_25_1),
		.out_wire_2_2(horizontal_tile_17_26_to_tile_17_25_2),
		.out_wire_2_3(horizontal_tile_17_26_to_tile_17_25_3),
		.in_wire_2_0(horizontal_tile_17_25_to_tile_17_26_0),
		.in_wire_2_1(horizontal_tile_17_25_to_tile_17_26_1),
		.in_wire_2_2(horizontal_tile_17_25_to_tile_17_26_2),
		.in_wire_2_3(horizontal_tile_17_25_to_tile_17_26_3),
		.out_wire_0_0(horizontal_tile_17_26_to_tile_17_27_0),
		.out_wire_0_1(horizontal_tile_17_26_to_tile_17_27_1),
		.out_wire_0_2(horizontal_tile_17_26_to_tile_17_27_2),
		.out_wire_0_3(horizontal_tile_17_26_to_tile_17_27_3),
		.in_wire_0_0(horizontal_tile_17_27_to_tile_17_26_0),
		.in_wire_0_1(horizontal_tile_17_27_to_tile_17_26_1),
		.in_wire_0_2(horizontal_tile_17_27_to_tile_17_26_2),
		.in_wire_0_3(horizontal_tile_17_27_to_tile_17_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(571)
	);

	pe_tile pe_tile_17_27(
		.out_wire_3_0(vertical_tile_17_27_to_tile_16_27_0),
		.out_wire_3_1(vertical_tile_17_27_to_tile_16_27_1),
		.out_wire_3_2(vertical_tile_17_27_to_tile_16_27_2),
		.out_wire_3_3(vertical_tile_17_27_to_tile_16_27_3),
		.in_wire_3_0(vertical_tile_16_27_to_tile_17_27_0),
		.in_wire_3_1(vertical_tile_16_27_to_tile_17_27_1),
		.in_wire_3_2(vertical_tile_16_27_to_tile_17_27_2),
		.in_wire_3_3(vertical_tile_16_27_to_tile_17_27_3),
		.out_wire_1_0(vertical_tile_17_27_to_tile_18_27_0),
		.out_wire_1_1(vertical_tile_17_27_to_tile_18_27_1),
		.out_wire_1_2(vertical_tile_17_27_to_tile_18_27_2),
		.out_wire_1_3(vertical_tile_17_27_to_tile_18_27_3),
		.in_wire_1_0(vertical_tile_18_27_to_tile_17_27_0),
		.in_wire_1_1(vertical_tile_18_27_to_tile_17_27_1),
		.in_wire_1_2(vertical_tile_18_27_to_tile_17_27_2),
		.in_wire_1_3(vertical_tile_18_27_to_tile_17_27_3),
		.out_wire_2_0(horizontal_tile_17_27_to_tile_17_26_0),
		.out_wire_2_1(horizontal_tile_17_27_to_tile_17_26_1),
		.out_wire_2_2(horizontal_tile_17_27_to_tile_17_26_2),
		.out_wire_2_3(horizontal_tile_17_27_to_tile_17_26_3),
		.in_wire_2_0(horizontal_tile_17_26_to_tile_17_27_0),
		.in_wire_2_1(horizontal_tile_17_26_to_tile_17_27_1),
		.in_wire_2_2(horizontal_tile_17_26_to_tile_17_27_2),
		.in_wire_2_3(horizontal_tile_17_26_to_tile_17_27_3),
		.out_wire_0_0(horizontal_tile_17_27_to_tile_17_28_0),
		.out_wire_0_1(horizontal_tile_17_27_to_tile_17_28_1),
		.out_wire_0_2(horizontal_tile_17_27_to_tile_17_28_2),
		.out_wire_0_3(horizontal_tile_17_27_to_tile_17_28_3),
		.in_wire_0_0(horizontal_tile_17_28_to_tile_17_27_0),
		.in_wire_0_1(horizontal_tile_17_28_to_tile_17_27_1),
		.in_wire_0_2(horizontal_tile_17_28_to_tile_17_27_2),
		.in_wire_0_3(horizontal_tile_17_28_to_tile_17_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(572)
	);

	pe_tile pe_tile_17_28(
		.out_wire_3_0(vertical_tile_17_28_to_tile_16_28_0),
		.out_wire_3_1(vertical_tile_17_28_to_tile_16_28_1),
		.out_wire_3_2(vertical_tile_17_28_to_tile_16_28_2),
		.out_wire_3_3(vertical_tile_17_28_to_tile_16_28_3),
		.in_wire_3_0(vertical_tile_16_28_to_tile_17_28_0),
		.in_wire_3_1(vertical_tile_16_28_to_tile_17_28_1),
		.in_wire_3_2(vertical_tile_16_28_to_tile_17_28_2),
		.in_wire_3_3(vertical_tile_16_28_to_tile_17_28_3),
		.out_wire_1_0(vertical_tile_17_28_to_tile_18_28_0),
		.out_wire_1_1(vertical_tile_17_28_to_tile_18_28_1),
		.out_wire_1_2(vertical_tile_17_28_to_tile_18_28_2),
		.out_wire_1_3(vertical_tile_17_28_to_tile_18_28_3),
		.in_wire_1_0(vertical_tile_18_28_to_tile_17_28_0),
		.in_wire_1_1(vertical_tile_18_28_to_tile_17_28_1),
		.in_wire_1_2(vertical_tile_18_28_to_tile_17_28_2),
		.in_wire_1_3(vertical_tile_18_28_to_tile_17_28_3),
		.out_wire_2_0(horizontal_tile_17_28_to_tile_17_27_0),
		.out_wire_2_1(horizontal_tile_17_28_to_tile_17_27_1),
		.out_wire_2_2(horizontal_tile_17_28_to_tile_17_27_2),
		.out_wire_2_3(horizontal_tile_17_28_to_tile_17_27_3),
		.in_wire_2_0(horizontal_tile_17_27_to_tile_17_28_0),
		.in_wire_2_1(horizontal_tile_17_27_to_tile_17_28_1),
		.in_wire_2_2(horizontal_tile_17_27_to_tile_17_28_2),
		.in_wire_2_3(horizontal_tile_17_27_to_tile_17_28_3),
		.out_wire_0_0(horizontal_tile_17_28_to_tile_17_29_0),
		.out_wire_0_1(horizontal_tile_17_28_to_tile_17_29_1),
		.out_wire_0_2(horizontal_tile_17_28_to_tile_17_29_2),
		.out_wire_0_3(horizontal_tile_17_28_to_tile_17_29_3),
		.in_wire_0_0(horizontal_tile_17_29_to_tile_17_28_0),
		.in_wire_0_1(horizontal_tile_17_29_to_tile_17_28_1),
		.in_wire_0_2(horizontal_tile_17_29_to_tile_17_28_2),
		.in_wire_0_3(horizontal_tile_17_29_to_tile_17_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(573)
	);

	pe_tile pe_tile_17_29(
		.out_wire_3_0(vertical_tile_17_29_to_tile_16_29_0),
		.out_wire_3_1(vertical_tile_17_29_to_tile_16_29_1),
		.out_wire_3_2(vertical_tile_17_29_to_tile_16_29_2),
		.out_wire_3_3(vertical_tile_17_29_to_tile_16_29_3),
		.in_wire_3_0(vertical_tile_16_29_to_tile_17_29_0),
		.in_wire_3_1(vertical_tile_16_29_to_tile_17_29_1),
		.in_wire_3_2(vertical_tile_16_29_to_tile_17_29_2),
		.in_wire_3_3(vertical_tile_16_29_to_tile_17_29_3),
		.out_wire_1_0(vertical_tile_17_29_to_tile_18_29_0),
		.out_wire_1_1(vertical_tile_17_29_to_tile_18_29_1),
		.out_wire_1_2(vertical_tile_17_29_to_tile_18_29_2),
		.out_wire_1_3(vertical_tile_17_29_to_tile_18_29_3),
		.in_wire_1_0(vertical_tile_18_29_to_tile_17_29_0),
		.in_wire_1_1(vertical_tile_18_29_to_tile_17_29_1),
		.in_wire_1_2(vertical_tile_18_29_to_tile_17_29_2),
		.in_wire_1_3(vertical_tile_18_29_to_tile_17_29_3),
		.out_wire_2_0(horizontal_tile_17_29_to_tile_17_28_0),
		.out_wire_2_1(horizontal_tile_17_29_to_tile_17_28_1),
		.out_wire_2_2(horizontal_tile_17_29_to_tile_17_28_2),
		.out_wire_2_3(horizontal_tile_17_29_to_tile_17_28_3),
		.in_wire_2_0(horizontal_tile_17_28_to_tile_17_29_0),
		.in_wire_2_1(horizontal_tile_17_28_to_tile_17_29_1),
		.in_wire_2_2(horizontal_tile_17_28_to_tile_17_29_2),
		.in_wire_2_3(horizontal_tile_17_28_to_tile_17_29_3),
		.out_wire_0_0(horizontal_tile_17_29_to_tile_17_30_0),
		.out_wire_0_1(horizontal_tile_17_29_to_tile_17_30_1),
		.out_wire_0_2(horizontal_tile_17_29_to_tile_17_30_2),
		.out_wire_0_3(horizontal_tile_17_29_to_tile_17_30_3),
		.in_wire_0_0(horizontal_tile_17_30_to_tile_17_29_0),
		.in_wire_0_1(horizontal_tile_17_30_to_tile_17_29_1),
		.in_wire_0_2(horizontal_tile_17_30_to_tile_17_29_2),
		.in_wire_0_3(horizontal_tile_17_30_to_tile_17_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(574)
	);

	pe_tile pe_tile_17_30(
		.out_wire_3_0(vertical_tile_17_30_to_tile_16_30_0),
		.out_wire_3_1(vertical_tile_17_30_to_tile_16_30_1),
		.out_wire_3_2(vertical_tile_17_30_to_tile_16_30_2),
		.out_wire_3_3(vertical_tile_17_30_to_tile_16_30_3),
		.in_wire_3_0(vertical_tile_16_30_to_tile_17_30_0),
		.in_wire_3_1(vertical_tile_16_30_to_tile_17_30_1),
		.in_wire_3_2(vertical_tile_16_30_to_tile_17_30_2),
		.in_wire_3_3(vertical_tile_16_30_to_tile_17_30_3),
		.out_wire_1_0(vertical_tile_17_30_to_tile_18_30_0),
		.out_wire_1_1(vertical_tile_17_30_to_tile_18_30_1),
		.out_wire_1_2(vertical_tile_17_30_to_tile_18_30_2),
		.out_wire_1_3(vertical_tile_17_30_to_tile_18_30_3),
		.in_wire_1_0(vertical_tile_18_30_to_tile_17_30_0),
		.in_wire_1_1(vertical_tile_18_30_to_tile_17_30_1),
		.in_wire_1_2(vertical_tile_18_30_to_tile_17_30_2),
		.in_wire_1_3(vertical_tile_18_30_to_tile_17_30_3),
		.out_wire_2_0(horizontal_tile_17_30_to_tile_17_29_0),
		.out_wire_2_1(horizontal_tile_17_30_to_tile_17_29_1),
		.out_wire_2_2(horizontal_tile_17_30_to_tile_17_29_2),
		.out_wire_2_3(horizontal_tile_17_30_to_tile_17_29_3),
		.in_wire_2_0(horizontal_tile_17_29_to_tile_17_30_0),
		.in_wire_2_1(horizontal_tile_17_29_to_tile_17_30_1),
		.in_wire_2_2(horizontal_tile_17_29_to_tile_17_30_2),
		.in_wire_2_3(horizontal_tile_17_29_to_tile_17_30_3),
		.out_wire_0_0(horizontal_tile_17_30_to_tile_17_31_0),
		.out_wire_0_1(horizontal_tile_17_30_to_tile_17_31_1),
		.out_wire_0_2(horizontal_tile_17_30_to_tile_17_31_2),
		.out_wire_0_3(horizontal_tile_17_30_to_tile_17_31_3),
		.in_wire_0_0(horizontal_tile_17_31_to_tile_17_30_0),
		.in_wire_0_1(horizontal_tile_17_31_to_tile_17_30_1),
		.in_wire_0_2(horizontal_tile_17_31_to_tile_17_30_2),
		.in_wire_0_3(horizontal_tile_17_31_to_tile_17_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(575)
	);

	pe_tile_right pe_tile_17_31(
		.out_wire_3_0(vertical_tile_17_31_to_tile_16_31_0),
		.out_wire_3_1(vertical_tile_17_31_to_tile_16_31_1),
		.out_wire_3_2(vertical_tile_17_31_to_tile_16_31_2),
		.out_wire_3_3(vertical_tile_17_31_to_tile_16_31_3),
		.in_wire_3_0(vertical_tile_16_31_to_tile_17_31_0),
		.in_wire_3_1(vertical_tile_16_31_to_tile_17_31_1),
		.in_wire_3_2(vertical_tile_16_31_to_tile_17_31_2),
		.in_wire_3_3(vertical_tile_16_31_to_tile_17_31_3),
		.out_wire_1_0(vertical_tile_17_31_to_tile_18_31_0),
		.out_wire_1_1(vertical_tile_17_31_to_tile_18_31_1),
		.out_wire_1_2(vertical_tile_17_31_to_tile_18_31_2),
		.out_wire_1_3(vertical_tile_17_31_to_tile_18_31_3),
		.in_wire_1_0(vertical_tile_18_31_to_tile_17_31_0),
		.in_wire_1_1(vertical_tile_18_31_to_tile_17_31_1),
		.in_wire_1_2(vertical_tile_18_31_to_tile_17_31_2),
		.in_wire_1_3(vertical_tile_18_31_to_tile_17_31_3),
		.out_wire_2_0(horizontal_tile_17_31_to_tile_17_30_0),
		.out_wire_2_1(horizontal_tile_17_31_to_tile_17_30_1),
		.out_wire_2_2(horizontal_tile_17_31_to_tile_17_30_2),
		.out_wire_2_3(horizontal_tile_17_31_to_tile_17_30_3),
		.in_wire_2_0(horizontal_tile_17_30_to_tile_17_31_0),
		.in_wire_2_1(horizontal_tile_17_30_to_tile_17_31_1),
		.in_wire_2_2(horizontal_tile_17_30_to_tile_17_31_2),
		.in_wire_2_3(horizontal_tile_17_30_to_tile_17_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(576)
	);

	pe_tile_left pe_tile_18_0(
		.out_wire_3_0(vertical_tile_18_0_to_tile_17_0_0),
		.out_wire_3_1(vertical_tile_18_0_to_tile_17_0_1),
		.out_wire_3_2(vertical_tile_18_0_to_tile_17_0_2),
		.out_wire_3_3(vertical_tile_18_0_to_tile_17_0_3),
		.in_wire_3_0(vertical_tile_17_0_to_tile_18_0_0),
		.in_wire_3_1(vertical_tile_17_0_to_tile_18_0_1),
		.in_wire_3_2(vertical_tile_17_0_to_tile_18_0_2),
		.in_wire_3_3(vertical_tile_17_0_to_tile_18_0_3),
		.out_wire_1_0(vertical_tile_18_0_to_tile_19_0_0),
		.out_wire_1_1(vertical_tile_18_0_to_tile_19_0_1),
		.out_wire_1_2(vertical_tile_18_0_to_tile_19_0_2),
		.out_wire_1_3(vertical_tile_18_0_to_tile_19_0_3),
		.in_wire_1_0(vertical_tile_19_0_to_tile_18_0_0),
		.in_wire_1_1(vertical_tile_19_0_to_tile_18_0_1),
		.in_wire_1_2(vertical_tile_19_0_to_tile_18_0_2),
		.in_wire_1_3(vertical_tile_19_0_to_tile_18_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_18_0_to_tile_18_1_0),
		.out_wire_0_1(horizontal_tile_18_0_to_tile_18_1_1),
		.out_wire_0_2(horizontal_tile_18_0_to_tile_18_1_2),
		.out_wire_0_3(horizontal_tile_18_0_to_tile_18_1_3),
		.in_wire_0_0(horizontal_tile_18_1_to_tile_18_0_0),
		.in_wire_0_1(horizontal_tile_18_1_to_tile_18_0_1),
		.in_wire_0_2(horizontal_tile_18_1_to_tile_18_0_2),
		.in_wire_0_3(horizontal_tile_18_1_to_tile_18_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(577)
	);

	pe_tile pe_tile_18_1(
		.out_wire_3_0(vertical_tile_18_1_to_tile_17_1_0),
		.out_wire_3_1(vertical_tile_18_1_to_tile_17_1_1),
		.out_wire_3_2(vertical_tile_18_1_to_tile_17_1_2),
		.out_wire_3_3(vertical_tile_18_1_to_tile_17_1_3),
		.in_wire_3_0(vertical_tile_17_1_to_tile_18_1_0),
		.in_wire_3_1(vertical_tile_17_1_to_tile_18_1_1),
		.in_wire_3_2(vertical_tile_17_1_to_tile_18_1_2),
		.in_wire_3_3(vertical_tile_17_1_to_tile_18_1_3),
		.out_wire_1_0(vertical_tile_18_1_to_tile_19_1_0),
		.out_wire_1_1(vertical_tile_18_1_to_tile_19_1_1),
		.out_wire_1_2(vertical_tile_18_1_to_tile_19_1_2),
		.out_wire_1_3(vertical_tile_18_1_to_tile_19_1_3),
		.in_wire_1_0(vertical_tile_19_1_to_tile_18_1_0),
		.in_wire_1_1(vertical_tile_19_1_to_tile_18_1_1),
		.in_wire_1_2(vertical_tile_19_1_to_tile_18_1_2),
		.in_wire_1_3(vertical_tile_19_1_to_tile_18_1_3),
		.out_wire_2_0(horizontal_tile_18_1_to_tile_18_0_0),
		.out_wire_2_1(horizontal_tile_18_1_to_tile_18_0_1),
		.out_wire_2_2(horizontal_tile_18_1_to_tile_18_0_2),
		.out_wire_2_3(horizontal_tile_18_1_to_tile_18_0_3),
		.in_wire_2_0(horizontal_tile_18_0_to_tile_18_1_0),
		.in_wire_2_1(horizontal_tile_18_0_to_tile_18_1_1),
		.in_wire_2_2(horizontal_tile_18_0_to_tile_18_1_2),
		.in_wire_2_3(horizontal_tile_18_0_to_tile_18_1_3),
		.out_wire_0_0(horizontal_tile_18_1_to_tile_18_2_0),
		.out_wire_0_1(horizontal_tile_18_1_to_tile_18_2_1),
		.out_wire_0_2(horizontal_tile_18_1_to_tile_18_2_2),
		.out_wire_0_3(horizontal_tile_18_1_to_tile_18_2_3),
		.in_wire_0_0(horizontal_tile_18_2_to_tile_18_1_0),
		.in_wire_0_1(horizontal_tile_18_2_to_tile_18_1_1),
		.in_wire_0_2(horizontal_tile_18_2_to_tile_18_1_2),
		.in_wire_0_3(horizontal_tile_18_2_to_tile_18_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(578)
	);

	pe_tile pe_tile_18_2(
		.out_wire_3_0(vertical_tile_18_2_to_tile_17_2_0),
		.out_wire_3_1(vertical_tile_18_2_to_tile_17_2_1),
		.out_wire_3_2(vertical_tile_18_2_to_tile_17_2_2),
		.out_wire_3_3(vertical_tile_18_2_to_tile_17_2_3),
		.in_wire_3_0(vertical_tile_17_2_to_tile_18_2_0),
		.in_wire_3_1(vertical_tile_17_2_to_tile_18_2_1),
		.in_wire_3_2(vertical_tile_17_2_to_tile_18_2_2),
		.in_wire_3_3(vertical_tile_17_2_to_tile_18_2_3),
		.out_wire_1_0(vertical_tile_18_2_to_tile_19_2_0),
		.out_wire_1_1(vertical_tile_18_2_to_tile_19_2_1),
		.out_wire_1_2(vertical_tile_18_2_to_tile_19_2_2),
		.out_wire_1_3(vertical_tile_18_2_to_tile_19_2_3),
		.in_wire_1_0(vertical_tile_19_2_to_tile_18_2_0),
		.in_wire_1_1(vertical_tile_19_2_to_tile_18_2_1),
		.in_wire_1_2(vertical_tile_19_2_to_tile_18_2_2),
		.in_wire_1_3(vertical_tile_19_2_to_tile_18_2_3),
		.out_wire_2_0(horizontal_tile_18_2_to_tile_18_1_0),
		.out_wire_2_1(horizontal_tile_18_2_to_tile_18_1_1),
		.out_wire_2_2(horizontal_tile_18_2_to_tile_18_1_2),
		.out_wire_2_3(horizontal_tile_18_2_to_tile_18_1_3),
		.in_wire_2_0(horizontal_tile_18_1_to_tile_18_2_0),
		.in_wire_2_1(horizontal_tile_18_1_to_tile_18_2_1),
		.in_wire_2_2(horizontal_tile_18_1_to_tile_18_2_2),
		.in_wire_2_3(horizontal_tile_18_1_to_tile_18_2_3),
		.out_wire_0_0(horizontal_tile_18_2_to_tile_18_3_0),
		.out_wire_0_1(horizontal_tile_18_2_to_tile_18_3_1),
		.out_wire_0_2(horizontal_tile_18_2_to_tile_18_3_2),
		.out_wire_0_3(horizontal_tile_18_2_to_tile_18_3_3),
		.in_wire_0_0(horizontal_tile_18_3_to_tile_18_2_0),
		.in_wire_0_1(horizontal_tile_18_3_to_tile_18_2_1),
		.in_wire_0_2(horizontal_tile_18_3_to_tile_18_2_2),
		.in_wire_0_3(horizontal_tile_18_3_to_tile_18_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(579)
	);

	pe_tile pe_tile_18_3(
		.out_wire_3_0(vertical_tile_18_3_to_tile_17_3_0),
		.out_wire_3_1(vertical_tile_18_3_to_tile_17_3_1),
		.out_wire_3_2(vertical_tile_18_3_to_tile_17_3_2),
		.out_wire_3_3(vertical_tile_18_3_to_tile_17_3_3),
		.in_wire_3_0(vertical_tile_17_3_to_tile_18_3_0),
		.in_wire_3_1(vertical_tile_17_3_to_tile_18_3_1),
		.in_wire_3_2(vertical_tile_17_3_to_tile_18_3_2),
		.in_wire_3_3(vertical_tile_17_3_to_tile_18_3_3),
		.out_wire_1_0(vertical_tile_18_3_to_tile_19_3_0),
		.out_wire_1_1(vertical_tile_18_3_to_tile_19_3_1),
		.out_wire_1_2(vertical_tile_18_3_to_tile_19_3_2),
		.out_wire_1_3(vertical_tile_18_3_to_tile_19_3_3),
		.in_wire_1_0(vertical_tile_19_3_to_tile_18_3_0),
		.in_wire_1_1(vertical_tile_19_3_to_tile_18_3_1),
		.in_wire_1_2(vertical_tile_19_3_to_tile_18_3_2),
		.in_wire_1_3(vertical_tile_19_3_to_tile_18_3_3),
		.out_wire_2_0(horizontal_tile_18_3_to_tile_18_2_0),
		.out_wire_2_1(horizontal_tile_18_3_to_tile_18_2_1),
		.out_wire_2_2(horizontal_tile_18_3_to_tile_18_2_2),
		.out_wire_2_3(horizontal_tile_18_3_to_tile_18_2_3),
		.in_wire_2_0(horizontal_tile_18_2_to_tile_18_3_0),
		.in_wire_2_1(horizontal_tile_18_2_to_tile_18_3_1),
		.in_wire_2_2(horizontal_tile_18_2_to_tile_18_3_2),
		.in_wire_2_3(horizontal_tile_18_2_to_tile_18_3_3),
		.out_wire_0_0(horizontal_tile_18_3_to_tile_18_4_0),
		.out_wire_0_1(horizontal_tile_18_3_to_tile_18_4_1),
		.out_wire_0_2(horizontal_tile_18_3_to_tile_18_4_2),
		.out_wire_0_3(horizontal_tile_18_3_to_tile_18_4_3),
		.in_wire_0_0(horizontal_tile_18_4_to_tile_18_3_0),
		.in_wire_0_1(horizontal_tile_18_4_to_tile_18_3_1),
		.in_wire_0_2(horizontal_tile_18_4_to_tile_18_3_2),
		.in_wire_0_3(horizontal_tile_18_4_to_tile_18_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(580)
	);

	pe_tile pe_tile_18_4(
		.out_wire_3_0(vertical_tile_18_4_to_tile_17_4_0),
		.out_wire_3_1(vertical_tile_18_4_to_tile_17_4_1),
		.out_wire_3_2(vertical_tile_18_4_to_tile_17_4_2),
		.out_wire_3_3(vertical_tile_18_4_to_tile_17_4_3),
		.in_wire_3_0(vertical_tile_17_4_to_tile_18_4_0),
		.in_wire_3_1(vertical_tile_17_4_to_tile_18_4_1),
		.in_wire_3_2(vertical_tile_17_4_to_tile_18_4_2),
		.in_wire_3_3(vertical_tile_17_4_to_tile_18_4_3),
		.out_wire_1_0(vertical_tile_18_4_to_tile_19_4_0),
		.out_wire_1_1(vertical_tile_18_4_to_tile_19_4_1),
		.out_wire_1_2(vertical_tile_18_4_to_tile_19_4_2),
		.out_wire_1_3(vertical_tile_18_4_to_tile_19_4_3),
		.in_wire_1_0(vertical_tile_19_4_to_tile_18_4_0),
		.in_wire_1_1(vertical_tile_19_4_to_tile_18_4_1),
		.in_wire_1_2(vertical_tile_19_4_to_tile_18_4_2),
		.in_wire_1_3(vertical_tile_19_4_to_tile_18_4_3),
		.out_wire_2_0(horizontal_tile_18_4_to_tile_18_3_0),
		.out_wire_2_1(horizontal_tile_18_4_to_tile_18_3_1),
		.out_wire_2_2(horizontal_tile_18_4_to_tile_18_3_2),
		.out_wire_2_3(horizontal_tile_18_4_to_tile_18_3_3),
		.in_wire_2_0(horizontal_tile_18_3_to_tile_18_4_0),
		.in_wire_2_1(horizontal_tile_18_3_to_tile_18_4_1),
		.in_wire_2_2(horizontal_tile_18_3_to_tile_18_4_2),
		.in_wire_2_3(horizontal_tile_18_3_to_tile_18_4_3),
		.out_wire_0_0(horizontal_tile_18_4_to_tile_18_5_0),
		.out_wire_0_1(horizontal_tile_18_4_to_tile_18_5_1),
		.out_wire_0_2(horizontal_tile_18_4_to_tile_18_5_2),
		.out_wire_0_3(horizontal_tile_18_4_to_tile_18_5_3),
		.in_wire_0_0(horizontal_tile_18_5_to_tile_18_4_0),
		.in_wire_0_1(horizontal_tile_18_5_to_tile_18_4_1),
		.in_wire_0_2(horizontal_tile_18_5_to_tile_18_4_2),
		.in_wire_0_3(horizontal_tile_18_5_to_tile_18_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(581)
	);

	pe_tile pe_tile_18_5(
		.out_wire_3_0(vertical_tile_18_5_to_tile_17_5_0),
		.out_wire_3_1(vertical_tile_18_5_to_tile_17_5_1),
		.out_wire_3_2(vertical_tile_18_5_to_tile_17_5_2),
		.out_wire_3_3(vertical_tile_18_5_to_tile_17_5_3),
		.in_wire_3_0(vertical_tile_17_5_to_tile_18_5_0),
		.in_wire_3_1(vertical_tile_17_5_to_tile_18_5_1),
		.in_wire_3_2(vertical_tile_17_5_to_tile_18_5_2),
		.in_wire_3_3(vertical_tile_17_5_to_tile_18_5_3),
		.out_wire_1_0(vertical_tile_18_5_to_tile_19_5_0),
		.out_wire_1_1(vertical_tile_18_5_to_tile_19_5_1),
		.out_wire_1_2(vertical_tile_18_5_to_tile_19_5_2),
		.out_wire_1_3(vertical_tile_18_5_to_tile_19_5_3),
		.in_wire_1_0(vertical_tile_19_5_to_tile_18_5_0),
		.in_wire_1_1(vertical_tile_19_5_to_tile_18_5_1),
		.in_wire_1_2(vertical_tile_19_5_to_tile_18_5_2),
		.in_wire_1_3(vertical_tile_19_5_to_tile_18_5_3),
		.out_wire_2_0(horizontal_tile_18_5_to_tile_18_4_0),
		.out_wire_2_1(horizontal_tile_18_5_to_tile_18_4_1),
		.out_wire_2_2(horizontal_tile_18_5_to_tile_18_4_2),
		.out_wire_2_3(horizontal_tile_18_5_to_tile_18_4_3),
		.in_wire_2_0(horizontal_tile_18_4_to_tile_18_5_0),
		.in_wire_2_1(horizontal_tile_18_4_to_tile_18_5_1),
		.in_wire_2_2(horizontal_tile_18_4_to_tile_18_5_2),
		.in_wire_2_3(horizontal_tile_18_4_to_tile_18_5_3),
		.out_wire_0_0(horizontal_tile_18_5_to_tile_18_6_0),
		.out_wire_0_1(horizontal_tile_18_5_to_tile_18_6_1),
		.out_wire_0_2(horizontal_tile_18_5_to_tile_18_6_2),
		.out_wire_0_3(horizontal_tile_18_5_to_tile_18_6_3),
		.in_wire_0_0(horizontal_tile_18_6_to_tile_18_5_0),
		.in_wire_0_1(horizontal_tile_18_6_to_tile_18_5_1),
		.in_wire_0_2(horizontal_tile_18_6_to_tile_18_5_2),
		.in_wire_0_3(horizontal_tile_18_6_to_tile_18_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(582)
	);

	pe_tile pe_tile_18_6(
		.out_wire_3_0(vertical_tile_18_6_to_tile_17_6_0),
		.out_wire_3_1(vertical_tile_18_6_to_tile_17_6_1),
		.out_wire_3_2(vertical_tile_18_6_to_tile_17_6_2),
		.out_wire_3_3(vertical_tile_18_6_to_tile_17_6_3),
		.in_wire_3_0(vertical_tile_17_6_to_tile_18_6_0),
		.in_wire_3_1(vertical_tile_17_6_to_tile_18_6_1),
		.in_wire_3_2(vertical_tile_17_6_to_tile_18_6_2),
		.in_wire_3_3(vertical_tile_17_6_to_tile_18_6_3),
		.out_wire_1_0(vertical_tile_18_6_to_tile_19_6_0),
		.out_wire_1_1(vertical_tile_18_6_to_tile_19_6_1),
		.out_wire_1_2(vertical_tile_18_6_to_tile_19_6_2),
		.out_wire_1_3(vertical_tile_18_6_to_tile_19_6_3),
		.in_wire_1_0(vertical_tile_19_6_to_tile_18_6_0),
		.in_wire_1_1(vertical_tile_19_6_to_tile_18_6_1),
		.in_wire_1_2(vertical_tile_19_6_to_tile_18_6_2),
		.in_wire_1_3(vertical_tile_19_6_to_tile_18_6_3),
		.out_wire_2_0(horizontal_tile_18_6_to_tile_18_5_0),
		.out_wire_2_1(horizontal_tile_18_6_to_tile_18_5_1),
		.out_wire_2_2(horizontal_tile_18_6_to_tile_18_5_2),
		.out_wire_2_3(horizontal_tile_18_6_to_tile_18_5_3),
		.in_wire_2_0(horizontal_tile_18_5_to_tile_18_6_0),
		.in_wire_2_1(horizontal_tile_18_5_to_tile_18_6_1),
		.in_wire_2_2(horizontal_tile_18_5_to_tile_18_6_2),
		.in_wire_2_3(horizontal_tile_18_5_to_tile_18_6_3),
		.out_wire_0_0(horizontal_tile_18_6_to_tile_18_7_0),
		.out_wire_0_1(horizontal_tile_18_6_to_tile_18_7_1),
		.out_wire_0_2(horizontal_tile_18_6_to_tile_18_7_2),
		.out_wire_0_3(horizontal_tile_18_6_to_tile_18_7_3),
		.in_wire_0_0(horizontal_tile_18_7_to_tile_18_6_0),
		.in_wire_0_1(horizontal_tile_18_7_to_tile_18_6_1),
		.in_wire_0_2(horizontal_tile_18_7_to_tile_18_6_2),
		.in_wire_0_3(horizontal_tile_18_7_to_tile_18_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(583)
	);

	pe_tile pe_tile_18_7(
		.out_wire_3_0(vertical_tile_18_7_to_tile_17_7_0),
		.out_wire_3_1(vertical_tile_18_7_to_tile_17_7_1),
		.out_wire_3_2(vertical_tile_18_7_to_tile_17_7_2),
		.out_wire_3_3(vertical_tile_18_7_to_tile_17_7_3),
		.in_wire_3_0(vertical_tile_17_7_to_tile_18_7_0),
		.in_wire_3_1(vertical_tile_17_7_to_tile_18_7_1),
		.in_wire_3_2(vertical_tile_17_7_to_tile_18_7_2),
		.in_wire_3_3(vertical_tile_17_7_to_tile_18_7_3),
		.out_wire_1_0(vertical_tile_18_7_to_tile_19_7_0),
		.out_wire_1_1(vertical_tile_18_7_to_tile_19_7_1),
		.out_wire_1_2(vertical_tile_18_7_to_tile_19_7_2),
		.out_wire_1_3(vertical_tile_18_7_to_tile_19_7_3),
		.in_wire_1_0(vertical_tile_19_7_to_tile_18_7_0),
		.in_wire_1_1(vertical_tile_19_7_to_tile_18_7_1),
		.in_wire_1_2(vertical_tile_19_7_to_tile_18_7_2),
		.in_wire_1_3(vertical_tile_19_7_to_tile_18_7_3),
		.out_wire_2_0(horizontal_tile_18_7_to_tile_18_6_0),
		.out_wire_2_1(horizontal_tile_18_7_to_tile_18_6_1),
		.out_wire_2_2(horizontal_tile_18_7_to_tile_18_6_2),
		.out_wire_2_3(horizontal_tile_18_7_to_tile_18_6_3),
		.in_wire_2_0(horizontal_tile_18_6_to_tile_18_7_0),
		.in_wire_2_1(horizontal_tile_18_6_to_tile_18_7_1),
		.in_wire_2_2(horizontal_tile_18_6_to_tile_18_7_2),
		.in_wire_2_3(horizontal_tile_18_6_to_tile_18_7_3),
		.out_wire_0_0(horizontal_tile_18_7_to_tile_18_8_0),
		.out_wire_0_1(horizontal_tile_18_7_to_tile_18_8_1),
		.out_wire_0_2(horizontal_tile_18_7_to_tile_18_8_2),
		.out_wire_0_3(horizontal_tile_18_7_to_tile_18_8_3),
		.in_wire_0_0(horizontal_tile_18_8_to_tile_18_7_0),
		.in_wire_0_1(horizontal_tile_18_8_to_tile_18_7_1),
		.in_wire_0_2(horizontal_tile_18_8_to_tile_18_7_2),
		.in_wire_0_3(horizontal_tile_18_8_to_tile_18_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(584)
	);

	pe_tile pe_tile_18_8(
		.out_wire_3_0(vertical_tile_18_8_to_tile_17_8_0),
		.out_wire_3_1(vertical_tile_18_8_to_tile_17_8_1),
		.out_wire_3_2(vertical_tile_18_8_to_tile_17_8_2),
		.out_wire_3_3(vertical_tile_18_8_to_tile_17_8_3),
		.in_wire_3_0(vertical_tile_17_8_to_tile_18_8_0),
		.in_wire_3_1(vertical_tile_17_8_to_tile_18_8_1),
		.in_wire_3_2(vertical_tile_17_8_to_tile_18_8_2),
		.in_wire_3_3(vertical_tile_17_8_to_tile_18_8_3),
		.out_wire_1_0(vertical_tile_18_8_to_tile_19_8_0),
		.out_wire_1_1(vertical_tile_18_8_to_tile_19_8_1),
		.out_wire_1_2(vertical_tile_18_8_to_tile_19_8_2),
		.out_wire_1_3(vertical_tile_18_8_to_tile_19_8_3),
		.in_wire_1_0(vertical_tile_19_8_to_tile_18_8_0),
		.in_wire_1_1(vertical_tile_19_8_to_tile_18_8_1),
		.in_wire_1_2(vertical_tile_19_8_to_tile_18_8_2),
		.in_wire_1_3(vertical_tile_19_8_to_tile_18_8_3),
		.out_wire_2_0(horizontal_tile_18_8_to_tile_18_7_0),
		.out_wire_2_1(horizontal_tile_18_8_to_tile_18_7_1),
		.out_wire_2_2(horizontal_tile_18_8_to_tile_18_7_2),
		.out_wire_2_3(horizontal_tile_18_8_to_tile_18_7_3),
		.in_wire_2_0(horizontal_tile_18_7_to_tile_18_8_0),
		.in_wire_2_1(horizontal_tile_18_7_to_tile_18_8_1),
		.in_wire_2_2(horizontal_tile_18_7_to_tile_18_8_2),
		.in_wire_2_3(horizontal_tile_18_7_to_tile_18_8_3),
		.out_wire_0_0(horizontal_tile_18_8_to_tile_18_9_0),
		.out_wire_0_1(horizontal_tile_18_8_to_tile_18_9_1),
		.out_wire_0_2(horizontal_tile_18_8_to_tile_18_9_2),
		.out_wire_0_3(horizontal_tile_18_8_to_tile_18_9_3),
		.in_wire_0_0(horizontal_tile_18_9_to_tile_18_8_0),
		.in_wire_0_1(horizontal_tile_18_9_to_tile_18_8_1),
		.in_wire_0_2(horizontal_tile_18_9_to_tile_18_8_2),
		.in_wire_0_3(horizontal_tile_18_9_to_tile_18_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(585)
	);

	pe_tile pe_tile_18_9(
		.out_wire_3_0(vertical_tile_18_9_to_tile_17_9_0),
		.out_wire_3_1(vertical_tile_18_9_to_tile_17_9_1),
		.out_wire_3_2(vertical_tile_18_9_to_tile_17_9_2),
		.out_wire_3_3(vertical_tile_18_9_to_tile_17_9_3),
		.in_wire_3_0(vertical_tile_17_9_to_tile_18_9_0),
		.in_wire_3_1(vertical_tile_17_9_to_tile_18_9_1),
		.in_wire_3_2(vertical_tile_17_9_to_tile_18_9_2),
		.in_wire_3_3(vertical_tile_17_9_to_tile_18_9_3),
		.out_wire_1_0(vertical_tile_18_9_to_tile_19_9_0),
		.out_wire_1_1(vertical_tile_18_9_to_tile_19_9_1),
		.out_wire_1_2(vertical_tile_18_9_to_tile_19_9_2),
		.out_wire_1_3(vertical_tile_18_9_to_tile_19_9_3),
		.in_wire_1_0(vertical_tile_19_9_to_tile_18_9_0),
		.in_wire_1_1(vertical_tile_19_9_to_tile_18_9_1),
		.in_wire_1_2(vertical_tile_19_9_to_tile_18_9_2),
		.in_wire_1_3(vertical_tile_19_9_to_tile_18_9_3),
		.out_wire_2_0(horizontal_tile_18_9_to_tile_18_8_0),
		.out_wire_2_1(horizontal_tile_18_9_to_tile_18_8_1),
		.out_wire_2_2(horizontal_tile_18_9_to_tile_18_8_2),
		.out_wire_2_3(horizontal_tile_18_9_to_tile_18_8_3),
		.in_wire_2_0(horizontal_tile_18_8_to_tile_18_9_0),
		.in_wire_2_1(horizontal_tile_18_8_to_tile_18_9_1),
		.in_wire_2_2(horizontal_tile_18_8_to_tile_18_9_2),
		.in_wire_2_3(horizontal_tile_18_8_to_tile_18_9_3),
		.out_wire_0_0(horizontal_tile_18_9_to_tile_18_10_0),
		.out_wire_0_1(horizontal_tile_18_9_to_tile_18_10_1),
		.out_wire_0_2(horizontal_tile_18_9_to_tile_18_10_2),
		.out_wire_0_3(horizontal_tile_18_9_to_tile_18_10_3),
		.in_wire_0_0(horizontal_tile_18_10_to_tile_18_9_0),
		.in_wire_0_1(horizontal_tile_18_10_to_tile_18_9_1),
		.in_wire_0_2(horizontal_tile_18_10_to_tile_18_9_2),
		.in_wire_0_3(horizontal_tile_18_10_to_tile_18_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(586)
	);

	pe_tile pe_tile_18_10(
		.out_wire_3_0(vertical_tile_18_10_to_tile_17_10_0),
		.out_wire_3_1(vertical_tile_18_10_to_tile_17_10_1),
		.out_wire_3_2(vertical_tile_18_10_to_tile_17_10_2),
		.out_wire_3_3(vertical_tile_18_10_to_tile_17_10_3),
		.in_wire_3_0(vertical_tile_17_10_to_tile_18_10_0),
		.in_wire_3_1(vertical_tile_17_10_to_tile_18_10_1),
		.in_wire_3_2(vertical_tile_17_10_to_tile_18_10_2),
		.in_wire_3_3(vertical_tile_17_10_to_tile_18_10_3),
		.out_wire_1_0(vertical_tile_18_10_to_tile_19_10_0),
		.out_wire_1_1(vertical_tile_18_10_to_tile_19_10_1),
		.out_wire_1_2(vertical_tile_18_10_to_tile_19_10_2),
		.out_wire_1_3(vertical_tile_18_10_to_tile_19_10_3),
		.in_wire_1_0(vertical_tile_19_10_to_tile_18_10_0),
		.in_wire_1_1(vertical_tile_19_10_to_tile_18_10_1),
		.in_wire_1_2(vertical_tile_19_10_to_tile_18_10_2),
		.in_wire_1_3(vertical_tile_19_10_to_tile_18_10_3),
		.out_wire_2_0(horizontal_tile_18_10_to_tile_18_9_0),
		.out_wire_2_1(horizontal_tile_18_10_to_tile_18_9_1),
		.out_wire_2_2(horizontal_tile_18_10_to_tile_18_9_2),
		.out_wire_2_3(horizontal_tile_18_10_to_tile_18_9_3),
		.in_wire_2_0(horizontal_tile_18_9_to_tile_18_10_0),
		.in_wire_2_1(horizontal_tile_18_9_to_tile_18_10_1),
		.in_wire_2_2(horizontal_tile_18_9_to_tile_18_10_2),
		.in_wire_2_3(horizontal_tile_18_9_to_tile_18_10_3),
		.out_wire_0_0(horizontal_tile_18_10_to_tile_18_11_0),
		.out_wire_0_1(horizontal_tile_18_10_to_tile_18_11_1),
		.out_wire_0_2(horizontal_tile_18_10_to_tile_18_11_2),
		.out_wire_0_3(horizontal_tile_18_10_to_tile_18_11_3),
		.in_wire_0_0(horizontal_tile_18_11_to_tile_18_10_0),
		.in_wire_0_1(horizontal_tile_18_11_to_tile_18_10_1),
		.in_wire_0_2(horizontal_tile_18_11_to_tile_18_10_2),
		.in_wire_0_3(horizontal_tile_18_11_to_tile_18_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(587)
	);

	pe_tile pe_tile_18_11(
		.out_wire_3_0(vertical_tile_18_11_to_tile_17_11_0),
		.out_wire_3_1(vertical_tile_18_11_to_tile_17_11_1),
		.out_wire_3_2(vertical_tile_18_11_to_tile_17_11_2),
		.out_wire_3_3(vertical_tile_18_11_to_tile_17_11_3),
		.in_wire_3_0(vertical_tile_17_11_to_tile_18_11_0),
		.in_wire_3_1(vertical_tile_17_11_to_tile_18_11_1),
		.in_wire_3_2(vertical_tile_17_11_to_tile_18_11_2),
		.in_wire_3_3(vertical_tile_17_11_to_tile_18_11_3),
		.out_wire_1_0(vertical_tile_18_11_to_tile_19_11_0),
		.out_wire_1_1(vertical_tile_18_11_to_tile_19_11_1),
		.out_wire_1_2(vertical_tile_18_11_to_tile_19_11_2),
		.out_wire_1_3(vertical_tile_18_11_to_tile_19_11_3),
		.in_wire_1_0(vertical_tile_19_11_to_tile_18_11_0),
		.in_wire_1_1(vertical_tile_19_11_to_tile_18_11_1),
		.in_wire_1_2(vertical_tile_19_11_to_tile_18_11_2),
		.in_wire_1_3(vertical_tile_19_11_to_tile_18_11_3),
		.out_wire_2_0(horizontal_tile_18_11_to_tile_18_10_0),
		.out_wire_2_1(horizontal_tile_18_11_to_tile_18_10_1),
		.out_wire_2_2(horizontal_tile_18_11_to_tile_18_10_2),
		.out_wire_2_3(horizontal_tile_18_11_to_tile_18_10_3),
		.in_wire_2_0(horizontal_tile_18_10_to_tile_18_11_0),
		.in_wire_2_1(horizontal_tile_18_10_to_tile_18_11_1),
		.in_wire_2_2(horizontal_tile_18_10_to_tile_18_11_2),
		.in_wire_2_3(horizontal_tile_18_10_to_tile_18_11_3),
		.out_wire_0_0(horizontal_tile_18_11_to_tile_18_12_0),
		.out_wire_0_1(horizontal_tile_18_11_to_tile_18_12_1),
		.out_wire_0_2(horizontal_tile_18_11_to_tile_18_12_2),
		.out_wire_0_3(horizontal_tile_18_11_to_tile_18_12_3),
		.in_wire_0_0(horizontal_tile_18_12_to_tile_18_11_0),
		.in_wire_0_1(horizontal_tile_18_12_to_tile_18_11_1),
		.in_wire_0_2(horizontal_tile_18_12_to_tile_18_11_2),
		.in_wire_0_3(horizontal_tile_18_12_to_tile_18_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(588)
	);

	pe_tile pe_tile_18_12(
		.out_wire_3_0(vertical_tile_18_12_to_tile_17_12_0),
		.out_wire_3_1(vertical_tile_18_12_to_tile_17_12_1),
		.out_wire_3_2(vertical_tile_18_12_to_tile_17_12_2),
		.out_wire_3_3(vertical_tile_18_12_to_tile_17_12_3),
		.in_wire_3_0(vertical_tile_17_12_to_tile_18_12_0),
		.in_wire_3_1(vertical_tile_17_12_to_tile_18_12_1),
		.in_wire_3_2(vertical_tile_17_12_to_tile_18_12_2),
		.in_wire_3_3(vertical_tile_17_12_to_tile_18_12_3),
		.out_wire_1_0(vertical_tile_18_12_to_tile_19_12_0),
		.out_wire_1_1(vertical_tile_18_12_to_tile_19_12_1),
		.out_wire_1_2(vertical_tile_18_12_to_tile_19_12_2),
		.out_wire_1_3(vertical_tile_18_12_to_tile_19_12_3),
		.in_wire_1_0(vertical_tile_19_12_to_tile_18_12_0),
		.in_wire_1_1(vertical_tile_19_12_to_tile_18_12_1),
		.in_wire_1_2(vertical_tile_19_12_to_tile_18_12_2),
		.in_wire_1_3(vertical_tile_19_12_to_tile_18_12_3),
		.out_wire_2_0(horizontal_tile_18_12_to_tile_18_11_0),
		.out_wire_2_1(horizontal_tile_18_12_to_tile_18_11_1),
		.out_wire_2_2(horizontal_tile_18_12_to_tile_18_11_2),
		.out_wire_2_3(horizontal_tile_18_12_to_tile_18_11_3),
		.in_wire_2_0(horizontal_tile_18_11_to_tile_18_12_0),
		.in_wire_2_1(horizontal_tile_18_11_to_tile_18_12_1),
		.in_wire_2_2(horizontal_tile_18_11_to_tile_18_12_2),
		.in_wire_2_3(horizontal_tile_18_11_to_tile_18_12_3),
		.out_wire_0_0(horizontal_tile_18_12_to_tile_18_13_0),
		.out_wire_0_1(horizontal_tile_18_12_to_tile_18_13_1),
		.out_wire_0_2(horizontal_tile_18_12_to_tile_18_13_2),
		.out_wire_0_3(horizontal_tile_18_12_to_tile_18_13_3),
		.in_wire_0_0(horizontal_tile_18_13_to_tile_18_12_0),
		.in_wire_0_1(horizontal_tile_18_13_to_tile_18_12_1),
		.in_wire_0_2(horizontal_tile_18_13_to_tile_18_12_2),
		.in_wire_0_3(horizontal_tile_18_13_to_tile_18_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(589)
	);

	pe_tile pe_tile_18_13(
		.out_wire_3_0(vertical_tile_18_13_to_tile_17_13_0),
		.out_wire_3_1(vertical_tile_18_13_to_tile_17_13_1),
		.out_wire_3_2(vertical_tile_18_13_to_tile_17_13_2),
		.out_wire_3_3(vertical_tile_18_13_to_tile_17_13_3),
		.in_wire_3_0(vertical_tile_17_13_to_tile_18_13_0),
		.in_wire_3_1(vertical_tile_17_13_to_tile_18_13_1),
		.in_wire_3_2(vertical_tile_17_13_to_tile_18_13_2),
		.in_wire_3_3(vertical_tile_17_13_to_tile_18_13_3),
		.out_wire_1_0(vertical_tile_18_13_to_tile_19_13_0),
		.out_wire_1_1(vertical_tile_18_13_to_tile_19_13_1),
		.out_wire_1_2(vertical_tile_18_13_to_tile_19_13_2),
		.out_wire_1_3(vertical_tile_18_13_to_tile_19_13_3),
		.in_wire_1_0(vertical_tile_19_13_to_tile_18_13_0),
		.in_wire_1_1(vertical_tile_19_13_to_tile_18_13_1),
		.in_wire_1_2(vertical_tile_19_13_to_tile_18_13_2),
		.in_wire_1_3(vertical_tile_19_13_to_tile_18_13_3),
		.out_wire_2_0(horizontal_tile_18_13_to_tile_18_12_0),
		.out_wire_2_1(horizontal_tile_18_13_to_tile_18_12_1),
		.out_wire_2_2(horizontal_tile_18_13_to_tile_18_12_2),
		.out_wire_2_3(horizontal_tile_18_13_to_tile_18_12_3),
		.in_wire_2_0(horizontal_tile_18_12_to_tile_18_13_0),
		.in_wire_2_1(horizontal_tile_18_12_to_tile_18_13_1),
		.in_wire_2_2(horizontal_tile_18_12_to_tile_18_13_2),
		.in_wire_2_3(horizontal_tile_18_12_to_tile_18_13_3),
		.out_wire_0_0(horizontal_tile_18_13_to_tile_18_14_0),
		.out_wire_0_1(horizontal_tile_18_13_to_tile_18_14_1),
		.out_wire_0_2(horizontal_tile_18_13_to_tile_18_14_2),
		.out_wire_0_3(horizontal_tile_18_13_to_tile_18_14_3),
		.in_wire_0_0(horizontal_tile_18_14_to_tile_18_13_0),
		.in_wire_0_1(horizontal_tile_18_14_to_tile_18_13_1),
		.in_wire_0_2(horizontal_tile_18_14_to_tile_18_13_2),
		.in_wire_0_3(horizontal_tile_18_14_to_tile_18_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(590)
	);

	pe_tile pe_tile_18_14(
		.out_wire_3_0(vertical_tile_18_14_to_tile_17_14_0),
		.out_wire_3_1(vertical_tile_18_14_to_tile_17_14_1),
		.out_wire_3_2(vertical_tile_18_14_to_tile_17_14_2),
		.out_wire_3_3(vertical_tile_18_14_to_tile_17_14_3),
		.in_wire_3_0(vertical_tile_17_14_to_tile_18_14_0),
		.in_wire_3_1(vertical_tile_17_14_to_tile_18_14_1),
		.in_wire_3_2(vertical_tile_17_14_to_tile_18_14_2),
		.in_wire_3_3(vertical_tile_17_14_to_tile_18_14_3),
		.out_wire_1_0(vertical_tile_18_14_to_tile_19_14_0),
		.out_wire_1_1(vertical_tile_18_14_to_tile_19_14_1),
		.out_wire_1_2(vertical_tile_18_14_to_tile_19_14_2),
		.out_wire_1_3(vertical_tile_18_14_to_tile_19_14_3),
		.in_wire_1_0(vertical_tile_19_14_to_tile_18_14_0),
		.in_wire_1_1(vertical_tile_19_14_to_tile_18_14_1),
		.in_wire_1_2(vertical_tile_19_14_to_tile_18_14_2),
		.in_wire_1_3(vertical_tile_19_14_to_tile_18_14_3),
		.out_wire_2_0(horizontal_tile_18_14_to_tile_18_13_0),
		.out_wire_2_1(horizontal_tile_18_14_to_tile_18_13_1),
		.out_wire_2_2(horizontal_tile_18_14_to_tile_18_13_2),
		.out_wire_2_3(horizontal_tile_18_14_to_tile_18_13_3),
		.in_wire_2_0(horizontal_tile_18_13_to_tile_18_14_0),
		.in_wire_2_1(horizontal_tile_18_13_to_tile_18_14_1),
		.in_wire_2_2(horizontal_tile_18_13_to_tile_18_14_2),
		.in_wire_2_3(horizontal_tile_18_13_to_tile_18_14_3),
		.out_wire_0_0(horizontal_tile_18_14_to_tile_18_15_0),
		.out_wire_0_1(horizontal_tile_18_14_to_tile_18_15_1),
		.out_wire_0_2(horizontal_tile_18_14_to_tile_18_15_2),
		.out_wire_0_3(horizontal_tile_18_14_to_tile_18_15_3),
		.in_wire_0_0(horizontal_tile_18_15_to_tile_18_14_0),
		.in_wire_0_1(horizontal_tile_18_15_to_tile_18_14_1),
		.in_wire_0_2(horizontal_tile_18_15_to_tile_18_14_2),
		.in_wire_0_3(horizontal_tile_18_15_to_tile_18_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(591)
	);

	pe_tile pe_tile_18_15(
		.out_wire_3_0(vertical_tile_18_15_to_tile_17_15_0),
		.out_wire_3_1(vertical_tile_18_15_to_tile_17_15_1),
		.out_wire_3_2(vertical_tile_18_15_to_tile_17_15_2),
		.out_wire_3_3(vertical_tile_18_15_to_tile_17_15_3),
		.in_wire_3_0(vertical_tile_17_15_to_tile_18_15_0),
		.in_wire_3_1(vertical_tile_17_15_to_tile_18_15_1),
		.in_wire_3_2(vertical_tile_17_15_to_tile_18_15_2),
		.in_wire_3_3(vertical_tile_17_15_to_tile_18_15_3),
		.out_wire_1_0(vertical_tile_18_15_to_tile_19_15_0),
		.out_wire_1_1(vertical_tile_18_15_to_tile_19_15_1),
		.out_wire_1_2(vertical_tile_18_15_to_tile_19_15_2),
		.out_wire_1_3(vertical_tile_18_15_to_tile_19_15_3),
		.in_wire_1_0(vertical_tile_19_15_to_tile_18_15_0),
		.in_wire_1_1(vertical_tile_19_15_to_tile_18_15_1),
		.in_wire_1_2(vertical_tile_19_15_to_tile_18_15_2),
		.in_wire_1_3(vertical_tile_19_15_to_tile_18_15_3),
		.out_wire_2_0(horizontal_tile_18_15_to_tile_18_14_0),
		.out_wire_2_1(horizontal_tile_18_15_to_tile_18_14_1),
		.out_wire_2_2(horizontal_tile_18_15_to_tile_18_14_2),
		.out_wire_2_3(horizontal_tile_18_15_to_tile_18_14_3),
		.in_wire_2_0(horizontal_tile_18_14_to_tile_18_15_0),
		.in_wire_2_1(horizontal_tile_18_14_to_tile_18_15_1),
		.in_wire_2_2(horizontal_tile_18_14_to_tile_18_15_2),
		.in_wire_2_3(horizontal_tile_18_14_to_tile_18_15_3),
		.out_wire_0_0(horizontal_tile_18_15_to_tile_18_16_0),
		.out_wire_0_1(horizontal_tile_18_15_to_tile_18_16_1),
		.out_wire_0_2(horizontal_tile_18_15_to_tile_18_16_2),
		.out_wire_0_3(horizontal_tile_18_15_to_tile_18_16_3),
		.in_wire_0_0(horizontal_tile_18_16_to_tile_18_15_0),
		.in_wire_0_1(horizontal_tile_18_16_to_tile_18_15_1),
		.in_wire_0_2(horizontal_tile_18_16_to_tile_18_15_2),
		.in_wire_0_3(horizontal_tile_18_16_to_tile_18_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(592)
	);

	pe_tile pe_tile_18_16(
		.out_wire_3_0(vertical_tile_18_16_to_tile_17_16_0),
		.out_wire_3_1(vertical_tile_18_16_to_tile_17_16_1),
		.out_wire_3_2(vertical_tile_18_16_to_tile_17_16_2),
		.out_wire_3_3(vertical_tile_18_16_to_tile_17_16_3),
		.in_wire_3_0(vertical_tile_17_16_to_tile_18_16_0),
		.in_wire_3_1(vertical_tile_17_16_to_tile_18_16_1),
		.in_wire_3_2(vertical_tile_17_16_to_tile_18_16_2),
		.in_wire_3_3(vertical_tile_17_16_to_tile_18_16_3),
		.out_wire_1_0(vertical_tile_18_16_to_tile_19_16_0),
		.out_wire_1_1(vertical_tile_18_16_to_tile_19_16_1),
		.out_wire_1_2(vertical_tile_18_16_to_tile_19_16_2),
		.out_wire_1_3(vertical_tile_18_16_to_tile_19_16_3),
		.in_wire_1_0(vertical_tile_19_16_to_tile_18_16_0),
		.in_wire_1_1(vertical_tile_19_16_to_tile_18_16_1),
		.in_wire_1_2(vertical_tile_19_16_to_tile_18_16_2),
		.in_wire_1_3(vertical_tile_19_16_to_tile_18_16_3),
		.out_wire_2_0(horizontal_tile_18_16_to_tile_18_15_0),
		.out_wire_2_1(horizontal_tile_18_16_to_tile_18_15_1),
		.out_wire_2_2(horizontal_tile_18_16_to_tile_18_15_2),
		.out_wire_2_3(horizontal_tile_18_16_to_tile_18_15_3),
		.in_wire_2_0(horizontal_tile_18_15_to_tile_18_16_0),
		.in_wire_2_1(horizontal_tile_18_15_to_tile_18_16_1),
		.in_wire_2_2(horizontal_tile_18_15_to_tile_18_16_2),
		.in_wire_2_3(horizontal_tile_18_15_to_tile_18_16_3),
		.out_wire_0_0(horizontal_tile_18_16_to_tile_18_17_0),
		.out_wire_0_1(horizontal_tile_18_16_to_tile_18_17_1),
		.out_wire_0_2(horizontal_tile_18_16_to_tile_18_17_2),
		.out_wire_0_3(horizontal_tile_18_16_to_tile_18_17_3),
		.in_wire_0_0(horizontal_tile_18_17_to_tile_18_16_0),
		.in_wire_0_1(horizontal_tile_18_17_to_tile_18_16_1),
		.in_wire_0_2(horizontal_tile_18_17_to_tile_18_16_2),
		.in_wire_0_3(horizontal_tile_18_17_to_tile_18_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(593)
	);

	pe_tile pe_tile_18_17(
		.out_wire_3_0(vertical_tile_18_17_to_tile_17_17_0),
		.out_wire_3_1(vertical_tile_18_17_to_tile_17_17_1),
		.out_wire_3_2(vertical_tile_18_17_to_tile_17_17_2),
		.out_wire_3_3(vertical_tile_18_17_to_tile_17_17_3),
		.in_wire_3_0(vertical_tile_17_17_to_tile_18_17_0),
		.in_wire_3_1(vertical_tile_17_17_to_tile_18_17_1),
		.in_wire_3_2(vertical_tile_17_17_to_tile_18_17_2),
		.in_wire_3_3(vertical_tile_17_17_to_tile_18_17_3),
		.out_wire_1_0(vertical_tile_18_17_to_tile_19_17_0),
		.out_wire_1_1(vertical_tile_18_17_to_tile_19_17_1),
		.out_wire_1_2(vertical_tile_18_17_to_tile_19_17_2),
		.out_wire_1_3(vertical_tile_18_17_to_tile_19_17_3),
		.in_wire_1_0(vertical_tile_19_17_to_tile_18_17_0),
		.in_wire_1_1(vertical_tile_19_17_to_tile_18_17_1),
		.in_wire_1_2(vertical_tile_19_17_to_tile_18_17_2),
		.in_wire_1_3(vertical_tile_19_17_to_tile_18_17_3),
		.out_wire_2_0(horizontal_tile_18_17_to_tile_18_16_0),
		.out_wire_2_1(horizontal_tile_18_17_to_tile_18_16_1),
		.out_wire_2_2(horizontal_tile_18_17_to_tile_18_16_2),
		.out_wire_2_3(horizontal_tile_18_17_to_tile_18_16_3),
		.in_wire_2_0(horizontal_tile_18_16_to_tile_18_17_0),
		.in_wire_2_1(horizontal_tile_18_16_to_tile_18_17_1),
		.in_wire_2_2(horizontal_tile_18_16_to_tile_18_17_2),
		.in_wire_2_3(horizontal_tile_18_16_to_tile_18_17_3),
		.out_wire_0_0(horizontal_tile_18_17_to_tile_18_18_0),
		.out_wire_0_1(horizontal_tile_18_17_to_tile_18_18_1),
		.out_wire_0_2(horizontal_tile_18_17_to_tile_18_18_2),
		.out_wire_0_3(horizontal_tile_18_17_to_tile_18_18_3),
		.in_wire_0_0(horizontal_tile_18_18_to_tile_18_17_0),
		.in_wire_0_1(horizontal_tile_18_18_to_tile_18_17_1),
		.in_wire_0_2(horizontal_tile_18_18_to_tile_18_17_2),
		.in_wire_0_3(horizontal_tile_18_18_to_tile_18_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(594)
	);

	pe_tile pe_tile_18_18(
		.out_wire_3_0(vertical_tile_18_18_to_tile_17_18_0),
		.out_wire_3_1(vertical_tile_18_18_to_tile_17_18_1),
		.out_wire_3_2(vertical_tile_18_18_to_tile_17_18_2),
		.out_wire_3_3(vertical_tile_18_18_to_tile_17_18_3),
		.in_wire_3_0(vertical_tile_17_18_to_tile_18_18_0),
		.in_wire_3_1(vertical_tile_17_18_to_tile_18_18_1),
		.in_wire_3_2(vertical_tile_17_18_to_tile_18_18_2),
		.in_wire_3_3(vertical_tile_17_18_to_tile_18_18_3),
		.out_wire_1_0(vertical_tile_18_18_to_tile_19_18_0),
		.out_wire_1_1(vertical_tile_18_18_to_tile_19_18_1),
		.out_wire_1_2(vertical_tile_18_18_to_tile_19_18_2),
		.out_wire_1_3(vertical_tile_18_18_to_tile_19_18_3),
		.in_wire_1_0(vertical_tile_19_18_to_tile_18_18_0),
		.in_wire_1_1(vertical_tile_19_18_to_tile_18_18_1),
		.in_wire_1_2(vertical_tile_19_18_to_tile_18_18_2),
		.in_wire_1_3(vertical_tile_19_18_to_tile_18_18_3),
		.out_wire_2_0(horizontal_tile_18_18_to_tile_18_17_0),
		.out_wire_2_1(horizontal_tile_18_18_to_tile_18_17_1),
		.out_wire_2_2(horizontal_tile_18_18_to_tile_18_17_2),
		.out_wire_2_3(horizontal_tile_18_18_to_tile_18_17_3),
		.in_wire_2_0(horizontal_tile_18_17_to_tile_18_18_0),
		.in_wire_2_1(horizontal_tile_18_17_to_tile_18_18_1),
		.in_wire_2_2(horizontal_tile_18_17_to_tile_18_18_2),
		.in_wire_2_3(horizontal_tile_18_17_to_tile_18_18_3),
		.out_wire_0_0(horizontal_tile_18_18_to_tile_18_19_0),
		.out_wire_0_1(horizontal_tile_18_18_to_tile_18_19_1),
		.out_wire_0_2(horizontal_tile_18_18_to_tile_18_19_2),
		.out_wire_0_3(horizontal_tile_18_18_to_tile_18_19_3),
		.in_wire_0_0(horizontal_tile_18_19_to_tile_18_18_0),
		.in_wire_0_1(horizontal_tile_18_19_to_tile_18_18_1),
		.in_wire_0_2(horizontal_tile_18_19_to_tile_18_18_2),
		.in_wire_0_3(horizontal_tile_18_19_to_tile_18_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(595)
	);

	pe_tile pe_tile_18_19(
		.out_wire_3_0(vertical_tile_18_19_to_tile_17_19_0),
		.out_wire_3_1(vertical_tile_18_19_to_tile_17_19_1),
		.out_wire_3_2(vertical_tile_18_19_to_tile_17_19_2),
		.out_wire_3_3(vertical_tile_18_19_to_tile_17_19_3),
		.in_wire_3_0(vertical_tile_17_19_to_tile_18_19_0),
		.in_wire_3_1(vertical_tile_17_19_to_tile_18_19_1),
		.in_wire_3_2(vertical_tile_17_19_to_tile_18_19_2),
		.in_wire_3_3(vertical_tile_17_19_to_tile_18_19_3),
		.out_wire_1_0(vertical_tile_18_19_to_tile_19_19_0),
		.out_wire_1_1(vertical_tile_18_19_to_tile_19_19_1),
		.out_wire_1_2(vertical_tile_18_19_to_tile_19_19_2),
		.out_wire_1_3(vertical_tile_18_19_to_tile_19_19_3),
		.in_wire_1_0(vertical_tile_19_19_to_tile_18_19_0),
		.in_wire_1_1(vertical_tile_19_19_to_tile_18_19_1),
		.in_wire_1_2(vertical_tile_19_19_to_tile_18_19_2),
		.in_wire_1_3(vertical_tile_19_19_to_tile_18_19_3),
		.out_wire_2_0(horizontal_tile_18_19_to_tile_18_18_0),
		.out_wire_2_1(horizontal_tile_18_19_to_tile_18_18_1),
		.out_wire_2_2(horizontal_tile_18_19_to_tile_18_18_2),
		.out_wire_2_3(horizontal_tile_18_19_to_tile_18_18_3),
		.in_wire_2_0(horizontal_tile_18_18_to_tile_18_19_0),
		.in_wire_2_1(horizontal_tile_18_18_to_tile_18_19_1),
		.in_wire_2_2(horizontal_tile_18_18_to_tile_18_19_2),
		.in_wire_2_3(horizontal_tile_18_18_to_tile_18_19_3),
		.out_wire_0_0(horizontal_tile_18_19_to_tile_18_20_0),
		.out_wire_0_1(horizontal_tile_18_19_to_tile_18_20_1),
		.out_wire_0_2(horizontal_tile_18_19_to_tile_18_20_2),
		.out_wire_0_3(horizontal_tile_18_19_to_tile_18_20_3),
		.in_wire_0_0(horizontal_tile_18_20_to_tile_18_19_0),
		.in_wire_0_1(horizontal_tile_18_20_to_tile_18_19_1),
		.in_wire_0_2(horizontal_tile_18_20_to_tile_18_19_2),
		.in_wire_0_3(horizontal_tile_18_20_to_tile_18_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(596)
	);

	pe_tile pe_tile_18_20(
		.out_wire_3_0(vertical_tile_18_20_to_tile_17_20_0),
		.out_wire_3_1(vertical_tile_18_20_to_tile_17_20_1),
		.out_wire_3_2(vertical_tile_18_20_to_tile_17_20_2),
		.out_wire_3_3(vertical_tile_18_20_to_tile_17_20_3),
		.in_wire_3_0(vertical_tile_17_20_to_tile_18_20_0),
		.in_wire_3_1(vertical_tile_17_20_to_tile_18_20_1),
		.in_wire_3_2(vertical_tile_17_20_to_tile_18_20_2),
		.in_wire_3_3(vertical_tile_17_20_to_tile_18_20_3),
		.out_wire_1_0(vertical_tile_18_20_to_tile_19_20_0),
		.out_wire_1_1(vertical_tile_18_20_to_tile_19_20_1),
		.out_wire_1_2(vertical_tile_18_20_to_tile_19_20_2),
		.out_wire_1_3(vertical_tile_18_20_to_tile_19_20_3),
		.in_wire_1_0(vertical_tile_19_20_to_tile_18_20_0),
		.in_wire_1_1(vertical_tile_19_20_to_tile_18_20_1),
		.in_wire_1_2(vertical_tile_19_20_to_tile_18_20_2),
		.in_wire_1_3(vertical_tile_19_20_to_tile_18_20_3),
		.out_wire_2_0(horizontal_tile_18_20_to_tile_18_19_0),
		.out_wire_2_1(horizontal_tile_18_20_to_tile_18_19_1),
		.out_wire_2_2(horizontal_tile_18_20_to_tile_18_19_2),
		.out_wire_2_3(horizontal_tile_18_20_to_tile_18_19_3),
		.in_wire_2_0(horizontal_tile_18_19_to_tile_18_20_0),
		.in_wire_2_1(horizontal_tile_18_19_to_tile_18_20_1),
		.in_wire_2_2(horizontal_tile_18_19_to_tile_18_20_2),
		.in_wire_2_3(horizontal_tile_18_19_to_tile_18_20_3),
		.out_wire_0_0(horizontal_tile_18_20_to_tile_18_21_0),
		.out_wire_0_1(horizontal_tile_18_20_to_tile_18_21_1),
		.out_wire_0_2(horizontal_tile_18_20_to_tile_18_21_2),
		.out_wire_0_3(horizontal_tile_18_20_to_tile_18_21_3),
		.in_wire_0_0(horizontal_tile_18_21_to_tile_18_20_0),
		.in_wire_0_1(horizontal_tile_18_21_to_tile_18_20_1),
		.in_wire_0_2(horizontal_tile_18_21_to_tile_18_20_2),
		.in_wire_0_3(horizontal_tile_18_21_to_tile_18_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(597)
	);

	pe_tile pe_tile_18_21(
		.out_wire_3_0(vertical_tile_18_21_to_tile_17_21_0),
		.out_wire_3_1(vertical_tile_18_21_to_tile_17_21_1),
		.out_wire_3_2(vertical_tile_18_21_to_tile_17_21_2),
		.out_wire_3_3(vertical_tile_18_21_to_tile_17_21_3),
		.in_wire_3_0(vertical_tile_17_21_to_tile_18_21_0),
		.in_wire_3_1(vertical_tile_17_21_to_tile_18_21_1),
		.in_wire_3_2(vertical_tile_17_21_to_tile_18_21_2),
		.in_wire_3_3(vertical_tile_17_21_to_tile_18_21_3),
		.out_wire_1_0(vertical_tile_18_21_to_tile_19_21_0),
		.out_wire_1_1(vertical_tile_18_21_to_tile_19_21_1),
		.out_wire_1_2(vertical_tile_18_21_to_tile_19_21_2),
		.out_wire_1_3(vertical_tile_18_21_to_tile_19_21_3),
		.in_wire_1_0(vertical_tile_19_21_to_tile_18_21_0),
		.in_wire_1_1(vertical_tile_19_21_to_tile_18_21_1),
		.in_wire_1_2(vertical_tile_19_21_to_tile_18_21_2),
		.in_wire_1_3(vertical_tile_19_21_to_tile_18_21_3),
		.out_wire_2_0(horizontal_tile_18_21_to_tile_18_20_0),
		.out_wire_2_1(horizontal_tile_18_21_to_tile_18_20_1),
		.out_wire_2_2(horizontal_tile_18_21_to_tile_18_20_2),
		.out_wire_2_3(horizontal_tile_18_21_to_tile_18_20_3),
		.in_wire_2_0(horizontal_tile_18_20_to_tile_18_21_0),
		.in_wire_2_1(horizontal_tile_18_20_to_tile_18_21_1),
		.in_wire_2_2(horizontal_tile_18_20_to_tile_18_21_2),
		.in_wire_2_3(horizontal_tile_18_20_to_tile_18_21_3),
		.out_wire_0_0(horizontal_tile_18_21_to_tile_18_22_0),
		.out_wire_0_1(horizontal_tile_18_21_to_tile_18_22_1),
		.out_wire_0_2(horizontal_tile_18_21_to_tile_18_22_2),
		.out_wire_0_3(horizontal_tile_18_21_to_tile_18_22_3),
		.in_wire_0_0(horizontal_tile_18_22_to_tile_18_21_0),
		.in_wire_0_1(horizontal_tile_18_22_to_tile_18_21_1),
		.in_wire_0_2(horizontal_tile_18_22_to_tile_18_21_2),
		.in_wire_0_3(horizontal_tile_18_22_to_tile_18_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(598)
	);

	pe_tile pe_tile_18_22(
		.out_wire_3_0(vertical_tile_18_22_to_tile_17_22_0),
		.out_wire_3_1(vertical_tile_18_22_to_tile_17_22_1),
		.out_wire_3_2(vertical_tile_18_22_to_tile_17_22_2),
		.out_wire_3_3(vertical_tile_18_22_to_tile_17_22_3),
		.in_wire_3_0(vertical_tile_17_22_to_tile_18_22_0),
		.in_wire_3_1(vertical_tile_17_22_to_tile_18_22_1),
		.in_wire_3_2(vertical_tile_17_22_to_tile_18_22_2),
		.in_wire_3_3(vertical_tile_17_22_to_tile_18_22_3),
		.out_wire_1_0(vertical_tile_18_22_to_tile_19_22_0),
		.out_wire_1_1(vertical_tile_18_22_to_tile_19_22_1),
		.out_wire_1_2(vertical_tile_18_22_to_tile_19_22_2),
		.out_wire_1_3(vertical_tile_18_22_to_tile_19_22_3),
		.in_wire_1_0(vertical_tile_19_22_to_tile_18_22_0),
		.in_wire_1_1(vertical_tile_19_22_to_tile_18_22_1),
		.in_wire_1_2(vertical_tile_19_22_to_tile_18_22_2),
		.in_wire_1_3(vertical_tile_19_22_to_tile_18_22_3),
		.out_wire_2_0(horizontal_tile_18_22_to_tile_18_21_0),
		.out_wire_2_1(horizontal_tile_18_22_to_tile_18_21_1),
		.out_wire_2_2(horizontal_tile_18_22_to_tile_18_21_2),
		.out_wire_2_3(horizontal_tile_18_22_to_tile_18_21_3),
		.in_wire_2_0(horizontal_tile_18_21_to_tile_18_22_0),
		.in_wire_2_1(horizontal_tile_18_21_to_tile_18_22_1),
		.in_wire_2_2(horizontal_tile_18_21_to_tile_18_22_2),
		.in_wire_2_3(horizontal_tile_18_21_to_tile_18_22_3),
		.out_wire_0_0(horizontal_tile_18_22_to_tile_18_23_0),
		.out_wire_0_1(horizontal_tile_18_22_to_tile_18_23_1),
		.out_wire_0_2(horizontal_tile_18_22_to_tile_18_23_2),
		.out_wire_0_3(horizontal_tile_18_22_to_tile_18_23_3),
		.in_wire_0_0(horizontal_tile_18_23_to_tile_18_22_0),
		.in_wire_0_1(horizontal_tile_18_23_to_tile_18_22_1),
		.in_wire_0_2(horizontal_tile_18_23_to_tile_18_22_2),
		.in_wire_0_3(horizontal_tile_18_23_to_tile_18_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(599)
	);

	pe_tile pe_tile_18_23(
		.out_wire_3_0(vertical_tile_18_23_to_tile_17_23_0),
		.out_wire_3_1(vertical_tile_18_23_to_tile_17_23_1),
		.out_wire_3_2(vertical_tile_18_23_to_tile_17_23_2),
		.out_wire_3_3(vertical_tile_18_23_to_tile_17_23_3),
		.in_wire_3_0(vertical_tile_17_23_to_tile_18_23_0),
		.in_wire_3_1(vertical_tile_17_23_to_tile_18_23_1),
		.in_wire_3_2(vertical_tile_17_23_to_tile_18_23_2),
		.in_wire_3_3(vertical_tile_17_23_to_tile_18_23_3),
		.out_wire_1_0(vertical_tile_18_23_to_tile_19_23_0),
		.out_wire_1_1(vertical_tile_18_23_to_tile_19_23_1),
		.out_wire_1_2(vertical_tile_18_23_to_tile_19_23_2),
		.out_wire_1_3(vertical_tile_18_23_to_tile_19_23_3),
		.in_wire_1_0(vertical_tile_19_23_to_tile_18_23_0),
		.in_wire_1_1(vertical_tile_19_23_to_tile_18_23_1),
		.in_wire_1_2(vertical_tile_19_23_to_tile_18_23_2),
		.in_wire_1_3(vertical_tile_19_23_to_tile_18_23_3),
		.out_wire_2_0(horizontal_tile_18_23_to_tile_18_22_0),
		.out_wire_2_1(horizontal_tile_18_23_to_tile_18_22_1),
		.out_wire_2_2(horizontal_tile_18_23_to_tile_18_22_2),
		.out_wire_2_3(horizontal_tile_18_23_to_tile_18_22_3),
		.in_wire_2_0(horizontal_tile_18_22_to_tile_18_23_0),
		.in_wire_2_1(horizontal_tile_18_22_to_tile_18_23_1),
		.in_wire_2_2(horizontal_tile_18_22_to_tile_18_23_2),
		.in_wire_2_3(horizontal_tile_18_22_to_tile_18_23_3),
		.out_wire_0_0(horizontal_tile_18_23_to_tile_18_24_0),
		.out_wire_0_1(horizontal_tile_18_23_to_tile_18_24_1),
		.out_wire_0_2(horizontal_tile_18_23_to_tile_18_24_2),
		.out_wire_0_3(horizontal_tile_18_23_to_tile_18_24_3),
		.in_wire_0_0(horizontal_tile_18_24_to_tile_18_23_0),
		.in_wire_0_1(horizontal_tile_18_24_to_tile_18_23_1),
		.in_wire_0_2(horizontal_tile_18_24_to_tile_18_23_2),
		.in_wire_0_3(horizontal_tile_18_24_to_tile_18_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(600)
	);

	pe_tile pe_tile_18_24(
		.out_wire_3_0(vertical_tile_18_24_to_tile_17_24_0),
		.out_wire_3_1(vertical_tile_18_24_to_tile_17_24_1),
		.out_wire_3_2(vertical_tile_18_24_to_tile_17_24_2),
		.out_wire_3_3(vertical_tile_18_24_to_tile_17_24_3),
		.in_wire_3_0(vertical_tile_17_24_to_tile_18_24_0),
		.in_wire_3_1(vertical_tile_17_24_to_tile_18_24_1),
		.in_wire_3_2(vertical_tile_17_24_to_tile_18_24_2),
		.in_wire_3_3(vertical_tile_17_24_to_tile_18_24_3),
		.out_wire_1_0(vertical_tile_18_24_to_tile_19_24_0),
		.out_wire_1_1(vertical_tile_18_24_to_tile_19_24_1),
		.out_wire_1_2(vertical_tile_18_24_to_tile_19_24_2),
		.out_wire_1_3(vertical_tile_18_24_to_tile_19_24_3),
		.in_wire_1_0(vertical_tile_19_24_to_tile_18_24_0),
		.in_wire_1_1(vertical_tile_19_24_to_tile_18_24_1),
		.in_wire_1_2(vertical_tile_19_24_to_tile_18_24_2),
		.in_wire_1_3(vertical_tile_19_24_to_tile_18_24_3),
		.out_wire_2_0(horizontal_tile_18_24_to_tile_18_23_0),
		.out_wire_2_1(horizontal_tile_18_24_to_tile_18_23_1),
		.out_wire_2_2(horizontal_tile_18_24_to_tile_18_23_2),
		.out_wire_2_3(horizontal_tile_18_24_to_tile_18_23_3),
		.in_wire_2_0(horizontal_tile_18_23_to_tile_18_24_0),
		.in_wire_2_1(horizontal_tile_18_23_to_tile_18_24_1),
		.in_wire_2_2(horizontal_tile_18_23_to_tile_18_24_2),
		.in_wire_2_3(horizontal_tile_18_23_to_tile_18_24_3),
		.out_wire_0_0(horizontal_tile_18_24_to_tile_18_25_0),
		.out_wire_0_1(horizontal_tile_18_24_to_tile_18_25_1),
		.out_wire_0_2(horizontal_tile_18_24_to_tile_18_25_2),
		.out_wire_0_3(horizontal_tile_18_24_to_tile_18_25_3),
		.in_wire_0_0(horizontal_tile_18_25_to_tile_18_24_0),
		.in_wire_0_1(horizontal_tile_18_25_to_tile_18_24_1),
		.in_wire_0_2(horizontal_tile_18_25_to_tile_18_24_2),
		.in_wire_0_3(horizontal_tile_18_25_to_tile_18_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(601)
	);

	pe_tile pe_tile_18_25(
		.out_wire_3_0(vertical_tile_18_25_to_tile_17_25_0),
		.out_wire_3_1(vertical_tile_18_25_to_tile_17_25_1),
		.out_wire_3_2(vertical_tile_18_25_to_tile_17_25_2),
		.out_wire_3_3(vertical_tile_18_25_to_tile_17_25_3),
		.in_wire_3_0(vertical_tile_17_25_to_tile_18_25_0),
		.in_wire_3_1(vertical_tile_17_25_to_tile_18_25_1),
		.in_wire_3_2(vertical_tile_17_25_to_tile_18_25_2),
		.in_wire_3_3(vertical_tile_17_25_to_tile_18_25_3),
		.out_wire_1_0(vertical_tile_18_25_to_tile_19_25_0),
		.out_wire_1_1(vertical_tile_18_25_to_tile_19_25_1),
		.out_wire_1_2(vertical_tile_18_25_to_tile_19_25_2),
		.out_wire_1_3(vertical_tile_18_25_to_tile_19_25_3),
		.in_wire_1_0(vertical_tile_19_25_to_tile_18_25_0),
		.in_wire_1_1(vertical_tile_19_25_to_tile_18_25_1),
		.in_wire_1_2(vertical_tile_19_25_to_tile_18_25_2),
		.in_wire_1_3(vertical_tile_19_25_to_tile_18_25_3),
		.out_wire_2_0(horizontal_tile_18_25_to_tile_18_24_0),
		.out_wire_2_1(horizontal_tile_18_25_to_tile_18_24_1),
		.out_wire_2_2(horizontal_tile_18_25_to_tile_18_24_2),
		.out_wire_2_3(horizontal_tile_18_25_to_tile_18_24_3),
		.in_wire_2_0(horizontal_tile_18_24_to_tile_18_25_0),
		.in_wire_2_1(horizontal_tile_18_24_to_tile_18_25_1),
		.in_wire_2_2(horizontal_tile_18_24_to_tile_18_25_2),
		.in_wire_2_3(horizontal_tile_18_24_to_tile_18_25_3),
		.out_wire_0_0(horizontal_tile_18_25_to_tile_18_26_0),
		.out_wire_0_1(horizontal_tile_18_25_to_tile_18_26_1),
		.out_wire_0_2(horizontal_tile_18_25_to_tile_18_26_2),
		.out_wire_0_3(horizontal_tile_18_25_to_tile_18_26_3),
		.in_wire_0_0(horizontal_tile_18_26_to_tile_18_25_0),
		.in_wire_0_1(horizontal_tile_18_26_to_tile_18_25_1),
		.in_wire_0_2(horizontal_tile_18_26_to_tile_18_25_2),
		.in_wire_0_3(horizontal_tile_18_26_to_tile_18_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(602)
	);

	pe_tile pe_tile_18_26(
		.out_wire_3_0(vertical_tile_18_26_to_tile_17_26_0),
		.out_wire_3_1(vertical_tile_18_26_to_tile_17_26_1),
		.out_wire_3_2(vertical_tile_18_26_to_tile_17_26_2),
		.out_wire_3_3(vertical_tile_18_26_to_tile_17_26_3),
		.in_wire_3_0(vertical_tile_17_26_to_tile_18_26_0),
		.in_wire_3_1(vertical_tile_17_26_to_tile_18_26_1),
		.in_wire_3_2(vertical_tile_17_26_to_tile_18_26_2),
		.in_wire_3_3(vertical_tile_17_26_to_tile_18_26_3),
		.out_wire_1_0(vertical_tile_18_26_to_tile_19_26_0),
		.out_wire_1_1(vertical_tile_18_26_to_tile_19_26_1),
		.out_wire_1_2(vertical_tile_18_26_to_tile_19_26_2),
		.out_wire_1_3(vertical_tile_18_26_to_tile_19_26_3),
		.in_wire_1_0(vertical_tile_19_26_to_tile_18_26_0),
		.in_wire_1_1(vertical_tile_19_26_to_tile_18_26_1),
		.in_wire_1_2(vertical_tile_19_26_to_tile_18_26_2),
		.in_wire_1_3(vertical_tile_19_26_to_tile_18_26_3),
		.out_wire_2_0(horizontal_tile_18_26_to_tile_18_25_0),
		.out_wire_2_1(horizontal_tile_18_26_to_tile_18_25_1),
		.out_wire_2_2(horizontal_tile_18_26_to_tile_18_25_2),
		.out_wire_2_3(horizontal_tile_18_26_to_tile_18_25_3),
		.in_wire_2_0(horizontal_tile_18_25_to_tile_18_26_0),
		.in_wire_2_1(horizontal_tile_18_25_to_tile_18_26_1),
		.in_wire_2_2(horizontal_tile_18_25_to_tile_18_26_2),
		.in_wire_2_3(horizontal_tile_18_25_to_tile_18_26_3),
		.out_wire_0_0(horizontal_tile_18_26_to_tile_18_27_0),
		.out_wire_0_1(horizontal_tile_18_26_to_tile_18_27_1),
		.out_wire_0_2(horizontal_tile_18_26_to_tile_18_27_2),
		.out_wire_0_3(horizontal_tile_18_26_to_tile_18_27_3),
		.in_wire_0_0(horizontal_tile_18_27_to_tile_18_26_0),
		.in_wire_0_1(horizontal_tile_18_27_to_tile_18_26_1),
		.in_wire_0_2(horizontal_tile_18_27_to_tile_18_26_2),
		.in_wire_0_3(horizontal_tile_18_27_to_tile_18_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(603)
	);

	pe_tile pe_tile_18_27(
		.out_wire_3_0(vertical_tile_18_27_to_tile_17_27_0),
		.out_wire_3_1(vertical_tile_18_27_to_tile_17_27_1),
		.out_wire_3_2(vertical_tile_18_27_to_tile_17_27_2),
		.out_wire_3_3(vertical_tile_18_27_to_tile_17_27_3),
		.in_wire_3_0(vertical_tile_17_27_to_tile_18_27_0),
		.in_wire_3_1(vertical_tile_17_27_to_tile_18_27_1),
		.in_wire_3_2(vertical_tile_17_27_to_tile_18_27_2),
		.in_wire_3_3(vertical_tile_17_27_to_tile_18_27_3),
		.out_wire_1_0(vertical_tile_18_27_to_tile_19_27_0),
		.out_wire_1_1(vertical_tile_18_27_to_tile_19_27_1),
		.out_wire_1_2(vertical_tile_18_27_to_tile_19_27_2),
		.out_wire_1_3(vertical_tile_18_27_to_tile_19_27_3),
		.in_wire_1_0(vertical_tile_19_27_to_tile_18_27_0),
		.in_wire_1_1(vertical_tile_19_27_to_tile_18_27_1),
		.in_wire_1_2(vertical_tile_19_27_to_tile_18_27_2),
		.in_wire_1_3(vertical_tile_19_27_to_tile_18_27_3),
		.out_wire_2_0(horizontal_tile_18_27_to_tile_18_26_0),
		.out_wire_2_1(horizontal_tile_18_27_to_tile_18_26_1),
		.out_wire_2_2(horizontal_tile_18_27_to_tile_18_26_2),
		.out_wire_2_3(horizontal_tile_18_27_to_tile_18_26_3),
		.in_wire_2_0(horizontal_tile_18_26_to_tile_18_27_0),
		.in_wire_2_1(horizontal_tile_18_26_to_tile_18_27_1),
		.in_wire_2_2(horizontal_tile_18_26_to_tile_18_27_2),
		.in_wire_2_3(horizontal_tile_18_26_to_tile_18_27_3),
		.out_wire_0_0(horizontal_tile_18_27_to_tile_18_28_0),
		.out_wire_0_1(horizontal_tile_18_27_to_tile_18_28_1),
		.out_wire_0_2(horizontal_tile_18_27_to_tile_18_28_2),
		.out_wire_0_3(horizontal_tile_18_27_to_tile_18_28_3),
		.in_wire_0_0(horizontal_tile_18_28_to_tile_18_27_0),
		.in_wire_0_1(horizontal_tile_18_28_to_tile_18_27_1),
		.in_wire_0_2(horizontal_tile_18_28_to_tile_18_27_2),
		.in_wire_0_3(horizontal_tile_18_28_to_tile_18_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(604)
	);

	pe_tile pe_tile_18_28(
		.out_wire_3_0(vertical_tile_18_28_to_tile_17_28_0),
		.out_wire_3_1(vertical_tile_18_28_to_tile_17_28_1),
		.out_wire_3_2(vertical_tile_18_28_to_tile_17_28_2),
		.out_wire_3_3(vertical_tile_18_28_to_tile_17_28_3),
		.in_wire_3_0(vertical_tile_17_28_to_tile_18_28_0),
		.in_wire_3_1(vertical_tile_17_28_to_tile_18_28_1),
		.in_wire_3_2(vertical_tile_17_28_to_tile_18_28_2),
		.in_wire_3_3(vertical_tile_17_28_to_tile_18_28_3),
		.out_wire_1_0(vertical_tile_18_28_to_tile_19_28_0),
		.out_wire_1_1(vertical_tile_18_28_to_tile_19_28_1),
		.out_wire_1_2(vertical_tile_18_28_to_tile_19_28_2),
		.out_wire_1_3(vertical_tile_18_28_to_tile_19_28_3),
		.in_wire_1_0(vertical_tile_19_28_to_tile_18_28_0),
		.in_wire_1_1(vertical_tile_19_28_to_tile_18_28_1),
		.in_wire_1_2(vertical_tile_19_28_to_tile_18_28_2),
		.in_wire_1_3(vertical_tile_19_28_to_tile_18_28_3),
		.out_wire_2_0(horizontal_tile_18_28_to_tile_18_27_0),
		.out_wire_2_1(horizontal_tile_18_28_to_tile_18_27_1),
		.out_wire_2_2(horizontal_tile_18_28_to_tile_18_27_2),
		.out_wire_2_3(horizontal_tile_18_28_to_tile_18_27_3),
		.in_wire_2_0(horizontal_tile_18_27_to_tile_18_28_0),
		.in_wire_2_1(horizontal_tile_18_27_to_tile_18_28_1),
		.in_wire_2_2(horizontal_tile_18_27_to_tile_18_28_2),
		.in_wire_2_3(horizontal_tile_18_27_to_tile_18_28_3),
		.out_wire_0_0(horizontal_tile_18_28_to_tile_18_29_0),
		.out_wire_0_1(horizontal_tile_18_28_to_tile_18_29_1),
		.out_wire_0_2(horizontal_tile_18_28_to_tile_18_29_2),
		.out_wire_0_3(horizontal_tile_18_28_to_tile_18_29_3),
		.in_wire_0_0(horizontal_tile_18_29_to_tile_18_28_0),
		.in_wire_0_1(horizontal_tile_18_29_to_tile_18_28_1),
		.in_wire_0_2(horizontal_tile_18_29_to_tile_18_28_2),
		.in_wire_0_3(horizontal_tile_18_29_to_tile_18_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(605)
	);

	pe_tile pe_tile_18_29(
		.out_wire_3_0(vertical_tile_18_29_to_tile_17_29_0),
		.out_wire_3_1(vertical_tile_18_29_to_tile_17_29_1),
		.out_wire_3_2(vertical_tile_18_29_to_tile_17_29_2),
		.out_wire_3_3(vertical_tile_18_29_to_tile_17_29_3),
		.in_wire_3_0(vertical_tile_17_29_to_tile_18_29_0),
		.in_wire_3_1(vertical_tile_17_29_to_tile_18_29_1),
		.in_wire_3_2(vertical_tile_17_29_to_tile_18_29_2),
		.in_wire_3_3(vertical_tile_17_29_to_tile_18_29_3),
		.out_wire_1_0(vertical_tile_18_29_to_tile_19_29_0),
		.out_wire_1_1(vertical_tile_18_29_to_tile_19_29_1),
		.out_wire_1_2(vertical_tile_18_29_to_tile_19_29_2),
		.out_wire_1_3(vertical_tile_18_29_to_tile_19_29_3),
		.in_wire_1_0(vertical_tile_19_29_to_tile_18_29_0),
		.in_wire_1_1(vertical_tile_19_29_to_tile_18_29_1),
		.in_wire_1_2(vertical_tile_19_29_to_tile_18_29_2),
		.in_wire_1_3(vertical_tile_19_29_to_tile_18_29_3),
		.out_wire_2_0(horizontal_tile_18_29_to_tile_18_28_0),
		.out_wire_2_1(horizontal_tile_18_29_to_tile_18_28_1),
		.out_wire_2_2(horizontal_tile_18_29_to_tile_18_28_2),
		.out_wire_2_3(horizontal_tile_18_29_to_tile_18_28_3),
		.in_wire_2_0(horizontal_tile_18_28_to_tile_18_29_0),
		.in_wire_2_1(horizontal_tile_18_28_to_tile_18_29_1),
		.in_wire_2_2(horizontal_tile_18_28_to_tile_18_29_2),
		.in_wire_2_3(horizontal_tile_18_28_to_tile_18_29_3),
		.out_wire_0_0(horizontal_tile_18_29_to_tile_18_30_0),
		.out_wire_0_1(horizontal_tile_18_29_to_tile_18_30_1),
		.out_wire_0_2(horizontal_tile_18_29_to_tile_18_30_2),
		.out_wire_0_3(horizontal_tile_18_29_to_tile_18_30_3),
		.in_wire_0_0(horizontal_tile_18_30_to_tile_18_29_0),
		.in_wire_0_1(horizontal_tile_18_30_to_tile_18_29_1),
		.in_wire_0_2(horizontal_tile_18_30_to_tile_18_29_2),
		.in_wire_0_3(horizontal_tile_18_30_to_tile_18_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(606)
	);

	pe_tile pe_tile_18_30(
		.out_wire_3_0(vertical_tile_18_30_to_tile_17_30_0),
		.out_wire_3_1(vertical_tile_18_30_to_tile_17_30_1),
		.out_wire_3_2(vertical_tile_18_30_to_tile_17_30_2),
		.out_wire_3_3(vertical_tile_18_30_to_tile_17_30_3),
		.in_wire_3_0(vertical_tile_17_30_to_tile_18_30_0),
		.in_wire_3_1(vertical_tile_17_30_to_tile_18_30_1),
		.in_wire_3_2(vertical_tile_17_30_to_tile_18_30_2),
		.in_wire_3_3(vertical_tile_17_30_to_tile_18_30_3),
		.out_wire_1_0(vertical_tile_18_30_to_tile_19_30_0),
		.out_wire_1_1(vertical_tile_18_30_to_tile_19_30_1),
		.out_wire_1_2(vertical_tile_18_30_to_tile_19_30_2),
		.out_wire_1_3(vertical_tile_18_30_to_tile_19_30_3),
		.in_wire_1_0(vertical_tile_19_30_to_tile_18_30_0),
		.in_wire_1_1(vertical_tile_19_30_to_tile_18_30_1),
		.in_wire_1_2(vertical_tile_19_30_to_tile_18_30_2),
		.in_wire_1_3(vertical_tile_19_30_to_tile_18_30_3),
		.out_wire_2_0(horizontal_tile_18_30_to_tile_18_29_0),
		.out_wire_2_1(horizontal_tile_18_30_to_tile_18_29_1),
		.out_wire_2_2(horizontal_tile_18_30_to_tile_18_29_2),
		.out_wire_2_3(horizontal_tile_18_30_to_tile_18_29_3),
		.in_wire_2_0(horizontal_tile_18_29_to_tile_18_30_0),
		.in_wire_2_1(horizontal_tile_18_29_to_tile_18_30_1),
		.in_wire_2_2(horizontal_tile_18_29_to_tile_18_30_2),
		.in_wire_2_3(horizontal_tile_18_29_to_tile_18_30_3),
		.out_wire_0_0(horizontal_tile_18_30_to_tile_18_31_0),
		.out_wire_0_1(horizontal_tile_18_30_to_tile_18_31_1),
		.out_wire_0_2(horizontal_tile_18_30_to_tile_18_31_2),
		.out_wire_0_3(horizontal_tile_18_30_to_tile_18_31_3),
		.in_wire_0_0(horizontal_tile_18_31_to_tile_18_30_0),
		.in_wire_0_1(horizontal_tile_18_31_to_tile_18_30_1),
		.in_wire_0_2(horizontal_tile_18_31_to_tile_18_30_2),
		.in_wire_0_3(horizontal_tile_18_31_to_tile_18_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(607)
	);

	pe_tile_right pe_tile_18_31(
		.out_wire_3_0(vertical_tile_18_31_to_tile_17_31_0),
		.out_wire_3_1(vertical_tile_18_31_to_tile_17_31_1),
		.out_wire_3_2(vertical_tile_18_31_to_tile_17_31_2),
		.out_wire_3_3(vertical_tile_18_31_to_tile_17_31_3),
		.in_wire_3_0(vertical_tile_17_31_to_tile_18_31_0),
		.in_wire_3_1(vertical_tile_17_31_to_tile_18_31_1),
		.in_wire_3_2(vertical_tile_17_31_to_tile_18_31_2),
		.in_wire_3_3(vertical_tile_17_31_to_tile_18_31_3),
		.out_wire_1_0(vertical_tile_18_31_to_tile_19_31_0),
		.out_wire_1_1(vertical_tile_18_31_to_tile_19_31_1),
		.out_wire_1_2(vertical_tile_18_31_to_tile_19_31_2),
		.out_wire_1_3(vertical_tile_18_31_to_tile_19_31_3),
		.in_wire_1_0(vertical_tile_19_31_to_tile_18_31_0),
		.in_wire_1_1(vertical_tile_19_31_to_tile_18_31_1),
		.in_wire_1_2(vertical_tile_19_31_to_tile_18_31_2),
		.in_wire_1_3(vertical_tile_19_31_to_tile_18_31_3),
		.out_wire_2_0(horizontal_tile_18_31_to_tile_18_30_0),
		.out_wire_2_1(horizontal_tile_18_31_to_tile_18_30_1),
		.out_wire_2_2(horizontal_tile_18_31_to_tile_18_30_2),
		.out_wire_2_3(horizontal_tile_18_31_to_tile_18_30_3),
		.in_wire_2_0(horizontal_tile_18_30_to_tile_18_31_0),
		.in_wire_2_1(horizontal_tile_18_30_to_tile_18_31_1),
		.in_wire_2_2(horizontal_tile_18_30_to_tile_18_31_2),
		.in_wire_2_3(horizontal_tile_18_30_to_tile_18_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(608)
	);

	pe_tile_left pe_tile_19_0(
		.out_wire_3_0(vertical_tile_19_0_to_tile_18_0_0),
		.out_wire_3_1(vertical_tile_19_0_to_tile_18_0_1),
		.out_wire_3_2(vertical_tile_19_0_to_tile_18_0_2),
		.out_wire_3_3(vertical_tile_19_0_to_tile_18_0_3),
		.in_wire_3_0(vertical_tile_18_0_to_tile_19_0_0),
		.in_wire_3_1(vertical_tile_18_0_to_tile_19_0_1),
		.in_wire_3_2(vertical_tile_18_0_to_tile_19_0_2),
		.in_wire_3_3(vertical_tile_18_0_to_tile_19_0_3),
		.out_wire_1_0(vertical_tile_19_0_to_tile_20_0_0),
		.out_wire_1_1(vertical_tile_19_0_to_tile_20_0_1),
		.out_wire_1_2(vertical_tile_19_0_to_tile_20_0_2),
		.out_wire_1_3(vertical_tile_19_0_to_tile_20_0_3),
		.in_wire_1_0(vertical_tile_20_0_to_tile_19_0_0),
		.in_wire_1_1(vertical_tile_20_0_to_tile_19_0_1),
		.in_wire_1_2(vertical_tile_20_0_to_tile_19_0_2),
		.in_wire_1_3(vertical_tile_20_0_to_tile_19_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_19_0_to_tile_19_1_0),
		.out_wire_0_1(horizontal_tile_19_0_to_tile_19_1_1),
		.out_wire_0_2(horizontal_tile_19_0_to_tile_19_1_2),
		.out_wire_0_3(horizontal_tile_19_0_to_tile_19_1_3),
		.in_wire_0_0(horizontal_tile_19_1_to_tile_19_0_0),
		.in_wire_0_1(horizontal_tile_19_1_to_tile_19_0_1),
		.in_wire_0_2(horizontal_tile_19_1_to_tile_19_0_2),
		.in_wire_0_3(horizontal_tile_19_1_to_tile_19_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(609)
	);

	pe_tile pe_tile_19_1(
		.out_wire_3_0(vertical_tile_19_1_to_tile_18_1_0),
		.out_wire_3_1(vertical_tile_19_1_to_tile_18_1_1),
		.out_wire_3_2(vertical_tile_19_1_to_tile_18_1_2),
		.out_wire_3_3(vertical_tile_19_1_to_tile_18_1_3),
		.in_wire_3_0(vertical_tile_18_1_to_tile_19_1_0),
		.in_wire_3_1(vertical_tile_18_1_to_tile_19_1_1),
		.in_wire_3_2(vertical_tile_18_1_to_tile_19_1_2),
		.in_wire_3_3(vertical_tile_18_1_to_tile_19_1_3),
		.out_wire_1_0(vertical_tile_19_1_to_tile_20_1_0),
		.out_wire_1_1(vertical_tile_19_1_to_tile_20_1_1),
		.out_wire_1_2(vertical_tile_19_1_to_tile_20_1_2),
		.out_wire_1_3(vertical_tile_19_1_to_tile_20_1_3),
		.in_wire_1_0(vertical_tile_20_1_to_tile_19_1_0),
		.in_wire_1_1(vertical_tile_20_1_to_tile_19_1_1),
		.in_wire_1_2(vertical_tile_20_1_to_tile_19_1_2),
		.in_wire_1_3(vertical_tile_20_1_to_tile_19_1_3),
		.out_wire_2_0(horizontal_tile_19_1_to_tile_19_0_0),
		.out_wire_2_1(horizontal_tile_19_1_to_tile_19_0_1),
		.out_wire_2_2(horizontal_tile_19_1_to_tile_19_0_2),
		.out_wire_2_3(horizontal_tile_19_1_to_tile_19_0_3),
		.in_wire_2_0(horizontal_tile_19_0_to_tile_19_1_0),
		.in_wire_2_1(horizontal_tile_19_0_to_tile_19_1_1),
		.in_wire_2_2(horizontal_tile_19_0_to_tile_19_1_2),
		.in_wire_2_3(horizontal_tile_19_0_to_tile_19_1_3),
		.out_wire_0_0(horizontal_tile_19_1_to_tile_19_2_0),
		.out_wire_0_1(horizontal_tile_19_1_to_tile_19_2_1),
		.out_wire_0_2(horizontal_tile_19_1_to_tile_19_2_2),
		.out_wire_0_3(horizontal_tile_19_1_to_tile_19_2_3),
		.in_wire_0_0(horizontal_tile_19_2_to_tile_19_1_0),
		.in_wire_0_1(horizontal_tile_19_2_to_tile_19_1_1),
		.in_wire_0_2(horizontal_tile_19_2_to_tile_19_1_2),
		.in_wire_0_3(horizontal_tile_19_2_to_tile_19_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(610)
	);

	pe_tile pe_tile_19_2(
		.out_wire_3_0(vertical_tile_19_2_to_tile_18_2_0),
		.out_wire_3_1(vertical_tile_19_2_to_tile_18_2_1),
		.out_wire_3_2(vertical_tile_19_2_to_tile_18_2_2),
		.out_wire_3_3(vertical_tile_19_2_to_tile_18_2_3),
		.in_wire_3_0(vertical_tile_18_2_to_tile_19_2_0),
		.in_wire_3_1(vertical_tile_18_2_to_tile_19_2_1),
		.in_wire_3_2(vertical_tile_18_2_to_tile_19_2_2),
		.in_wire_3_3(vertical_tile_18_2_to_tile_19_2_3),
		.out_wire_1_0(vertical_tile_19_2_to_tile_20_2_0),
		.out_wire_1_1(vertical_tile_19_2_to_tile_20_2_1),
		.out_wire_1_2(vertical_tile_19_2_to_tile_20_2_2),
		.out_wire_1_3(vertical_tile_19_2_to_tile_20_2_3),
		.in_wire_1_0(vertical_tile_20_2_to_tile_19_2_0),
		.in_wire_1_1(vertical_tile_20_2_to_tile_19_2_1),
		.in_wire_1_2(vertical_tile_20_2_to_tile_19_2_2),
		.in_wire_1_3(vertical_tile_20_2_to_tile_19_2_3),
		.out_wire_2_0(horizontal_tile_19_2_to_tile_19_1_0),
		.out_wire_2_1(horizontal_tile_19_2_to_tile_19_1_1),
		.out_wire_2_2(horizontal_tile_19_2_to_tile_19_1_2),
		.out_wire_2_3(horizontal_tile_19_2_to_tile_19_1_3),
		.in_wire_2_0(horizontal_tile_19_1_to_tile_19_2_0),
		.in_wire_2_1(horizontal_tile_19_1_to_tile_19_2_1),
		.in_wire_2_2(horizontal_tile_19_1_to_tile_19_2_2),
		.in_wire_2_3(horizontal_tile_19_1_to_tile_19_2_3),
		.out_wire_0_0(horizontal_tile_19_2_to_tile_19_3_0),
		.out_wire_0_1(horizontal_tile_19_2_to_tile_19_3_1),
		.out_wire_0_2(horizontal_tile_19_2_to_tile_19_3_2),
		.out_wire_0_3(horizontal_tile_19_2_to_tile_19_3_3),
		.in_wire_0_0(horizontal_tile_19_3_to_tile_19_2_0),
		.in_wire_0_1(horizontal_tile_19_3_to_tile_19_2_1),
		.in_wire_0_2(horizontal_tile_19_3_to_tile_19_2_2),
		.in_wire_0_3(horizontal_tile_19_3_to_tile_19_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(611)
	);

	pe_tile pe_tile_19_3(
		.out_wire_3_0(vertical_tile_19_3_to_tile_18_3_0),
		.out_wire_3_1(vertical_tile_19_3_to_tile_18_3_1),
		.out_wire_3_2(vertical_tile_19_3_to_tile_18_3_2),
		.out_wire_3_3(vertical_tile_19_3_to_tile_18_3_3),
		.in_wire_3_0(vertical_tile_18_3_to_tile_19_3_0),
		.in_wire_3_1(vertical_tile_18_3_to_tile_19_3_1),
		.in_wire_3_2(vertical_tile_18_3_to_tile_19_3_2),
		.in_wire_3_3(vertical_tile_18_3_to_tile_19_3_3),
		.out_wire_1_0(vertical_tile_19_3_to_tile_20_3_0),
		.out_wire_1_1(vertical_tile_19_3_to_tile_20_3_1),
		.out_wire_1_2(vertical_tile_19_3_to_tile_20_3_2),
		.out_wire_1_3(vertical_tile_19_3_to_tile_20_3_3),
		.in_wire_1_0(vertical_tile_20_3_to_tile_19_3_0),
		.in_wire_1_1(vertical_tile_20_3_to_tile_19_3_1),
		.in_wire_1_2(vertical_tile_20_3_to_tile_19_3_2),
		.in_wire_1_3(vertical_tile_20_3_to_tile_19_3_3),
		.out_wire_2_0(horizontal_tile_19_3_to_tile_19_2_0),
		.out_wire_2_1(horizontal_tile_19_3_to_tile_19_2_1),
		.out_wire_2_2(horizontal_tile_19_3_to_tile_19_2_2),
		.out_wire_2_3(horizontal_tile_19_3_to_tile_19_2_3),
		.in_wire_2_0(horizontal_tile_19_2_to_tile_19_3_0),
		.in_wire_2_1(horizontal_tile_19_2_to_tile_19_3_1),
		.in_wire_2_2(horizontal_tile_19_2_to_tile_19_3_2),
		.in_wire_2_3(horizontal_tile_19_2_to_tile_19_3_3),
		.out_wire_0_0(horizontal_tile_19_3_to_tile_19_4_0),
		.out_wire_0_1(horizontal_tile_19_3_to_tile_19_4_1),
		.out_wire_0_2(horizontal_tile_19_3_to_tile_19_4_2),
		.out_wire_0_3(horizontal_tile_19_3_to_tile_19_4_3),
		.in_wire_0_0(horizontal_tile_19_4_to_tile_19_3_0),
		.in_wire_0_1(horizontal_tile_19_4_to_tile_19_3_1),
		.in_wire_0_2(horizontal_tile_19_4_to_tile_19_3_2),
		.in_wire_0_3(horizontal_tile_19_4_to_tile_19_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(612)
	);

	pe_tile pe_tile_19_4(
		.out_wire_3_0(vertical_tile_19_4_to_tile_18_4_0),
		.out_wire_3_1(vertical_tile_19_4_to_tile_18_4_1),
		.out_wire_3_2(vertical_tile_19_4_to_tile_18_4_2),
		.out_wire_3_3(vertical_tile_19_4_to_tile_18_4_3),
		.in_wire_3_0(vertical_tile_18_4_to_tile_19_4_0),
		.in_wire_3_1(vertical_tile_18_4_to_tile_19_4_1),
		.in_wire_3_2(vertical_tile_18_4_to_tile_19_4_2),
		.in_wire_3_3(vertical_tile_18_4_to_tile_19_4_3),
		.out_wire_1_0(vertical_tile_19_4_to_tile_20_4_0),
		.out_wire_1_1(vertical_tile_19_4_to_tile_20_4_1),
		.out_wire_1_2(vertical_tile_19_4_to_tile_20_4_2),
		.out_wire_1_3(vertical_tile_19_4_to_tile_20_4_3),
		.in_wire_1_0(vertical_tile_20_4_to_tile_19_4_0),
		.in_wire_1_1(vertical_tile_20_4_to_tile_19_4_1),
		.in_wire_1_2(vertical_tile_20_4_to_tile_19_4_2),
		.in_wire_1_3(vertical_tile_20_4_to_tile_19_4_3),
		.out_wire_2_0(horizontal_tile_19_4_to_tile_19_3_0),
		.out_wire_2_1(horizontal_tile_19_4_to_tile_19_3_1),
		.out_wire_2_2(horizontal_tile_19_4_to_tile_19_3_2),
		.out_wire_2_3(horizontal_tile_19_4_to_tile_19_3_3),
		.in_wire_2_0(horizontal_tile_19_3_to_tile_19_4_0),
		.in_wire_2_1(horizontal_tile_19_3_to_tile_19_4_1),
		.in_wire_2_2(horizontal_tile_19_3_to_tile_19_4_2),
		.in_wire_2_3(horizontal_tile_19_3_to_tile_19_4_3),
		.out_wire_0_0(horizontal_tile_19_4_to_tile_19_5_0),
		.out_wire_0_1(horizontal_tile_19_4_to_tile_19_5_1),
		.out_wire_0_2(horizontal_tile_19_4_to_tile_19_5_2),
		.out_wire_0_3(horizontal_tile_19_4_to_tile_19_5_3),
		.in_wire_0_0(horizontal_tile_19_5_to_tile_19_4_0),
		.in_wire_0_1(horizontal_tile_19_5_to_tile_19_4_1),
		.in_wire_0_2(horizontal_tile_19_5_to_tile_19_4_2),
		.in_wire_0_3(horizontal_tile_19_5_to_tile_19_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(613)
	);

	pe_tile pe_tile_19_5(
		.out_wire_3_0(vertical_tile_19_5_to_tile_18_5_0),
		.out_wire_3_1(vertical_tile_19_5_to_tile_18_5_1),
		.out_wire_3_2(vertical_tile_19_5_to_tile_18_5_2),
		.out_wire_3_3(vertical_tile_19_5_to_tile_18_5_3),
		.in_wire_3_0(vertical_tile_18_5_to_tile_19_5_0),
		.in_wire_3_1(vertical_tile_18_5_to_tile_19_5_1),
		.in_wire_3_2(vertical_tile_18_5_to_tile_19_5_2),
		.in_wire_3_3(vertical_tile_18_5_to_tile_19_5_3),
		.out_wire_1_0(vertical_tile_19_5_to_tile_20_5_0),
		.out_wire_1_1(vertical_tile_19_5_to_tile_20_5_1),
		.out_wire_1_2(vertical_tile_19_5_to_tile_20_5_2),
		.out_wire_1_3(vertical_tile_19_5_to_tile_20_5_3),
		.in_wire_1_0(vertical_tile_20_5_to_tile_19_5_0),
		.in_wire_1_1(vertical_tile_20_5_to_tile_19_5_1),
		.in_wire_1_2(vertical_tile_20_5_to_tile_19_5_2),
		.in_wire_1_3(vertical_tile_20_5_to_tile_19_5_3),
		.out_wire_2_0(horizontal_tile_19_5_to_tile_19_4_0),
		.out_wire_2_1(horizontal_tile_19_5_to_tile_19_4_1),
		.out_wire_2_2(horizontal_tile_19_5_to_tile_19_4_2),
		.out_wire_2_3(horizontal_tile_19_5_to_tile_19_4_3),
		.in_wire_2_0(horizontal_tile_19_4_to_tile_19_5_0),
		.in_wire_2_1(horizontal_tile_19_4_to_tile_19_5_1),
		.in_wire_2_2(horizontal_tile_19_4_to_tile_19_5_2),
		.in_wire_2_3(horizontal_tile_19_4_to_tile_19_5_3),
		.out_wire_0_0(horizontal_tile_19_5_to_tile_19_6_0),
		.out_wire_0_1(horizontal_tile_19_5_to_tile_19_6_1),
		.out_wire_0_2(horizontal_tile_19_5_to_tile_19_6_2),
		.out_wire_0_3(horizontal_tile_19_5_to_tile_19_6_3),
		.in_wire_0_0(horizontal_tile_19_6_to_tile_19_5_0),
		.in_wire_0_1(horizontal_tile_19_6_to_tile_19_5_1),
		.in_wire_0_2(horizontal_tile_19_6_to_tile_19_5_2),
		.in_wire_0_3(horizontal_tile_19_6_to_tile_19_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(614)
	);

	pe_tile pe_tile_19_6(
		.out_wire_3_0(vertical_tile_19_6_to_tile_18_6_0),
		.out_wire_3_1(vertical_tile_19_6_to_tile_18_6_1),
		.out_wire_3_2(vertical_tile_19_6_to_tile_18_6_2),
		.out_wire_3_3(vertical_tile_19_6_to_tile_18_6_3),
		.in_wire_3_0(vertical_tile_18_6_to_tile_19_6_0),
		.in_wire_3_1(vertical_tile_18_6_to_tile_19_6_1),
		.in_wire_3_2(vertical_tile_18_6_to_tile_19_6_2),
		.in_wire_3_3(vertical_tile_18_6_to_tile_19_6_3),
		.out_wire_1_0(vertical_tile_19_6_to_tile_20_6_0),
		.out_wire_1_1(vertical_tile_19_6_to_tile_20_6_1),
		.out_wire_1_2(vertical_tile_19_6_to_tile_20_6_2),
		.out_wire_1_3(vertical_tile_19_6_to_tile_20_6_3),
		.in_wire_1_0(vertical_tile_20_6_to_tile_19_6_0),
		.in_wire_1_1(vertical_tile_20_6_to_tile_19_6_1),
		.in_wire_1_2(vertical_tile_20_6_to_tile_19_6_2),
		.in_wire_1_3(vertical_tile_20_6_to_tile_19_6_3),
		.out_wire_2_0(horizontal_tile_19_6_to_tile_19_5_0),
		.out_wire_2_1(horizontal_tile_19_6_to_tile_19_5_1),
		.out_wire_2_2(horizontal_tile_19_6_to_tile_19_5_2),
		.out_wire_2_3(horizontal_tile_19_6_to_tile_19_5_3),
		.in_wire_2_0(horizontal_tile_19_5_to_tile_19_6_0),
		.in_wire_2_1(horizontal_tile_19_5_to_tile_19_6_1),
		.in_wire_2_2(horizontal_tile_19_5_to_tile_19_6_2),
		.in_wire_2_3(horizontal_tile_19_5_to_tile_19_6_3),
		.out_wire_0_0(horizontal_tile_19_6_to_tile_19_7_0),
		.out_wire_0_1(horizontal_tile_19_6_to_tile_19_7_1),
		.out_wire_0_2(horizontal_tile_19_6_to_tile_19_7_2),
		.out_wire_0_3(horizontal_tile_19_6_to_tile_19_7_3),
		.in_wire_0_0(horizontal_tile_19_7_to_tile_19_6_0),
		.in_wire_0_1(horizontal_tile_19_7_to_tile_19_6_1),
		.in_wire_0_2(horizontal_tile_19_7_to_tile_19_6_2),
		.in_wire_0_3(horizontal_tile_19_7_to_tile_19_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(615)
	);

	pe_tile pe_tile_19_7(
		.out_wire_3_0(vertical_tile_19_7_to_tile_18_7_0),
		.out_wire_3_1(vertical_tile_19_7_to_tile_18_7_1),
		.out_wire_3_2(vertical_tile_19_7_to_tile_18_7_2),
		.out_wire_3_3(vertical_tile_19_7_to_tile_18_7_3),
		.in_wire_3_0(vertical_tile_18_7_to_tile_19_7_0),
		.in_wire_3_1(vertical_tile_18_7_to_tile_19_7_1),
		.in_wire_3_2(vertical_tile_18_7_to_tile_19_7_2),
		.in_wire_3_3(vertical_tile_18_7_to_tile_19_7_3),
		.out_wire_1_0(vertical_tile_19_7_to_tile_20_7_0),
		.out_wire_1_1(vertical_tile_19_7_to_tile_20_7_1),
		.out_wire_1_2(vertical_tile_19_7_to_tile_20_7_2),
		.out_wire_1_3(vertical_tile_19_7_to_tile_20_7_3),
		.in_wire_1_0(vertical_tile_20_7_to_tile_19_7_0),
		.in_wire_1_1(vertical_tile_20_7_to_tile_19_7_1),
		.in_wire_1_2(vertical_tile_20_7_to_tile_19_7_2),
		.in_wire_1_3(vertical_tile_20_7_to_tile_19_7_3),
		.out_wire_2_0(horizontal_tile_19_7_to_tile_19_6_0),
		.out_wire_2_1(horizontal_tile_19_7_to_tile_19_6_1),
		.out_wire_2_2(horizontal_tile_19_7_to_tile_19_6_2),
		.out_wire_2_3(horizontal_tile_19_7_to_tile_19_6_3),
		.in_wire_2_0(horizontal_tile_19_6_to_tile_19_7_0),
		.in_wire_2_1(horizontal_tile_19_6_to_tile_19_7_1),
		.in_wire_2_2(horizontal_tile_19_6_to_tile_19_7_2),
		.in_wire_2_3(horizontal_tile_19_6_to_tile_19_7_3),
		.out_wire_0_0(horizontal_tile_19_7_to_tile_19_8_0),
		.out_wire_0_1(horizontal_tile_19_7_to_tile_19_8_1),
		.out_wire_0_2(horizontal_tile_19_7_to_tile_19_8_2),
		.out_wire_0_3(horizontal_tile_19_7_to_tile_19_8_3),
		.in_wire_0_0(horizontal_tile_19_8_to_tile_19_7_0),
		.in_wire_0_1(horizontal_tile_19_8_to_tile_19_7_1),
		.in_wire_0_2(horizontal_tile_19_8_to_tile_19_7_2),
		.in_wire_0_3(horizontal_tile_19_8_to_tile_19_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(616)
	);

	pe_tile pe_tile_19_8(
		.out_wire_3_0(vertical_tile_19_8_to_tile_18_8_0),
		.out_wire_3_1(vertical_tile_19_8_to_tile_18_8_1),
		.out_wire_3_2(vertical_tile_19_8_to_tile_18_8_2),
		.out_wire_3_3(vertical_tile_19_8_to_tile_18_8_3),
		.in_wire_3_0(vertical_tile_18_8_to_tile_19_8_0),
		.in_wire_3_1(vertical_tile_18_8_to_tile_19_8_1),
		.in_wire_3_2(vertical_tile_18_8_to_tile_19_8_2),
		.in_wire_3_3(vertical_tile_18_8_to_tile_19_8_3),
		.out_wire_1_0(vertical_tile_19_8_to_tile_20_8_0),
		.out_wire_1_1(vertical_tile_19_8_to_tile_20_8_1),
		.out_wire_1_2(vertical_tile_19_8_to_tile_20_8_2),
		.out_wire_1_3(vertical_tile_19_8_to_tile_20_8_3),
		.in_wire_1_0(vertical_tile_20_8_to_tile_19_8_0),
		.in_wire_1_1(vertical_tile_20_8_to_tile_19_8_1),
		.in_wire_1_2(vertical_tile_20_8_to_tile_19_8_2),
		.in_wire_1_3(vertical_tile_20_8_to_tile_19_8_3),
		.out_wire_2_0(horizontal_tile_19_8_to_tile_19_7_0),
		.out_wire_2_1(horizontal_tile_19_8_to_tile_19_7_1),
		.out_wire_2_2(horizontal_tile_19_8_to_tile_19_7_2),
		.out_wire_2_3(horizontal_tile_19_8_to_tile_19_7_3),
		.in_wire_2_0(horizontal_tile_19_7_to_tile_19_8_0),
		.in_wire_2_1(horizontal_tile_19_7_to_tile_19_8_1),
		.in_wire_2_2(horizontal_tile_19_7_to_tile_19_8_2),
		.in_wire_2_3(horizontal_tile_19_7_to_tile_19_8_3),
		.out_wire_0_0(horizontal_tile_19_8_to_tile_19_9_0),
		.out_wire_0_1(horizontal_tile_19_8_to_tile_19_9_1),
		.out_wire_0_2(horizontal_tile_19_8_to_tile_19_9_2),
		.out_wire_0_3(horizontal_tile_19_8_to_tile_19_9_3),
		.in_wire_0_0(horizontal_tile_19_9_to_tile_19_8_0),
		.in_wire_0_1(horizontal_tile_19_9_to_tile_19_8_1),
		.in_wire_0_2(horizontal_tile_19_9_to_tile_19_8_2),
		.in_wire_0_3(horizontal_tile_19_9_to_tile_19_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(617)
	);

	pe_tile pe_tile_19_9(
		.out_wire_3_0(vertical_tile_19_9_to_tile_18_9_0),
		.out_wire_3_1(vertical_tile_19_9_to_tile_18_9_1),
		.out_wire_3_2(vertical_tile_19_9_to_tile_18_9_2),
		.out_wire_3_3(vertical_tile_19_9_to_tile_18_9_3),
		.in_wire_3_0(vertical_tile_18_9_to_tile_19_9_0),
		.in_wire_3_1(vertical_tile_18_9_to_tile_19_9_1),
		.in_wire_3_2(vertical_tile_18_9_to_tile_19_9_2),
		.in_wire_3_3(vertical_tile_18_9_to_tile_19_9_3),
		.out_wire_1_0(vertical_tile_19_9_to_tile_20_9_0),
		.out_wire_1_1(vertical_tile_19_9_to_tile_20_9_1),
		.out_wire_1_2(vertical_tile_19_9_to_tile_20_9_2),
		.out_wire_1_3(vertical_tile_19_9_to_tile_20_9_3),
		.in_wire_1_0(vertical_tile_20_9_to_tile_19_9_0),
		.in_wire_1_1(vertical_tile_20_9_to_tile_19_9_1),
		.in_wire_1_2(vertical_tile_20_9_to_tile_19_9_2),
		.in_wire_1_3(vertical_tile_20_9_to_tile_19_9_3),
		.out_wire_2_0(horizontal_tile_19_9_to_tile_19_8_0),
		.out_wire_2_1(horizontal_tile_19_9_to_tile_19_8_1),
		.out_wire_2_2(horizontal_tile_19_9_to_tile_19_8_2),
		.out_wire_2_3(horizontal_tile_19_9_to_tile_19_8_3),
		.in_wire_2_0(horizontal_tile_19_8_to_tile_19_9_0),
		.in_wire_2_1(horizontal_tile_19_8_to_tile_19_9_1),
		.in_wire_2_2(horizontal_tile_19_8_to_tile_19_9_2),
		.in_wire_2_3(horizontal_tile_19_8_to_tile_19_9_3),
		.out_wire_0_0(horizontal_tile_19_9_to_tile_19_10_0),
		.out_wire_0_1(horizontal_tile_19_9_to_tile_19_10_1),
		.out_wire_0_2(horizontal_tile_19_9_to_tile_19_10_2),
		.out_wire_0_3(horizontal_tile_19_9_to_tile_19_10_3),
		.in_wire_0_0(horizontal_tile_19_10_to_tile_19_9_0),
		.in_wire_0_1(horizontal_tile_19_10_to_tile_19_9_1),
		.in_wire_0_2(horizontal_tile_19_10_to_tile_19_9_2),
		.in_wire_0_3(horizontal_tile_19_10_to_tile_19_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(618)
	);

	pe_tile pe_tile_19_10(
		.out_wire_3_0(vertical_tile_19_10_to_tile_18_10_0),
		.out_wire_3_1(vertical_tile_19_10_to_tile_18_10_1),
		.out_wire_3_2(vertical_tile_19_10_to_tile_18_10_2),
		.out_wire_3_3(vertical_tile_19_10_to_tile_18_10_3),
		.in_wire_3_0(vertical_tile_18_10_to_tile_19_10_0),
		.in_wire_3_1(vertical_tile_18_10_to_tile_19_10_1),
		.in_wire_3_2(vertical_tile_18_10_to_tile_19_10_2),
		.in_wire_3_3(vertical_tile_18_10_to_tile_19_10_3),
		.out_wire_1_0(vertical_tile_19_10_to_tile_20_10_0),
		.out_wire_1_1(vertical_tile_19_10_to_tile_20_10_1),
		.out_wire_1_2(vertical_tile_19_10_to_tile_20_10_2),
		.out_wire_1_3(vertical_tile_19_10_to_tile_20_10_3),
		.in_wire_1_0(vertical_tile_20_10_to_tile_19_10_0),
		.in_wire_1_1(vertical_tile_20_10_to_tile_19_10_1),
		.in_wire_1_2(vertical_tile_20_10_to_tile_19_10_2),
		.in_wire_1_3(vertical_tile_20_10_to_tile_19_10_3),
		.out_wire_2_0(horizontal_tile_19_10_to_tile_19_9_0),
		.out_wire_2_1(horizontal_tile_19_10_to_tile_19_9_1),
		.out_wire_2_2(horizontal_tile_19_10_to_tile_19_9_2),
		.out_wire_2_3(horizontal_tile_19_10_to_tile_19_9_3),
		.in_wire_2_0(horizontal_tile_19_9_to_tile_19_10_0),
		.in_wire_2_1(horizontal_tile_19_9_to_tile_19_10_1),
		.in_wire_2_2(horizontal_tile_19_9_to_tile_19_10_2),
		.in_wire_2_3(horizontal_tile_19_9_to_tile_19_10_3),
		.out_wire_0_0(horizontal_tile_19_10_to_tile_19_11_0),
		.out_wire_0_1(horizontal_tile_19_10_to_tile_19_11_1),
		.out_wire_0_2(horizontal_tile_19_10_to_tile_19_11_2),
		.out_wire_0_3(horizontal_tile_19_10_to_tile_19_11_3),
		.in_wire_0_0(horizontal_tile_19_11_to_tile_19_10_0),
		.in_wire_0_1(horizontal_tile_19_11_to_tile_19_10_1),
		.in_wire_0_2(horizontal_tile_19_11_to_tile_19_10_2),
		.in_wire_0_3(horizontal_tile_19_11_to_tile_19_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(619)
	);

	pe_tile pe_tile_19_11(
		.out_wire_3_0(vertical_tile_19_11_to_tile_18_11_0),
		.out_wire_3_1(vertical_tile_19_11_to_tile_18_11_1),
		.out_wire_3_2(vertical_tile_19_11_to_tile_18_11_2),
		.out_wire_3_3(vertical_tile_19_11_to_tile_18_11_3),
		.in_wire_3_0(vertical_tile_18_11_to_tile_19_11_0),
		.in_wire_3_1(vertical_tile_18_11_to_tile_19_11_1),
		.in_wire_3_2(vertical_tile_18_11_to_tile_19_11_2),
		.in_wire_3_3(vertical_tile_18_11_to_tile_19_11_3),
		.out_wire_1_0(vertical_tile_19_11_to_tile_20_11_0),
		.out_wire_1_1(vertical_tile_19_11_to_tile_20_11_1),
		.out_wire_1_2(vertical_tile_19_11_to_tile_20_11_2),
		.out_wire_1_3(vertical_tile_19_11_to_tile_20_11_3),
		.in_wire_1_0(vertical_tile_20_11_to_tile_19_11_0),
		.in_wire_1_1(vertical_tile_20_11_to_tile_19_11_1),
		.in_wire_1_2(vertical_tile_20_11_to_tile_19_11_2),
		.in_wire_1_3(vertical_tile_20_11_to_tile_19_11_3),
		.out_wire_2_0(horizontal_tile_19_11_to_tile_19_10_0),
		.out_wire_2_1(horizontal_tile_19_11_to_tile_19_10_1),
		.out_wire_2_2(horizontal_tile_19_11_to_tile_19_10_2),
		.out_wire_2_3(horizontal_tile_19_11_to_tile_19_10_3),
		.in_wire_2_0(horizontal_tile_19_10_to_tile_19_11_0),
		.in_wire_2_1(horizontal_tile_19_10_to_tile_19_11_1),
		.in_wire_2_2(horizontal_tile_19_10_to_tile_19_11_2),
		.in_wire_2_3(horizontal_tile_19_10_to_tile_19_11_3),
		.out_wire_0_0(horizontal_tile_19_11_to_tile_19_12_0),
		.out_wire_0_1(horizontal_tile_19_11_to_tile_19_12_1),
		.out_wire_0_2(horizontal_tile_19_11_to_tile_19_12_2),
		.out_wire_0_3(horizontal_tile_19_11_to_tile_19_12_3),
		.in_wire_0_0(horizontal_tile_19_12_to_tile_19_11_0),
		.in_wire_0_1(horizontal_tile_19_12_to_tile_19_11_1),
		.in_wire_0_2(horizontal_tile_19_12_to_tile_19_11_2),
		.in_wire_0_3(horizontal_tile_19_12_to_tile_19_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(620)
	);

	pe_tile pe_tile_19_12(
		.out_wire_3_0(vertical_tile_19_12_to_tile_18_12_0),
		.out_wire_3_1(vertical_tile_19_12_to_tile_18_12_1),
		.out_wire_3_2(vertical_tile_19_12_to_tile_18_12_2),
		.out_wire_3_3(vertical_tile_19_12_to_tile_18_12_3),
		.in_wire_3_0(vertical_tile_18_12_to_tile_19_12_0),
		.in_wire_3_1(vertical_tile_18_12_to_tile_19_12_1),
		.in_wire_3_2(vertical_tile_18_12_to_tile_19_12_2),
		.in_wire_3_3(vertical_tile_18_12_to_tile_19_12_3),
		.out_wire_1_0(vertical_tile_19_12_to_tile_20_12_0),
		.out_wire_1_1(vertical_tile_19_12_to_tile_20_12_1),
		.out_wire_1_2(vertical_tile_19_12_to_tile_20_12_2),
		.out_wire_1_3(vertical_tile_19_12_to_tile_20_12_3),
		.in_wire_1_0(vertical_tile_20_12_to_tile_19_12_0),
		.in_wire_1_1(vertical_tile_20_12_to_tile_19_12_1),
		.in_wire_1_2(vertical_tile_20_12_to_tile_19_12_2),
		.in_wire_1_3(vertical_tile_20_12_to_tile_19_12_3),
		.out_wire_2_0(horizontal_tile_19_12_to_tile_19_11_0),
		.out_wire_2_1(horizontal_tile_19_12_to_tile_19_11_1),
		.out_wire_2_2(horizontal_tile_19_12_to_tile_19_11_2),
		.out_wire_2_3(horizontal_tile_19_12_to_tile_19_11_3),
		.in_wire_2_0(horizontal_tile_19_11_to_tile_19_12_0),
		.in_wire_2_1(horizontal_tile_19_11_to_tile_19_12_1),
		.in_wire_2_2(horizontal_tile_19_11_to_tile_19_12_2),
		.in_wire_2_3(horizontal_tile_19_11_to_tile_19_12_3),
		.out_wire_0_0(horizontal_tile_19_12_to_tile_19_13_0),
		.out_wire_0_1(horizontal_tile_19_12_to_tile_19_13_1),
		.out_wire_0_2(horizontal_tile_19_12_to_tile_19_13_2),
		.out_wire_0_3(horizontal_tile_19_12_to_tile_19_13_3),
		.in_wire_0_0(horizontal_tile_19_13_to_tile_19_12_0),
		.in_wire_0_1(horizontal_tile_19_13_to_tile_19_12_1),
		.in_wire_0_2(horizontal_tile_19_13_to_tile_19_12_2),
		.in_wire_0_3(horizontal_tile_19_13_to_tile_19_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(621)
	);

	pe_tile pe_tile_19_13(
		.out_wire_3_0(vertical_tile_19_13_to_tile_18_13_0),
		.out_wire_3_1(vertical_tile_19_13_to_tile_18_13_1),
		.out_wire_3_2(vertical_tile_19_13_to_tile_18_13_2),
		.out_wire_3_3(vertical_tile_19_13_to_tile_18_13_3),
		.in_wire_3_0(vertical_tile_18_13_to_tile_19_13_0),
		.in_wire_3_1(vertical_tile_18_13_to_tile_19_13_1),
		.in_wire_3_2(vertical_tile_18_13_to_tile_19_13_2),
		.in_wire_3_3(vertical_tile_18_13_to_tile_19_13_3),
		.out_wire_1_0(vertical_tile_19_13_to_tile_20_13_0),
		.out_wire_1_1(vertical_tile_19_13_to_tile_20_13_1),
		.out_wire_1_2(vertical_tile_19_13_to_tile_20_13_2),
		.out_wire_1_3(vertical_tile_19_13_to_tile_20_13_3),
		.in_wire_1_0(vertical_tile_20_13_to_tile_19_13_0),
		.in_wire_1_1(vertical_tile_20_13_to_tile_19_13_1),
		.in_wire_1_2(vertical_tile_20_13_to_tile_19_13_2),
		.in_wire_1_3(vertical_tile_20_13_to_tile_19_13_3),
		.out_wire_2_0(horizontal_tile_19_13_to_tile_19_12_0),
		.out_wire_2_1(horizontal_tile_19_13_to_tile_19_12_1),
		.out_wire_2_2(horizontal_tile_19_13_to_tile_19_12_2),
		.out_wire_2_3(horizontal_tile_19_13_to_tile_19_12_3),
		.in_wire_2_0(horizontal_tile_19_12_to_tile_19_13_0),
		.in_wire_2_1(horizontal_tile_19_12_to_tile_19_13_1),
		.in_wire_2_2(horizontal_tile_19_12_to_tile_19_13_2),
		.in_wire_2_3(horizontal_tile_19_12_to_tile_19_13_3),
		.out_wire_0_0(horizontal_tile_19_13_to_tile_19_14_0),
		.out_wire_0_1(horizontal_tile_19_13_to_tile_19_14_1),
		.out_wire_0_2(horizontal_tile_19_13_to_tile_19_14_2),
		.out_wire_0_3(horizontal_tile_19_13_to_tile_19_14_3),
		.in_wire_0_0(horizontal_tile_19_14_to_tile_19_13_0),
		.in_wire_0_1(horizontal_tile_19_14_to_tile_19_13_1),
		.in_wire_0_2(horizontal_tile_19_14_to_tile_19_13_2),
		.in_wire_0_3(horizontal_tile_19_14_to_tile_19_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(622)
	);

	pe_tile pe_tile_19_14(
		.out_wire_3_0(vertical_tile_19_14_to_tile_18_14_0),
		.out_wire_3_1(vertical_tile_19_14_to_tile_18_14_1),
		.out_wire_3_2(vertical_tile_19_14_to_tile_18_14_2),
		.out_wire_3_3(vertical_tile_19_14_to_tile_18_14_3),
		.in_wire_3_0(vertical_tile_18_14_to_tile_19_14_0),
		.in_wire_3_1(vertical_tile_18_14_to_tile_19_14_1),
		.in_wire_3_2(vertical_tile_18_14_to_tile_19_14_2),
		.in_wire_3_3(vertical_tile_18_14_to_tile_19_14_3),
		.out_wire_1_0(vertical_tile_19_14_to_tile_20_14_0),
		.out_wire_1_1(vertical_tile_19_14_to_tile_20_14_1),
		.out_wire_1_2(vertical_tile_19_14_to_tile_20_14_2),
		.out_wire_1_3(vertical_tile_19_14_to_tile_20_14_3),
		.in_wire_1_0(vertical_tile_20_14_to_tile_19_14_0),
		.in_wire_1_1(vertical_tile_20_14_to_tile_19_14_1),
		.in_wire_1_2(vertical_tile_20_14_to_tile_19_14_2),
		.in_wire_1_3(vertical_tile_20_14_to_tile_19_14_3),
		.out_wire_2_0(horizontal_tile_19_14_to_tile_19_13_0),
		.out_wire_2_1(horizontal_tile_19_14_to_tile_19_13_1),
		.out_wire_2_2(horizontal_tile_19_14_to_tile_19_13_2),
		.out_wire_2_3(horizontal_tile_19_14_to_tile_19_13_3),
		.in_wire_2_0(horizontal_tile_19_13_to_tile_19_14_0),
		.in_wire_2_1(horizontal_tile_19_13_to_tile_19_14_1),
		.in_wire_2_2(horizontal_tile_19_13_to_tile_19_14_2),
		.in_wire_2_3(horizontal_tile_19_13_to_tile_19_14_3),
		.out_wire_0_0(horizontal_tile_19_14_to_tile_19_15_0),
		.out_wire_0_1(horizontal_tile_19_14_to_tile_19_15_1),
		.out_wire_0_2(horizontal_tile_19_14_to_tile_19_15_2),
		.out_wire_0_3(horizontal_tile_19_14_to_tile_19_15_3),
		.in_wire_0_0(horizontal_tile_19_15_to_tile_19_14_0),
		.in_wire_0_1(horizontal_tile_19_15_to_tile_19_14_1),
		.in_wire_0_2(horizontal_tile_19_15_to_tile_19_14_2),
		.in_wire_0_3(horizontal_tile_19_15_to_tile_19_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(623)
	);

	pe_tile pe_tile_19_15(
		.out_wire_3_0(vertical_tile_19_15_to_tile_18_15_0),
		.out_wire_3_1(vertical_tile_19_15_to_tile_18_15_1),
		.out_wire_3_2(vertical_tile_19_15_to_tile_18_15_2),
		.out_wire_3_3(vertical_tile_19_15_to_tile_18_15_3),
		.in_wire_3_0(vertical_tile_18_15_to_tile_19_15_0),
		.in_wire_3_1(vertical_tile_18_15_to_tile_19_15_1),
		.in_wire_3_2(vertical_tile_18_15_to_tile_19_15_2),
		.in_wire_3_3(vertical_tile_18_15_to_tile_19_15_3),
		.out_wire_1_0(vertical_tile_19_15_to_tile_20_15_0),
		.out_wire_1_1(vertical_tile_19_15_to_tile_20_15_1),
		.out_wire_1_2(vertical_tile_19_15_to_tile_20_15_2),
		.out_wire_1_3(vertical_tile_19_15_to_tile_20_15_3),
		.in_wire_1_0(vertical_tile_20_15_to_tile_19_15_0),
		.in_wire_1_1(vertical_tile_20_15_to_tile_19_15_1),
		.in_wire_1_2(vertical_tile_20_15_to_tile_19_15_2),
		.in_wire_1_3(vertical_tile_20_15_to_tile_19_15_3),
		.out_wire_2_0(horizontal_tile_19_15_to_tile_19_14_0),
		.out_wire_2_1(horizontal_tile_19_15_to_tile_19_14_1),
		.out_wire_2_2(horizontal_tile_19_15_to_tile_19_14_2),
		.out_wire_2_3(horizontal_tile_19_15_to_tile_19_14_3),
		.in_wire_2_0(horizontal_tile_19_14_to_tile_19_15_0),
		.in_wire_2_1(horizontal_tile_19_14_to_tile_19_15_1),
		.in_wire_2_2(horizontal_tile_19_14_to_tile_19_15_2),
		.in_wire_2_3(horizontal_tile_19_14_to_tile_19_15_3),
		.out_wire_0_0(horizontal_tile_19_15_to_tile_19_16_0),
		.out_wire_0_1(horizontal_tile_19_15_to_tile_19_16_1),
		.out_wire_0_2(horizontal_tile_19_15_to_tile_19_16_2),
		.out_wire_0_3(horizontal_tile_19_15_to_tile_19_16_3),
		.in_wire_0_0(horizontal_tile_19_16_to_tile_19_15_0),
		.in_wire_0_1(horizontal_tile_19_16_to_tile_19_15_1),
		.in_wire_0_2(horizontal_tile_19_16_to_tile_19_15_2),
		.in_wire_0_3(horizontal_tile_19_16_to_tile_19_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(624)
	);

	pe_tile pe_tile_19_16(
		.out_wire_3_0(vertical_tile_19_16_to_tile_18_16_0),
		.out_wire_3_1(vertical_tile_19_16_to_tile_18_16_1),
		.out_wire_3_2(vertical_tile_19_16_to_tile_18_16_2),
		.out_wire_3_3(vertical_tile_19_16_to_tile_18_16_3),
		.in_wire_3_0(vertical_tile_18_16_to_tile_19_16_0),
		.in_wire_3_1(vertical_tile_18_16_to_tile_19_16_1),
		.in_wire_3_2(vertical_tile_18_16_to_tile_19_16_2),
		.in_wire_3_3(vertical_tile_18_16_to_tile_19_16_3),
		.out_wire_1_0(vertical_tile_19_16_to_tile_20_16_0),
		.out_wire_1_1(vertical_tile_19_16_to_tile_20_16_1),
		.out_wire_1_2(vertical_tile_19_16_to_tile_20_16_2),
		.out_wire_1_3(vertical_tile_19_16_to_tile_20_16_3),
		.in_wire_1_0(vertical_tile_20_16_to_tile_19_16_0),
		.in_wire_1_1(vertical_tile_20_16_to_tile_19_16_1),
		.in_wire_1_2(vertical_tile_20_16_to_tile_19_16_2),
		.in_wire_1_3(vertical_tile_20_16_to_tile_19_16_3),
		.out_wire_2_0(horizontal_tile_19_16_to_tile_19_15_0),
		.out_wire_2_1(horizontal_tile_19_16_to_tile_19_15_1),
		.out_wire_2_2(horizontal_tile_19_16_to_tile_19_15_2),
		.out_wire_2_3(horizontal_tile_19_16_to_tile_19_15_3),
		.in_wire_2_0(horizontal_tile_19_15_to_tile_19_16_0),
		.in_wire_2_1(horizontal_tile_19_15_to_tile_19_16_1),
		.in_wire_2_2(horizontal_tile_19_15_to_tile_19_16_2),
		.in_wire_2_3(horizontal_tile_19_15_to_tile_19_16_3),
		.out_wire_0_0(horizontal_tile_19_16_to_tile_19_17_0),
		.out_wire_0_1(horizontal_tile_19_16_to_tile_19_17_1),
		.out_wire_0_2(horizontal_tile_19_16_to_tile_19_17_2),
		.out_wire_0_3(horizontal_tile_19_16_to_tile_19_17_3),
		.in_wire_0_0(horizontal_tile_19_17_to_tile_19_16_0),
		.in_wire_0_1(horizontal_tile_19_17_to_tile_19_16_1),
		.in_wire_0_2(horizontal_tile_19_17_to_tile_19_16_2),
		.in_wire_0_3(horizontal_tile_19_17_to_tile_19_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(625)
	);

	pe_tile pe_tile_19_17(
		.out_wire_3_0(vertical_tile_19_17_to_tile_18_17_0),
		.out_wire_3_1(vertical_tile_19_17_to_tile_18_17_1),
		.out_wire_3_2(vertical_tile_19_17_to_tile_18_17_2),
		.out_wire_3_3(vertical_tile_19_17_to_tile_18_17_3),
		.in_wire_3_0(vertical_tile_18_17_to_tile_19_17_0),
		.in_wire_3_1(vertical_tile_18_17_to_tile_19_17_1),
		.in_wire_3_2(vertical_tile_18_17_to_tile_19_17_2),
		.in_wire_3_3(vertical_tile_18_17_to_tile_19_17_3),
		.out_wire_1_0(vertical_tile_19_17_to_tile_20_17_0),
		.out_wire_1_1(vertical_tile_19_17_to_tile_20_17_1),
		.out_wire_1_2(vertical_tile_19_17_to_tile_20_17_2),
		.out_wire_1_3(vertical_tile_19_17_to_tile_20_17_3),
		.in_wire_1_0(vertical_tile_20_17_to_tile_19_17_0),
		.in_wire_1_1(vertical_tile_20_17_to_tile_19_17_1),
		.in_wire_1_2(vertical_tile_20_17_to_tile_19_17_2),
		.in_wire_1_3(vertical_tile_20_17_to_tile_19_17_3),
		.out_wire_2_0(horizontal_tile_19_17_to_tile_19_16_0),
		.out_wire_2_1(horizontal_tile_19_17_to_tile_19_16_1),
		.out_wire_2_2(horizontal_tile_19_17_to_tile_19_16_2),
		.out_wire_2_3(horizontal_tile_19_17_to_tile_19_16_3),
		.in_wire_2_0(horizontal_tile_19_16_to_tile_19_17_0),
		.in_wire_2_1(horizontal_tile_19_16_to_tile_19_17_1),
		.in_wire_2_2(horizontal_tile_19_16_to_tile_19_17_2),
		.in_wire_2_3(horizontal_tile_19_16_to_tile_19_17_3),
		.out_wire_0_0(horizontal_tile_19_17_to_tile_19_18_0),
		.out_wire_0_1(horizontal_tile_19_17_to_tile_19_18_1),
		.out_wire_0_2(horizontal_tile_19_17_to_tile_19_18_2),
		.out_wire_0_3(horizontal_tile_19_17_to_tile_19_18_3),
		.in_wire_0_0(horizontal_tile_19_18_to_tile_19_17_0),
		.in_wire_0_1(horizontal_tile_19_18_to_tile_19_17_1),
		.in_wire_0_2(horizontal_tile_19_18_to_tile_19_17_2),
		.in_wire_0_3(horizontal_tile_19_18_to_tile_19_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(626)
	);

	pe_tile pe_tile_19_18(
		.out_wire_3_0(vertical_tile_19_18_to_tile_18_18_0),
		.out_wire_3_1(vertical_tile_19_18_to_tile_18_18_1),
		.out_wire_3_2(vertical_tile_19_18_to_tile_18_18_2),
		.out_wire_3_3(vertical_tile_19_18_to_tile_18_18_3),
		.in_wire_3_0(vertical_tile_18_18_to_tile_19_18_0),
		.in_wire_3_1(vertical_tile_18_18_to_tile_19_18_1),
		.in_wire_3_2(vertical_tile_18_18_to_tile_19_18_2),
		.in_wire_3_3(vertical_tile_18_18_to_tile_19_18_3),
		.out_wire_1_0(vertical_tile_19_18_to_tile_20_18_0),
		.out_wire_1_1(vertical_tile_19_18_to_tile_20_18_1),
		.out_wire_1_2(vertical_tile_19_18_to_tile_20_18_2),
		.out_wire_1_3(vertical_tile_19_18_to_tile_20_18_3),
		.in_wire_1_0(vertical_tile_20_18_to_tile_19_18_0),
		.in_wire_1_1(vertical_tile_20_18_to_tile_19_18_1),
		.in_wire_1_2(vertical_tile_20_18_to_tile_19_18_2),
		.in_wire_1_3(vertical_tile_20_18_to_tile_19_18_3),
		.out_wire_2_0(horizontal_tile_19_18_to_tile_19_17_0),
		.out_wire_2_1(horizontal_tile_19_18_to_tile_19_17_1),
		.out_wire_2_2(horizontal_tile_19_18_to_tile_19_17_2),
		.out_wire_2_3(horizontal_tile_19_18_to_tile_19_17_3),
		.in_wire_2_0(horizontal_tile_19_17_to_tile_19_18_0),
		.in_wire_2_1(horizontal_tile_19_17_to_tile_19_18_1),
		.in_wire_2_2(horizontal_tile_19_17_to_tile_19_18_2),
		.in_wire_2_3(horizontal_tile_19_17_to_tile_19_18_3),
		.out_wire_0_0(horizontal_tile_19_18_to_tile_19_19_0),
		.out_wire_0_1(horizontal_tile_19_18_to_tile_19_19_1),
		.out_wire_0_2(horizontal_tile_19_18_to_tile_19_19_2),
		.out_wire_0_3(horizontal_tile_19_18_to_tile_19_19_3),
		.in_wire_0_0(horizontal_tile_19_19_to_tile_19_18_0),
		.in_wire_0_1(horizontal_tile_19_19_to_tile_19_18_1),
		.in_wire_0_2(horizontal_tile_19_19_to_tile_19_18_2),
		.in_wire_0_3(horizontal_tile_19_19_to_tile_19_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(627)
	);

	pe_tile pe_tile_19_19(
		.out_wire_3_0(vertical_tile_19_19_to_tile_18_19_0),
		.out_wire_3_1(vertical_tile_19_19_to_tile_18_19_1),
		.out_wire_3_2(vertical_tile_19_19_to_tile_18_19_2),
		.out_wire_3_3(vertical_tile_19_19_to_tile_18_19_3),
		.in_wire_3_0(vertical_tile_18_19_to_tile_19_19_0),
		.in_wire_3_1(vertical_tile_18_19_to_tile_19_19_1),
		.in_wire_3_2(vertical_tile_18_19_to_tile_19_19_2),
		.in_wire_3_3(vertical_tile_18_19_to_tile_19_19_3),
		.out_wire_1_0(vertical_tile_19_19_to_tile_20_19_0),
		.out_wire_1_1(vertical_tile_19_19_to_tile_20_19_1),
		.out_wire_1_2(vertical_tile_19_19_to_tile_20_19_2),
		.out_wire_1_3(vertical_tile_19_19_to_tile_20_19_3),
		.in_wire_1_0(vertical_tile_20_19_to_tile_19_19_0),
		.in_wire_1_1(vertical_tile_20_19_to_tile_19_19_1),
		.in_wire_1_2(vertical_tile_20_19_to_tile_19_19_2),
		.in_wire_1_3(vertical_tile_20_19_to_tile_19_19_3),
		.out_wire_2_0(horizontal_tile_19_19_to_tile_19_18_0),
		.out_wire_2_1(horizontal_tile_19_19_to_tile_19_18_1),
		.out_wire_2_2(horizontal_tile_19_19_to_tile_19_18_2),
		.out_wire_2_3(horizontal_tile_19_19_to_tile_19_18_3),
		.in_wire_2_0(horizontal_tile_19_18_to_tile_19_19_0),
		.in_wire_2_1(horizontal_tile_19_18_to_tile_19_19_1),
		.in_wire_2_2(horizontal_tile_19_18_to_tile_19_19_2),
		.in_wire_2_3(horizontal_tile_19_18_to_tile_19_19_3),
		.out_wire_0_0(horizontal_tile_19_19_to_tile_19_20_0),
		.out_wire_0_1(horizontal_tile_19_19_to_tile_19_20_1),
		.out_wire_0_2(horizontal_tile_19_19_to_tile_19_20_2),
		.out_wire_0_3(horizontal_tile_19_19_to_tile_19_20_3),
		.in_wire_0_0(horizontal_tile_19_20_to_tile_19_19_0),
		.in_wire_0_1(horizontal_tile_19_20_to_tile_19_19_1),
		.in_wire_0_2(horizontal_tile_19_20_to_tile_19_19_2),
		.in_wire_0_3(horizontal_tile_19_20_to_tile_19_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(628)
	);

	pe_tile pe_tile_19_20(
		.out_wire_3_0(vertical_tile_19_20_to_tile_18_20_0),
		.out_wire_3_1(vertical_tile_19_20_to_tile_18_20_1),
		.out_wire_3_2(vertical_tile_19_20_to_tile_18_20_2),
		.out_wire_3_3(vertical_tile_19_20_to_tile_18_20_3),
		.in_wire_3_0(vertical_tile_18_20_to_tile_19_20_0),
		.in_wire_3_1(vertical_tile_18_20_to_tile_19_20_1),
		.in_wire_3_2(vertical_tile_18_20_to_tile_19_20_2),
		.in_wire_3_3(vertical_tile_18_20_to_tile_19_20_3),
		.out_wire_1_0(vertical_tile_19_20_to_tile_20_20_0),
		.out_wire_1_1(vertical_tile_19_20_to_tile_20_20_1),
		.out_wire_1_2(vertical_tile_19_20_to_tile_20_20_2),
		.out_wire_1_3(vertical_tile_19_20_to_tile_20_20_3),
		.in_wire_1_0(vertical_tile_20_20_to_tile_19_20_0),
		.in_wire_1_1(vertical_tile_20_20_to_tile_19_20_1),
		.in_wire_1_2(vertical_tile_20_20_to_tile_19_20_2),
		.in_wire_1_3(vertical_tile_20_20_to_tile_19_20_3),
		.out_wire_2_0(horizontal_tile_19_20_to_tile_19_19_0),
		.out_wire_2_1(horizontal_tile_19_20_to_tile_19_19_1),
		.out_wire_2_2(horizontal_tile_19_20_to_tile_19_19_2),
		.out_wire_2_3(horizontal_tile_19_20_to_tile_19_19_3),
		.in_wire_2_0(horizontal_tile_19_19_to_tile_19_20_0),
		.in_wire_2_1(horizontal_tile_19_19_to_tile_19_20_1),
		.in_wire_2_2(horizontal_tile_19_19_to_tile_19_20_2),
		.in_wire_2_3(horizontal_tile_19_19_to_tile_19_20_3),
		.out_wire_0_0(horizontal_tile_19_20_to_tile_19_21_0),
		.out_wire_0_1(horizontal_tile_19_20_to_tile_19_21_1),
		.out_wire_0_2(horizontal_tile_19_20_to_tile_19_21_2),
		.out_wire_0_3(horizontal_tile_19_20_to_tile_19_21_3),
		.in_wire_0_0(horizontal_tile_19_21_to_tile_19_20_0),
		.in_wire_0_1(horizontal_tile_19_21_to_tile_19_20_1),
		.in_wire_0_2(horizontal_tile_19_21_to_tile_19_20_2),
		.in_wire_0_3(horizontal_tile_19_21_to_tile_19_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(629)
	);

	pe_tile pe_tile_19_21(
		.out_wire_3_0(vertical_tile_19_21_to_tile_18_21_0),
		.out_wire_3_1(vertical_tile_19_21_to_tile_18_21_1),
		.out_wire_3_2(vertical_tile_19_21_to_tile_18_21_2),
		.out_wire_3_3(vertical_tile_19_21_to_tile_18_21_3),
		.in_wire_3_0(vertical_tile_18_21_to_tile_19_21_0),
		.in_wire_3_1(vertical_tile_18_21_to_tile_19_21_1),
		.in_wire_3_2(vertical_tile_18_21_to_tile_19_21_2),
		.in_wire_3_3(vertical_tile_18_21_to_tile_19_21_3),
		.out_wire_1_0(vertical_tile_19_21_to_tile_20_21_0),
		.out_wire_1_1(vertical_tile_19_21_to_tile_20_21_1),
		.out_wire_1_2(vertical_tile_19_21_to_tile_20_21_2),
		.out_wire_1_3(vertical_tile_19_21_to_tile_20_21_3),
		.in_wire_1_0(vertical_tile_20_21_to_tile_19_21_0),
		.in_wire_1_1(vertical_tile_20_21_to_tile_19_21_1),
		.in_wire_1_2(vertical_tile_20_21_to_tile_19_21_2),
		.in_wire_1_3(vertical_tile_20_21_to_tile_19_21_3),
		.out_wire_2_0(horizontal_tile_19_21_to_tile_19_20_0),
		.out_wire_2_1(horizontal_tile_19_21_to_tile_19_20_1),
		.out_wire_2_2(horizontal_tile_19_21_to_tile_19_20_2),
		.out_wire_2_3(horizontal_tile_19_21_to_tile_19_20_3),
		.in_wire_2_0(horizontal_tile_19_20_to_tile_19_21_0),
		.in_wire_2_1(horizontal_tile_19_20_to_tile_19_21_1),
		.in_wire_2_2(horizontal_tile_19_20_to_tile_19_21_2),
		.in_wire_2_3(horizontal_tile_19_20_to_tile_19_21_3),
		.out_wire_0_0(horizontal_tile_19_21_to_tile_19_22_0),
		.out_wire_0_1(horizontal_tile_19_21_to_tile_19_22_1),
		.out_wire_0_2(horizontal_tile_19_21_to_tile_19_22_2),
		.out_wire_0_3(horizontal_tile_19_21_to_tile_19_22_3),
		.in_wire_0_0(horizontal_tile_19_22_to_tile_19_21_0),
		.in_wire_0_1(horizontal_tile_19_22_to_tile_19_21_1),
		.in_wire_0_2(horizontal_tile_19_22_to_tile_19_21_2),
		.in_wire_0_3(horizontal_tile_19_22_to_tile_19_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(630)
	);

	pe_tile pe_tile_19_22(
		.out_wire_3_0(vertical_tile_19_22_to_tile_18_22_0),
		.out_wire_3_1(vertical_tile_19_22_to_tile_18_22_1),
		.out_wire_3_2(vertical_tile_19_22_to_tile_18_22_2),
		.out_wire_3_3(vertical_tile_19_22_to_tile_18_22_3),
		.in_wire_3_0(vertical_tile_18_22_to_tile_19_22_0),
		.in_wire_3_1(vertical_tile_18_22_to_tile_19_22_1),
		.in_wire_3_2(vertical_tile_18_22_to_tile_19_22_2),
		.in_wire_3_3(vertical_tile_18_22_to_tile_19_22_3),
		.out_wire_1_0(vertical_tile_19_22_to_tile_20_22_0),
		.out_wire_1_1(vertical_tile_19_22_to_tile_20_22_1),
		.out_wire_1_2(vertical_tile_19_22_to_tile_20_22_2),
		.out_wire_1_3(vertical_tile_19_22_to_tile_20_22_3),
		.in_wire_1_0(vertical_tile_20_22_to_tile_19_22_0),
		.in_wire_1_1(vertical_tile_20_22_to_tile_19_22_1),
		.in_wire_1_2(vertical_tile_20_22_to_tile_19_22_2),
		.in_wire_1_3(vertical_tile_20_22_to_tile_19_22_3),
		.out_wire_2_0(horizontal_tile_19_22_to_tile_19_21_0),
		.out_wire_2_1(horizontal_tile_19_22_to_tile_19_21_1),
		.out_wire_2_2(horizontal_tile_19_22_to_tile_19_21_2),
		.out_wire_2_3(horizontal_tile_19_22_to_tile_19_21_3),
		.in_wire_2_0(horizontal_tile_19_21_to_tile_19_22_0),
		.in_wire_2_1(horizontal_tile_19_21_to_tile_19_22_1),
		.in_wire_2_2(horizontal_tile_19_21_to_tile_19_22_2),
		.in_wire_2_3(horizontal_tile_19_21_to_tile_19_22_3),
		.out_wire_0_0(horizontal_tile_19_22_to_tile_19_23_0),
		.out_wire_0_1(horizontal_tile_19_22_to_tile_19_23_1),
		.out_wire_0_2(horizontal_tile_19_22_to_tile_19_23_2),
		.out_wire_0_3(horizontal_tile_19_22_to_tile_19_23_3),
		.in_wire_0_0(horizontal_tile_19_23_to_tile_19_22_0),
		.in_wire_0_1(horizontal_tile_19_23_to_tile_19_22_1),
		.in_wire_0_2(horizontal_tile_19_23_to_tile_19_22_2),
		.in_wire_0_3(horizontal_tile_19_23_to_tile_19_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(631)
	);

	pe_tile pe_tile_19_23(
		.out_wire_3_0(vertical_tile_19_23_to_tile_18_23_0),
		.out_wire_3_1(vertical_tile_19_23_to_tile_18_23_1),
		.out_wire_3_2(vertical_tile_19_23_to_tile_18_23_2),
		.out_wire_3_3(vertical_tile_19_23_to_tile_18_23_3),
		.in_wire_3_0(vertical_tile_18_23_to_tile_19_23_0),
		.in_wire_3_1(vertical_tile_18_23_to_tile_19_23_1),
		.in_wire_3_2(vertical_tile_18_23_to_tile_19_23_2),
		.in_wire_3_3(vertical_tile_18_23_to_tile_19_23_3),
		.out_wire_1_0(vertical_tile_19_23_to_tile_20_23_0),
		.out_wire_1_1(vertical_tile_19_23_to_tile_20_23_1),
		.out_wire_1_2(vertical_tile_19_23_to_tile_20_23_2),
		.out_wire_1_3(vertical_tile_19_23_to_tile_20_23_3),
		.in_wire_1_0(vertical_tile_20_23_to_tile_19_23_0),
		.in_wire_1_1(vertical_tile_20_23_to_tile_19_23_1),
		.in_wire_1_2(vertical_tile_20_23_to_tile_19_23_2),
		.in_wire_1_3(vertical_tile_20_23_to_tile_19_23_3),
		.out_wire_2_0(horizontal_tile_19_23_to_tile_19_22_0),
		.out_wire_2_1(horizontal_tile_19_23_to_tile_19_22_1),
		.out_wire_2_2(horizontal_tile_19_23_to_tile_19_22_2),
		.out_wire_2_3(horizontal_tile_19_23_to_tile_19_22_3),
		.in_wire_2_0(horizontal_tile_19_22_to_tile_19_23_0),
		.in_wire_2_1(horizontal_tile_19_22_to_tile_19_23_1),
		.in_wire_2_2(horizontal_tile_19_22_to_tile_19_23_2),
		.in_wire_2_3(horizontal_tile_19_22_to_tile_19_23_3),
		.out_wire_0_0(horizontal_tile_19_23_to_tile_19_24_0),
		.out_wire_0_1(horizontal_tile_19_23_to_tile_19_24_1),
		.out_wire_0_2(horizontal_tile_19_23_to_tile_19_24_2),
		.out_wire_0_3(horizontal_tile_19_23_to_tile_19_24_3),
		.in_wire_0_0(horizontal_tile_19_24_to_tile_19_23_0),
		.in_wire_0_1(horizontal_tile_19_24_to_tile_19_23_1),
		.in_wire_0_2(horizontal_tile_19_24_to_tile_19_23_2),
		.in_wire_0_3(horizontal_tile_19_24_to_tile_19_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(632)
	);

	pe_tile pe_tile_19_24(
		.out_wire_3_0(vertical_tile_19_24_to_tile_18_24_0),
		.out_wire_3_1(vertical_tile_19_24_to_tile_18_24_1),
		.out_wire_3_2(vertical_tile_19_24_to_tile_18_24_2),
		.out_wire_3_3(vertical_tile_19_24_to_tile_18_24_3),
		.in_wire_3_0(vertical_tile_18_24_to_tile_19_24_0),
		.in_wire_3_1(vertical_tile_18_24_to_tile_19_24_1),
		.in_wire_3_2(vertical_tile_18_24_to_tile_19_24_2),
		.in_wire_3_3(vertical_tile_18_24_to_tile_19_24_3),
		.out_wire_1_0(vertical_tile_19_24_to_tile_20_24_0),
		.out_wire_1_1(vertical_tile_19_24_to_tile_20_24_1),
		.out_wire_1_2(vertical_tile_19_24_to_tile_20_24_2),
		.out_wire_1_3(vertical_tile_19_24_to_tile_20_24_3),
		.in_wire_1_0(vertical_tile_20_24_to_tile_19_24_0),
		.in_wire_1_1(vertical_tile_20_24_to_tile_19_24_1),
		.in_wire_1_2(vertical_tile_20_24_to_tile_19_24_2),
		.in_wire_1_3(vertical_tile_20_24_to_tile_19_24_3),
		.out_wire_2_0(horizontal_tile_19_24_to_tile_19_23_0),
		.out_wire_2_1(horizontal_tile_19_24_to_tile_19_23_1),
		.out_wire_2_2(horizontal_tile_19_24_to_tile_19_23_2),
		.out_wire_2_3(horizontal_tile_19_24_to_tile_19_23_3),
		.in_wire_2_0(horizontal_tile_19_23_to_tile_19_24_0),
		.in_wire_2_1(horizontal_tile_19_23_to_tile_19_24_1),
		.in_wire_2_2(horizontal_tile_19_23_to_tile_19_24_2),
		.in_wire_2_3(horizontal_tile_19_23_to_tile_19_24_3),
		.out_wire_0_0(horizontal_tile_19_24_to_tile_19_25_0),
		.out_wire_0_1(horizontal_tile_19_24_to_tile_19_25_1),
		.out_wire_0_2(horizontal_tile_19_24_to_tile_19_25_2),
		.out_wire_0_3(horizontal_tile_19_24_to_tile_19_25_3),
		.in_wire_0_0(horizontal_tile_19_25_to_tile_19_24_0),
		.in_wire_0_1(horizontal_tile_19_25_to_tile_19_24_1),
		.in_wire_0_2(horizontal_tile_19_25_to_tile_19_24_2),
		.in_wire_0_3(horizontal_tile_19_25_to_tile_19_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(633)
	);

	pe_tile pe_tile_19_25(
		.out_wire_3_0(vertical_tile_19_25_to_tile_18_25_0),
		.out_wire_3_1(vertical_tile_19_25_to_tile_18_25_1),
		.out_wire_3_2(vertical_tile_19_25_to_tile_18_25_2),
		.out_wire_3_3(vertical_tile_19_25_to_tile_18_25_3),
		.in_wire_3_0(vertical_tile_18_25_to_tile_19_25_0),
		.in_wire_3_1(vertical_tile_18_25_to_tile_19_25_1),
		.in_wire_3_2(vertical_tile_18_25_to_tile_19_25_2),
		.in_wire_3_3(vertical_tile_18_25_to_tile_19_25_3),
		.out_wire_1_0(vertical_tile_19_25_to_tile_20_25_0),
		.out_wire_1_1(vertical_tile_19_25_to_tile_20_25_1),
		.out_wire_1_2(vertical_tile_19_25_to_tile_20_25_2),
		.out_wire_1_3(vertical_tile_19_25_to_tile_20_25_3),
		.in_wire_1_0(vertical_tile_20_25_to_tile_19_25_0),
		.in_wire_1_1(vertical_tile_20_25_to_tile_19_25_1),
		.in_wire_1_2(vertical_tile_20_25_to_tile_19_25_2),
		.in_wire_1_3(vertical_tile_20_25_to_tile_19_25_3),
		.out_wire_2_0(horizontal_tile_19_25_to_tile_19_24_0),
		.out_wire_2_1(horizontal_tile_19_25_to_tile_19_24_1),
		.out_wire_2_2(horizontal_tile_19_25_to_tile_19_24_2),
		.out_wire_2_3(horizontal_tile_19_25_to_tile_19_24_3),
		.in_wire_2_0(horizontal_tile_19_24_to_tile_19_25_0),
		.in_wire_2_1(horizontal_tile_19_24_to_tile_19_25_1),
		.in_wire_2_2(horizontal_tile_19_24_to_tile_19_25_2),
		.in_wire_2_3(horizontal_tile_19_24_to_tile_19_25_3),
		.out_wire_0_0(horizontal_tile_19_25_to_tile_19_26_0),
		.out_wire_0_1(horizontal_tile_19_25_to_tile_19_26_1),
		.out_wire_0_2(horizontal_tile_19_25_to_tile_19_26_2),
		.out_wire_0_3(horizontal_tile_19_25_to_tile_19_26_3),
		.in_wire_0_0(horizontal_tile_19_26_to_tile_19_25_0),
		.in_wire_0_1(horizontal_tile_19_26_to_tile_19_25_1),
		.in_wire_0_2(horizontal_tile_19_26_to_tile_19_25_2),
		.in_wire_0_3(horizontal_tile_19_26_to_tile_19_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(634)
	);

	pe_tile pe_tile_19_26(
		.out_wire_3_0(vertical_tile_19_26_to_tile_18_26_0),
		.out_wire_3_1(vertical_tile_19_26_to_tile_18_26_1),
		.out_wire_3_2(vertical_tile_19_26_to_tile_18_26_2),
		.out_wire_3_3(vertical_tile_19_26_to_tile_18_26_3),
		.in_wire_3_0(vertical_tile_18_26_to_tile_19_26_0),
		.in_wire_3_1(vertical_tile_18_26_to_tile_19_26_1),
		.in_wire_3_2(vertical_tile_18_26_to_tile_19_26_2),
		.in_wire_3_3(vertical_tile_18_26_to_tile_19_26_3),
		.out_wire_1_0(vertical_tile_19_26_to_tile_20_26_0),
		.out_wire_1_1(vertical_tile_19_26_to_tile_20_26_1),
		.out_wire_1_2(vertical_tile_19_26_to_tile_20_26_2),
		.out_wire_1_3(vertical_tile_19_26_to_tile_20_26_3),
		.in_wire_1_0(vertical_tile_20_26_to_tile_19_26_0),
		.in_wire_1_1(vertical_tile_20_26_to_tile_19_26_1),
		.in_wire_1_2(vertical_tile_20_26_to_tile_19_26_2),
		.in_wire_1_3(vertical_tile_20_26_to_tile_19_26_3),
		.out_wire_2_0(horizontal_tile_19_26_to_tile_19_25_0),
		.out_wire_2_1(horizontal_tile_19_26_to_tile_19_25_1),
		.out_wire_2_2(horizontal_tile_19_26_to_tile_19_25_2),
		.out_wire_2_3(horizontal_tile_19_26_to_tile_19_25_3),
		.in_wire_2_0(horizontal_tile_19_25_to_tile_19_26_0),
		.in_wire_2_1(horizontal_tile_19_25_to_tile_19_26_1),
		.in_wire_2_2(horizontal_tile_19_25_to_tile_19_26_2),
		.in_wire_2_3(horizontal_tile_19_25_to_tile_19_26_3),
		.out_wire_0_0(horizontal_tile_19_26_to_tile_19_27_0),
		.out_wire_0_1(horizontal_tile_19_26_to_tile_19_27_1),
		.out_wire_0_2(horizontal_tile_19_26_to_tile_19_27_2),
		.out_wire_0_3(horizontal_tile_19_26_to_tile_19_27_3),
		.in_wire_0_0(horizontal_tile_19_27_to_tile_19_26_0),
		.in_wire_0_1(horizontal_tile_19_27_to_tile_19_26_1),
		.in_wire_0_2(horizontal_tile_19_27_to_tile_19_26_2),
		.in_wire_0_3(horizontal_tile_19_27_to_tile_19_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(635)
	);

	pe_tile pe_tile_19_27(
		.out_wire_3_0(vertical_tile_19_27_to_tile_18_27_0),
		.out_wire_3_1(vertical_tile_19_27_to_tile_18_27_1),
		.out_wire_3_2(vertical_tile_19_27_to_tile_18_27_2),
		.out_wire_3_3(vertical_tile_19_27_to_tile_18_27_3),
		.in_wire_3_0(vertical_tile_18_27_to_tile_19_27_0),
		.in_wire_3_1(vertical_tile_18_27_to_tile_19_27_1),
		.in_wire_3_2(vertical_tile_18_27_to_tile_19_27_2),
		.in_wire_3_3(vertical_tile_18_27_to_tile_19_27_3),
		.out_wire_1_0(vertical_tile_19_27_to_tile_20_27_0),
		.out_wire_1_1(vertical_tile_19_27_to_tile_20_27_1),
		.out_wire_1_2(vertical_tile_19_27_to_tile_20_27_2),
		.out_wire_1_3(vertical_tile_19_27_to_tile_20_27_3),
		.in_wire_1_0(vertical_tile_20_27_to_tile_19_27_0),
		.in_wire_1_1(vertical_tile_20_27_to_tile_19_27_1),
		.in_wire_1_2(vertical_tile_20_27_to_tile_19_27_2),
		.in_wire_1_3(vertical_tile_20_27_to_tile_19_27_3),
		.out_wire_2_0(horizontal_tile_19_27_to_tile_19_26_0),
		.out_wire_2_1(horizontal_tile_19_27_to_tile_19_26_1),
		.out_wire_2_2(horizontal_tile_19_27_to_tile_19_26_2),
		.out_wire_2_3(horizontal_tile_19_27_to_tile_19_26_3),
		.in_wire_2_0(horizontal_tile_19_26_to_tile_19_27_0),
		.in_wire_2_1(horizontal_tile_19_26_to_tile_19_27_1),
		.in_wire_2_2(horizontal_tile_19_26_to_tile_19_27_2),
		.in_wire_2_3(horizontal_tile_19_26_to_tile_19_27_3),
		.out_wire_0_0(horizontal_tile_19_27_to_tile_19_28_0),
		.out_wire_0_1(horizontal_tile_19_27_to_tile_19_28_1),
		.out_wire_0_2(horizontal_tile_19_27_to_tile_19_28_2),
		.out_wire_0_3(horizontal_tile_19_27_to_tile_19_28_3),
		.in_wire_0_0(horizontal_tile_19_28_to_tile_19_27_0),
		.in_wire_0_1(horizontal_tile_19_28_to_tile_19_27_1),
		.in_wire_0_2(horizontal_tile_19_28_to_tile_19_27_2),
		.in_wire_0_3(horizontal_tile_19_28_to_tile_19_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(636)
	);

	pe_tile pe_tile_19_28(
		.out_wire_3_0(vertical_tile_19_28_to_tile_18_28_0),
		.out_wire_3_1(vertical_tile_19_28_to_tile_18_28_1),
		.out_wire_3_2(vertical_tile_19_28_to_tile_18_28_2),
		.out_wire_3_3(vertical_tile_19_28_to_tile_18_28_3),
		.in_wire_3_0(vertical_tile_18_28_to_tile_19_28_0),
		.in_wire_3_1(vertical_tile_18_28_to_tile_19_28_1),
		.in_wire_3_2(vertical_tile_18_28_to_tile_19_28_2),
		.in_wire_3_3(vertical_tile_18_28_to_tile_19_28_3),
		.out_wire_1_0(vertical_tile_19_28_to_tile_20_28_0),
		.out_wire_1_1(vertical_tile_19_28_to_tile_20_28_1),
		.out_wire_1_2(vertical_tile_19_28_to_tile_20_28_2),
		.out_wire_1_3(vertical_tile_19_28_to_tile_20_28_3),
		.in_wire_1_0(vertical_tile_20_28_to_tile_19_28_0),
		.in_wire_1_1(vertical_tile_20_28_to_tile_19_28_1),
		.in_wire_1_2(vertical_tile_20_28_to_tile_19_28_2),
		.in_wire_1_3(vertical_tile_20_28_to_tile_19_28_3),
		.out_wire_2_0(horizontal_tile_19_28_to_tile_19_27_0),
		.out_wire_2_1(horizontal_tile_19_28_to_tile_19_27_1),
		.out_wire_2_2(horizontal_tile_19_28_to_tile_19_27_2),
		.out_wire_2_3(horizontal_tile_19_28_to_tile_19_27_3),
		.in_wire_2_0(horizontal_tile_19_27_to_tile_19_28_0),
		.in_wire_2_1(horizontal_tile_19_27_to_tile_19_28_1),
		.in_wire_2_2(horizontal_tile_19_27_to_tile_19_28_2),
		.in_wire_2_3(horizontal_tile_19_27_to_tile_19_28_3),
		.out_wire_0_0(horizontal_tile_19_28_to_tile_19_29_0),
		.out_wire_0_1(horizontal_tile_19_28_to_tile_19_29_1),
		.out_wire_0_2(horizontal_tile_19_28_to_tile_19_29_2),
		.out_wire_0_3(horizontal_tile_19_28_to_tile_19_29_3),
		.in_wire_0_0(horizontal_tile_19_29_to_tile_19_28_0),
		.in_wire_0_1(horizontal_tile_19_29_to_tile_19_28_1),
		.in_wire_0_2(horizontal_tile_19_29_to_tile_19_28_2),
		.in_wire_0_3(horizontal_tile_19_29_to_tile_19_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(637)
	);

	pe_tile pe_tile_19_29(
		.out_wire_3_0(vertical_tile_19_29_to_tile_18_29_0),
		.out_wire_3_1(vertical_tile_19_29_to_tile_18_29_1),
		.out_wire_3_2(vertical_tile_19_29_to_tile_18_29_2),
		.out_wire_3_3(vertical_tile_19_29_to_tile_18_29_3),
		.in_wire_3_0(vertical_tile_18_29_to_tile_19_29_0),
		.in_wire_3_1(vertical_tile_18_29_to_tile_19_29_1),
		.in_wire_3_2(vertical_tile_18_29_to_tile_19_29_2),
		.in_wire_3_3(vertical_tile_18_29_to_tile_19_29_3),
		.out_wire_1_0(vertical_tile_19_29_to_tile_20_29_0),
		.out_wire_1_1(vertical_tile_19_29_to_tile_20_29_1),
		.out_wire_1_2(vertical_tile_19_29_to_tile_20_29_2),
		.out_wire_1_3(vertical_tile_19_29_to_tile_20_29_3),
		.in_wire_1_0(vertical_tile_20_29_to_tile_19_29_0),
		.in_wire_1_1(vertical_tile_20_29_to_tile_19_29_1),
		.in_wire_1_2(vertical_tile_20_29_to_tile_19_29_2),
		.in_wire_1_3(vertical_tile_20_29_to_tile_19_29_3),
		.out_wire_2_0(horizontal_tile_19_29_to_tile_19_28_0),
		.out_wire_2_1(horizontal_tile_19_29_to_tile_19_28_1),
		.out_wire_2_2(horizontal_tile_19_29_to_tile_19_28_2),
		.out_wire_2_3(horizontal_tile_19_29_to_tile_19_28_3),
		.in_wire_2_0(horizontal_tile_19_28_to_tile_19_29_0),
		.in_wire_2_1(horizontal_tile_19_28_to_tile_19_29_1),
		.in_wire_2_2(horizontal_tile_19_28_to_tile_19_29_2),
		.in_wire_2_3(horizontal_tile_19_28_to_tile_19_29_3),
		.out_wire_0_0(horizontal_tile_19_29_to_tile_19_30_0),
		.out_wire_0_1(horizontal_tile_19_29_to_tile_19_30_1),
		.out_wire_0_2(horizontal_tile_19_29_to_tile_19_30_2),
		.out_wire_0_3(horizontal_tile_19_29_to_tile_19_30_3),
		.in_wire_0_0(horizontal_tile_19_30_to_tile_19_29_0),
		.in_wire_0_1(horizontal_tile_19_30_to_tile_19_29_1),
		.in_wire_0_2(horizontal_tile_19_30_to_tile_19_29_2),
		.in_wire_0_3(horizontal_tile_19_30_to_tile_19_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(638)
	);

	pe_tile pe_tile_19_30(
		.out_wire_3_0(vertical_tile_19_30_to_tile_18_30_0),
		.out_wire_3_1(vertical_tile_19_30_to_tile_18_30_1),
		.out_wire_3_2(vertical_tile_19_30_to_tile_18_30_2),
		.out_wire_3_3(vertical_tile_19_30_to_tile_18_30_3),
		.in_wire_3_0(vertical_tile_18_30_to_tile_19_30_0),
		.in_wire_3_1(vertical_tile_18_30_to_tile_19_30_1),
		.in_wire_3_2(vertical_tile_18_30_to_tile_19_30_2),
		.in_wire_3_3(vertical_tile_18_30_to_tile_19_30_3),
		.out_wire_1_0(vertical_tile_19_30_to_tile_20_30_0),
		.out_wire_1_1(vertical_tile_19_30_to_tile_20_30_1),
		.out_wire_1_2(vertical_tile_19_30_to_tile_20_30_2),
		.out_wire_1_3(vertical_tile_19_30_to_tile_20_30_3),
		.in_wire_1_0(vertical_tile_20_30_to_tile_19_30_0),
		.in_wire_1_1(vertical_tile_20_30_to_tile_19_30_1),
		.in_wire_1_2(vertical_tile_20_30_to_tile_19_30_2),
		.in_wire_1_3(vertical_tile_20_30_to_tile_19_30_3),
		.out_wire_2_0(horizontal_tile_19_30_to_tile_19_29_0),
		.out_wire_2_1(horizontal_tile_19_30_to_tile_19_29_1),
		.out_wire_2_2(horizontal_tile_19_30_to_tile_19_29_2),
		.out_wire_2_3(horizontal_tile_19_30_to_tile_19_29_3),
		.in_wire_2_0(horizontal_tile_19_29_to_tile_19_30_0),
		.in_wire_2_1(horizontal_tile_19_29_to_tile_19_30_1),
		.in_wire_2_2(horizontal_tile_19_29_to_tile_19_30_2),
		.in_wire_2_3(horizontal_tile_19_29_to_tile_19_30_3),
		.out_wire_0_0(horizontal_tile_19_30_to_tile_19_31_0),
		.out_wire_0_1(horizontal_tile_19_30_to_tile_19_31_1),
		.out_wire_0_2(horizontal_tile_19_30_to_tile_19_31_2),
		.out_wire_0_3(horizontal_tile_19_30_to_tile_19_31_3),
		.in_wire_0_0(horizontal_tile_19_31_to_tile_19_30_0),
		.in_wire_0_1(horizontal_tile_19_31_to_tile_19_30_1),
		.in_wire_0_2(horizontal_tile_19_31_to_tile_19_30_2),
		.in_wire_0_3(horizontal_tile_19_31_to_tile_19_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(639)
	);

	pe_tile_right pe_tile_19_31(
		.out_wire_3_0(vertical_tile_19_31_to_tile_18_31_0),
		.out_wire_3_1(vertical_tile_19_31_to_tile_18_31_1),
		.out_wire_3_2(vertical_tile_19_31_to_tile_18_31_2),
		.out_wire_3_3(vertical_tile_19_31_to_tile_18_31_3),
		.in_wire_3_0(vertical_tile_18_31_to_tile_19_31_0),
		.in_wire_3_1(vertical_tile_18_31_to_tile_19_31_1),
		.in_wire_3_2(vertical_tile_18_31_to_tile_19_31_2),
		.in_wire_3_3(vertical_tile_18_31_to_tile_19_31_3),
		.out_wire_1_0(vertical_tile_19_31_to_tile_20_31_0),
		.out_wire_1_1(vertical_tile_19_31_to_tile_20_31_1),
		.out_wire_1_2(vertical_tile_19_31_to_tile_20_31_2),
		.out_wire_1_3(vertical_tile_19_31_to_tile_20_31_3),
		.in_wire_1_0(vertical_tile_20_31_to_tile_19_31_0),
		.in_wire_1_1(vertical_tile_20_31_to_tile_19_31_1),
		.in_wire_1_2(vertical_tile_20_31_to_tile_19_31_2),
		.in_wire_1_3(vertical_tile_20_31_to_tile_19_31_3),
		.out_wire_2_0(horizontal_tile_19_31_to_tile_19_30_0),
		.out_wire_2_1(horizontal_tile_19_31_to_tile_19_30_1),
		.out_wire_2_2(horizontal_tile_19_31_to_tile_19_30_2),
		.out_wire_2_3(horizontal_tile_19_31_to_tile_19_30_3),
		.in_wire_2_0(horizontal_tile_19_30_to_tile_19_31_0),
		.in_wire_2_1(horizontal_tile_19_30_to_tile_19_31_1),
		.in_wire_2_2(horizontal_tile_19_30_to_tile_19_31_2),
		.in_wire_2_3(horizontal_tile_19_30_to_tile_19_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(640)
	);

	pe_tile_left pe_tile_20_0(
		.out_wire_3_0(vertical_tile_20_0_to_tile_19_0_0),
		.out_wire_3_1(vertical_tile_20_0_to_tile_19_0_1),
		.out_wire_3_2(vertical_tile_20_0_to_tile_19_0_2),
		.out_wire_3_3(vertical_tile_20_0_to_tile_19_0_3),
		.in_wire_3_0(vertical_tile_19_0_to_tile_20_0_0),
		.in_wire_3_1(vertical_tile_19_0_to_tile_20_0_1),
		.in_wire_3_2(vertical_tile_19_0_to_tile_20_0_2),
		.in_wire_3_3(vertical_tile_19_0_to_tile_20_0_3),
		.out_wire_1_0(vertical_tile_20_0_to_tile_21_0_0),
		.out_wire_1_1(vertical_tile_20_0_to_tile_21_0_1),
		.out_wire_1_2(vertical_tile_20_0_to_tile_21_0_2),
		.out_wire_1_3(vertical_tile_20_0_to_tile_21_0_3),
		.in_wire_1_0(vertical_tile_21_0_to_tile_20_0_0),
		.in_wire_1_1(vertical_tile_21_0_to_tile_20_0_1),
		.in_wire_1_2(vertical_tile_21_0_to_tile_20_0_2),
		.in_wire_1_3(vertical_tile_21_0_to_tile_20_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_20_0_to_tile_20_1_0),
		.out_wire_0_1(horizontal_tile_20_0_to_tile_20_1_1),
		.out_wire_0_2(horizontal_tile_20_0_to_tile_20_1_2),
		.out_wire_0_3(horizontal_tile_20_0_to_tile_20_1_3),
		.in_wire_0_0(horizontal_tile_20_1_to_tile_20_0_0),
		.in_wire_0_1(horizontal_tile_20_1_to_tile_20_0_1),
		.in_wire_0_2(horizontal_tile_20_1_to_tile_20_0_2),
		.in_wire_0_3(horizontal_tile_20_1_to_tile_20_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(641)
	);

	pe_tile pe_tile_20_1(
		.out_wire_3_0(vertical_tile_20_1_to_tile_19_1_0),
		.out_wire_3_1(vertical_tile_20_1_to_tile_19_1_1),
		.out_wire_3_2(vertical_tile_20_1_to_tile_19_1_2),
		.out_wire_3_3(vertical_tile_20_1_to_tile_19_1_3),
		.in_wire_3_0(vertical_tile_19_1_to_tile_20_1_0),
		.in_wire_3_1(vertical_tile_19_1_to_tile_20_1_1),
		.in_wire_3_2(vertical_tile_19_1_to_tile_20_1_2),
		.in_wire_3_3(vertical_tile_19_1_to_tile_20_1_3),
		.out_wire_1_0(vertical_tile_20_1_to_tile_21_1_0),
		.out_wire_1_1(vertical_tile_20_1_to_tile_21_1_1),
		.out_wire_1_2(vertical_tile_20_1_to_tile_21_1_2),
		.out_wire_1_3(vertical_tile_20_1_to_tile_21_1_3),
		.in_wire_1_0(vertical_tile_21_1_to_tile_20_1_0),
		.in_wire_1_1(vertical_tile_21_1_to_tile_20_1_1),
		.in_wire_1_2(vertical_tile_21_1_to_tile_20_1_2),
		.in_wire_1_3(vertical_tile_21_1_to_tile_20_1_3),
		.out_wire_2_0(horizontal_tile_20_1_to_tile_20_0_0),
		.out_wire_2_1(horizontal_tile_20_1_to_tile_20_0_1),
		.out_wire_2_2(horizontal_tile_20_1_to_tile_20_0_2),
		.out_wire_2_3(horizontal_tile_20_1_to_tile_20_0_3),
		.in_wire_2_0(horizontal_tile_20_0_to_tile_20_1_0),
		.in_wire_2_1(horizontal_tile_20_0_to_tile_20_1_1),
		.in_wire_2_2(horizontal_tile_20_0_to_tile_20_1_2),
		.in_wire_2_3(horizontal_tile_20_0_to_tile_20_1_3),
		.out_wire_0_0(horizontal_tile_20_1_to_tile_20_2_0),
		.out_wire_0_1(horizontal_tile_20_1_to_tile_20_2_1),
		.out_wire_0_2(horizontal_tile_20_1_to_tile_20_2_2),
		.out_wire_0_3(horizontal_tile_20_1_to_tile_20_2_3),
		.in_wire_0_0(horizontal_tile_20_2_to_tile_20_1_0),
		.in_wire_0_1(horizontal_tile_20_2_to_tile_20_1_1),
		.in_wire_0_2(horizontal_tile_20_2_to_tile_20_1_2),
		.in_wire_0_3(horizontal_tile_20_2_to_tile_20_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(642)
	);

	pe_tile pe_tile_20_2(
		.out_wire_3_0(vertical_tile_20_2_to_tile_19_2_0),
		.out_wire_3_1(vertical_tile_20_2_to_tile_19_2_1),
		.out_wire_3_2(vertical_tile_20_2_to_tile_19_2_2),
		.out_wire_3_3(vertical_tile_20_2_to_tile_19_2_3),
		.in_wire_3_0(vertical_tile_19_2_to_tile_20_2_0),
		.in_wire_3_1(vertical_tile_19_2_to_tile_20_2_1),
		.in_wire_3_2(vertical_tile_19_2_to_tile_20_2_2),
		.in_wire_3_3(vertical_tile_19_2_to_tile_20_2_3),
		.out_wire_1_0(vertical_tile_20_2_to_tile_21_2_0),
		.out_wire_1_1(vertical_tile_20_2_to_tile_21_2_1),
		.out_wire_1_2(vertical_tile_20_2_to_tile_21_2_2),
		.out_wire_1_3(vertical_tile_20_2_to_tile_21_2_3),
		.in_wire_1_0(vertical_tile_21_2_to_tile_20_2_0),
		.in_wire_1_1(vertical_tile_21_2_to_tile_20_2_1),
		.in_wire_1_2(vertical_tile_21_2_to_tile_20_2_2),
		.in_wire_1_3(vertical_tile_21_2_to_tile_20_2_3),
		.out_wire_2_0(horizontal_tile_20_2_to_tile_20_1_0),
		.out_wire_2_1(horizontal_tile_20_2_to_tile_20_1_1),
		.out_wire_2_2(horizontal_tile_20_2_to_tile_20_1_2),
		.out_wire_2_3(horizontal_tile_20_2_to_tile_20_1_3),
		.in_wire_2_0(horizontal_tile_20_1_to_tile_20_2_0),
		.in_wire_2_1(horizontal_tile_20_1_to_tile_20_2_1),
		.in_wire_2_2(horizontal_tile_20_1_to_tile_20_2_2),
		.in_wire_2_3(horizontal_tile_20_1_to_tile_20_2_3),
		.out_wire_0_0(horizontal_tile_20_2_to_tile_20_3_0),
		.out_wire_0_1(horizontal_tile_20_2_to_tile_20_3_1),
		.out_wire_0_2(horizontal_tile_20_2_to_tile_20_3_2),
		.out_wire_0_3(horizontal_tile_20_2_to_tile_20_3_3),
		.in_wire_0_0(horizontal_tile_20_3_to_tile_20_2_0),
		.in_wire_0_1(horizontal_tile_20_3_to_tile_20_2_1),
		.in_wire_0_2(horizontal_tile_20_3_to_tile_20_2_2),
		.in_wire_0_3(horizontal_tile_20_3_to_tile_20_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(643)
	);

	pe_tile pe_tile_20_3(
		.out_wire_3_0(vertical_tile_20_3_to_tile_19_3_0),
		.out_wire_3_1(vertical_tile_20_3_to_tile_19_3_1),
		.out_wire_3_2(vertical_tile_20_3_to_tile_19_3_2),
		.out_wire_3_3(vertical_tile_20_3_to_tile_19_3_3),
		.in_wire_3_0(vertical_tile_19_3_to_tile_20_3_0),
		.in_wire_3_1(vertical_tile_19_3_to_tile_20_3_1),
		.in_wire_3_2(vertical_tile_19_3_to_tile_20_3_2),
		.in_wire_3_3(vertical_tile_19_3_to_tile_20_3_3),
		.out_wire_1_0(vertical_tile_20_3_to_tile_21_3_0),
		.out_wire_1_1(vertical_tile_20_3_to_tile_21_3_1),
		.out_wire_1_2(vertical_tile_20_3_to_tile_21_3_2),
		.out_wire_1_3(vertical_tile_20_3_to_tile_21_3_3),
		.in_wire_1_0(vertical_tile_21_3_to_tile_20_3_0),
		.in_wire_1_1(vertical_tile_21_3_to_tile_20_3_1),
		.in_wire_1_2(vertical_tile_21_3_to_tile_20_3_2),
		.in_wire_1_3(vertical_tile_21_3_to_tile_20_3_3),
		.out_wire_2_0(horizontal_tile_20_3_to_tile_20_2_0),
		.out_wire_2_1(horizontal_tile_20_3_to_tile_20_2_1),
		.out_wire_2_2(horizontal_tile_20_3_to_tile_20_2_2),
		.out_wire_2_3(horizontal_tile_20_3_to_tile_20_2_3),
		.in_wire_2_0(horizontal_tile_20_2_to_tile_20_3_0),
		.in_wire_2_1(horizontal_tile_20_2_to_tile_20_3_1),
		.in_wire_2_2(horizontal_tile_20_2_to_tile_20_3_2),
		.in_wire_2_3(horizontal_tile_20_2_to_tile_20_3_3),
		.out_wire_0_0(horizontal_tile_20_3_to_tile_20_4_0),
		.out_wire_0_1(horizontal_tile_20_3_to_tile_20_4_1),
		.out_wire_0_2(horizontal_tile_20_3_to_tile_20_4_2),
		.out_wire_0_3(horizontal_tile_20_3_to_tile_20_4_3),
		.in_wire_0_0(horizontal_tile_20_4_to_tile_20_3_0),
		.in_wire_0_1(horizontal_tile_20_4_to_tile_20_3_1),
		.in_wire_0_2(horizontal_tile_20_4_to_tile_20_3_2),
		.in_wire_0_3(horizontal_tile_20_4_to_tile_20_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(644)
	);

	pe_tile pe_tile_20_4(
		.out_wire_3_0(vertical_tile_20_4_to_tile_19_4_0),
		.out_wire_3_1(vertical_tile_20_4_to_tile_19_4_1),
		.out_wire_3_2(vertical_tile_20_4_to_tile_19_4_2),
		.out_wire_3_3(vertical_tile_20_4_to_tile_19_4_3),
		.in_wire_3_0(vertical_tile_19_4_to_tile_20_4_0),
		.in_wire_3_1(vertical_tile_19_4_to_tile_20_4_1),
		.in_wire_3_2(vertical_tile_19_4_to_tile_20_4_2),
		.in_wire_3_3(vertical_tile_19_4_to_tile_20_4_3),
		.out_wire_1_0(vertical_tile_20_4_to_tile_21_4_0),
		.out_wire_1_1(vertical_tile_20_4_to_tile_21_4_1),
		.out_wire_1_2(vertical_tile_20_4_to_tile_21_4_2),
		.out_wire_1_3(vertical_tile_20_4_to_tile_21_4_3),
		.in_wire_1_0(vertical_tile_21_4_to_tile_20_4_0),
		.in_wire_1_1(vertical_tile_21_4_to_tile_20_4_1),
		.in_wire_1_2(vertical_tile_21_4_to_tile_20_4_2),
		.in_wire_1_3(vertical_tile_21_4_to_tile_20_4_3),
		.out_wire_2_0(horizontal_tile_20_4_to_tile_20_3_0),
		.out_wire_2_1(horizontal_tile_20_4_to_tile_20_3_1),
		.out_wire_2_2(horizontal_tile_20_4_to_tile_20_3_2),
		.out_wire_2_3(horizontal_tile_20_4_to_tile_20_3_3),
		.in_wire_2_0(horizontal_tile_20_3_to_tile_20_4_0),
		.in_wire_2_1(horizontal_tile_20_3_to_tile_20_4_1),
		.in_wire_2_2(horizontal_tile_20_3_to_tile_20_4_2),
		.in_wire_2_3(horizontal_tile_20_3_to_tile_20_4_3),
		.out_wire_0_0(horizontal_tile_20_4_to_tile_20_5_0),
		.out_wire_0_1(horizontal_tile_20_4_to_tile_20_5_1),
		.out_wire_0_2(horizontal_tile_20_4_to_tile_20_5_2),
		.out_wire_0_3(horizontal_tile_20_4_to_tile_20_5_3),
		.in_wire_0_0(horizontal_tile_20_5_to_tile_20_4_0),
		.in_wire_0_1(horizontal_tile_20_5_to_tile_20_4_1),
		.in_wire_0_2(horizontal_tile_20_5_to_tile_20_4_2),
		.in_wire_0_3(horizontal_tile_20_5_to_tile_20_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(645)
	);

	pe_tile pe_tile_20_5(
		.out_wire_3_0(vertical_tile_20_5_to_tile_19_5_0),
		.out_wire_3_1(vertical_tile_20_5_to_tile_19_5_1),
		.out_wire_3_2(vertical_tile_20_5_to_tile_19_5_2),
		.out_wire_3_3(vertical_tile_20_5_to_tile_19_5_3),
		.in_wire_3_0(vertical_tile_19_5_to_tile_20_5_0),
		.in_wire_3_1(vertical_tile_19_5_to_tile_20_5_1),
		.in_wire_3_2(vertical_tile_19_5_to_tile_20_5_2),
		.in_wire_3_3(vertical_tile_19_5_to_tile_20_5_3),
		.out_wire_1_0(vertical_tile_20_5_to_tile_21_5_0),
		.out_wire_1_1(vertical_tile_20_5_to_tile_21_5_1),
		.out_wire_1_2(vertical_tile_20_5_to_tile_21_5_2),
		.out_wire_1_3(vertical_tile_20_5_to_tile_21_5_3),
		.in_wire_1_0(vertical_tile_21_5_to_tile_20_5_0),
		.in_wire_1_1(vertical_tile_21_5_to_tile_20_5_1),
		.in_wire_1_2(vertical_tile_21_5_to_tile_20_5_2),
		.in_wire_1_3(vertical_tile_21_5_to_tile_20_5_3),
		.out_wire_2_0(horizontal_tile_20_5_to_tile_20_4_0),
		.out_wire_2_1(horizontal_tile_20_5_to_tile_20_4_1),
		.out_wire_2_2(horizontal_tile_20_5_to_tile_20_4_2),
		.out_wire_2_3(horizontal_tile_20_5_to_tile_20_4_3),
		.in_wire_2_0(horizontal_tile_20_4_to_tile_20_5_0),
		.in_wire_2_1(horizontal_tile_20_4_to_tile_20_5_1),
		.in_wire_2_2(horizontal_tile_20_4_to_tile_20_5_2),
		.in_wire_2_3(horizontal_tile_20_4_to_tile_20_5_3),
		.out_wire_0_0(horizontal_tile_20_5_to_tile_20_6_0),
		.out_wire_0_1(horizontal_tile_20_5_to_tile_20_6_1),
		.out_wire_0_2(horizontal_tile_20_5_to_tile_20_6_2),
		.out_wire_0_3(horizontal_tile_20_5_to_tile_20_6_3),
		.in_wire_0_0(horizontal_tile_20_6_to_tile_20_5_0),
		.in_wire_0_1(horizontal_tile_20_6_to_tile_20_5_1),
		.in_wire_0_2(horizontal_tile_20_6_to_tile_20_5_2),
		.in_wire_0_3(horizontal_tile_20_6_to_tile_20_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(646)
	);

	pe_tile pe_tile_20_6(
		.out_wire_3_0(vertical_tile_20_6_to_tile_19_6_0),
		.out_wire_3_1(vertical_tile_20_6_to_tile_19_6_1),
		.out_wire_3_2(vertical_tile_20_6_to_tile_19_6_2),
		.out_wire_3_3(vertical_tile_20_6_to_tile_19_6_3),
		.in_wire_3_0(vertical_tile_19_6_to_tile_20_6_0),
		.in_wire_3_1(vertical_tile_19_6_to_tile_20_6_1),
		.in_wire_3_2(vertical_tile_19_6_to_tile_20_6_2),
		.in_wire_3_3(vertical_tile_19_6_to_tile_20_6_3),
		.out_wire_1_0(vertical_tile_20_6_to_tile_21_6_0),
		.out_wire_1_1(vertical_tile_20_6_to_tile_21_6_1),
		.out_wire_1_2(vertical_tile_20_6_to_tile_21_6_2),
		.out_wire_1_3(vertical_tile_20_6_to_tile_21_6_3),
		.in_wire_1_0(vertical_tile_21_6_to_tile_20_6_0),
		.in_wire_1_1(vertical_tile_21_6_to_tile_20_6_1),
		.in_wire_1_2(vertical_tile_21_6_to_tile_20_6_2),
		.in_wire_1_3(vertical_tile_21_6_to_tile_20_6_3),
		.out_wire_2_0(horizontal_tile_20_6_to_tile_20_5_0),
		.out_wire_2_1(horizontal_tile_20_6_to_tile_20_5_1),
		.out_wire_2_2(horizontal_tile_20_6_to_tile_20_5_2),
		.out_wire_2_3(horizontal_tile_20_6_to_tile_20_5_3),
		.in_wire_2_0(horizontal_tile_20_5_to_tile_20_6_0),
		.in_wire_2_1(horizontal_tile_20_5_to_tile_20_6_1),
		.in_wire_2_2(horizontal_tile_20_5_to_tile_20_6_2),
		.in_wire_2_3(horizontal_tile_20_5_to_tile_20_6_3),
		.out_wire_0_0(horizontal_tile_20_6_to_tile_20_7_0),
		.out_wire_0_1(horizontal_tile_20_6_to_tile_20_7_1),
		.out_wire_0_2(horizontal_tile_20_6_to_tile_20_7_2),
		.out_wire_0_3(horizontal_tile_20_6_to_tile_20_7_3),
		.in_wire_0_0(horizontal_tile_20_7_to_tile_20_6_0),
		.in_wire_0_1(horizontal_tile_20_7_to_tile_20_6_1),
		.in_wire_0_2(horizontal_tile_20_7_to_tile_20_6_2),
		.in_wire_0_3(horizontal_tile_20_7_to_tile_20_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(647)
	);

	pe_tile pe_tile_20_7(
		.out_wire_3_0(vertical_tile_20_7_to_tile_19_7_0),
		.out_wire_3_1(vertical_tile_20_7_to_tile_19_7_1),
		.out_wire_3_2(vertical_tile_20_7_to_tile_19_7_2),
		.out_wire_3_3(vertical_tile_20_7_to_tile_19_7_3),
		.in_wire_3_0(vertical_tile_19_7_to_tile_20_7_0),
		.in_wire_3_1(vertical_tile_19_7_to_tile_20_7_1),
		.in_wire_3_2(vertical_tile_19_7_to_tile_20_7_2),
		.in_wire_3_3(vertical_tile_19_7_to_tile_20_7_3),
		.out_wire_1_0(vertical_tile_20_7_to_tile_21_7_0),
		.out_wire_1_1(vertical_tile_20_7_to_tile_21_7_1),
		.out_wire_1_2(vertical_tile_20_7_to_tile_21_7_2),
		.out_wire_1_3(vertical_tile_20_7_to_tile_21_7_3),
		.in_wire_1_0(vertical_tile_21_7_to_tile_20_7_0),
		.in_wire_1_1(vertical_tile_21_7_to_tile_20_7_1),
		.in_wire_1_2(vertical_tile_21_7_to_tile_20_7_2),
		.in_wire_1_3(vertical_tile_21_7_to_tile_20_7_3),
		.out_wire_2_0(horizontal_tile_20_7_to_tile_20_6_0),
		.out_wire_2_1(horizontal_tile_20_7_to_tile_20_6_1),
		.out_wire_2_2(horizontal_tile_20_7_to_tile_20_6_2),
		.out_wire_2_3(horizontal_tile_20_7_to_tile_20_6_3),
		.in_wire_2_0(horizontal_tile_20_6_to_tile_20_7_0),
		.in_wire_2_1(horizontal_tile_20_6_to_tile_20_7_1),
		.in_wire_2_2(horizontal_tile_20_6_to_tile_20_7_2),
		.in_wire_2_3(horizontal_tile_20_6_to_tile_20_7_3),
		.out_wire_0_0(horizontal_tile_20_7_to_tile_20_8_0),
		.out_wire_0_1(horizontal_tile_20_7_to_tile_20_8_1),
		.out_wire_0_2(horizontal_tile_20_7_to_tile_20_8_2),
		.out_wire_0_3(horizontal_tile_20_7_to_tile_20_8_3),
		.in_wire_0_0(horizontal_tile_20_8_to_tile_20_7_0),
		.in_wire_0_1(horizontal_tile_20_8_to_tile_20_7_1),
		.in_wire_0_2(horizontal_tile_20_8_to_tile_20_7_2),
		.in_wire_0_3(horizontal_tile_20_8_to_tile_20_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(648)
	);

	pe_tile pe_tile_20_8(
		.out_wire_3_0(vertical_tile_20_8_to_tile_19_8_0),
		.out_wire_3_1(vertical_tile_20_8_to_tile_19_8_1),
		.out_wire_3_2(vertical_tile_20_8_to_tile_19_8_2),
		.out_wire_3_3(vertical_tile_20_8_to_tile_19_8_3),
		.in_wire_3_0(vertical_tile_19_8_to_tile_20_8_0),
		.in_wire_3_1(vertical_tile_19_8_to_tile_20_8_1),
		.in_wire_3_2(vertical_tile_19_8_to_tile_20_8_2),
		.in_wire_3_3(vertical_tile_19_8_to_tile_20_8_3),
		.out_wire_1_0(vertical_tile_20_8_to_tile_21_8_0),
		.out_wire_1_1(vertical_tile_20_8_to_tile_21_8_1),
		.out_wire_1_2(vertical_tile_20_8_to_tile_21_8_2),
		.out_wire_1_3(vertical_tile_20_8_to_tile_21_8_3),
		.in_wire_1_0(vertical_tile_21_8_to_tile_20_8_0),
		.in_wire_1_1(vertical_tile_21_8_to_tile_20_8_1),
		.in_wire_1_2(vertical_tile_21_8_to_tile_20_8_2),
		.in_wire_1_3(vertical_tile_21_8_to_tile_20_8_3),
		.out_wire_2_0(horizontal_tile_20_8_to_tile_20_7_0),
		.out_wire_2_1(horizontal_tile_20_8_to_tile_20_7_1),
		.out_wire_2_2(horizontal_tile_20_8_to_tile_20_7_2),
		.out_wire_2_3(horizontal_tile_20_8_to_tile_20_7_3),
		.in_wire_2_0(horizontal_tile_20_7_to_tile_20_8_0),
		.in_wire_2_1(horizontal_tile_20_7_to_tile_20_8_1),
		.in_wire_2_2(horizontal_tile_20_7_to_tile_20_8_2),
		.in_wire_2_3(horizontal_tile_20_7_to_tile_20_8_3),
		.out_wire_0_0(horizontal_tile_20_8_to_tile_20_9_0),
		.out_wire_0_1(horizontal_tile_20_8_to_tile_20_9_1),
		.out_wire_0_2(horizontal_tile_20_8_to_tile_20_9_2),
		.out_wire_0_3(horizontal_tile_20_8_to_tile_20_9_3),
		.in_wire_0_0(horizontal_tile_20_9_to_tile_20_8_0),
		.in_wire_0_1(horizontal_tile_20_9_to_tile_20_8_1),
		.in_wire_0_2(horizontal_tile_20_9_to_tile_20_8_2),
		.in_wire_0_3(horizontal_tile_20_9_to_tile_20_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(649)
	);

	pe_tile pe_tile_20_9(
		.out_wire_3_0(vertical_tile_20_9_to_tile_19_9_0),
		.out_wire_3_1(vertical_tile_20_9_to_tile_19_9_1),
		.out_wire_3_2(vertical_tile_20_9_to_tile_19_9_2),
		.out_wire_3_3(vertical_tile_20_9_to_tile_19_9_3),
		.in_wire_3_0(vertical_tile_19_9_to_tile_20_9_0),
		.in_wire_3_1(vertical_tile_19_9_to_tile_20_9_1),
		.in_wire_3_2(vertical_tile_19_9_to_tile_20_9_2),
		.in_wire_3_3(vertical_tile_19_9_to_tile_20_9_3),
		.out_wire_1_0(vertical_tile_20_9_to_tile_21_9_0),
		.out_wire_1_1(vertical_tile_20_9_to_tile_21_9_1),
		.out_wire_1_2(vertical_tile_20_9_to_tile_21_9_2),
		.out_wire_1_3(vertical_tile_20_9_to_tile_21_9_3),
		.in_wire_1_0(vertical_tile_21_9_to_tile_20_9_0),
		.in_wire_1_1(vertical_tile_21_9_to_tile_20_9_1),
		.in_wire_1_2(vertical_tile_21_9_to_tile_20_9_2),
		.in_wire_1_3(vertical_tile_21_9_to_tile_20_9_3),
		.out_wire_2_0(horizontal_tile_20_9_to_tile_20_8_0),
		.out_wire_2_1(horizontal_tile_20_9_to_tile_20_8_1),
		.out_wire_2_2(horizontal_tile_20_9_to_tile_20_8_2),
		.out_wire_2_3(horizontal_tile_20_9_to_tile_20_8_3),
		.in_wire_2_0(horizontal_tile_20_8_to_tile_20_9_0),
		.in_wire_2_1(horizontal_tile_20_8_to_tile_20_9_1),
		.in_wire_2_2(horizontal_tile_20_8_to_tile_20_9_2),
		.in_wire_2_3(horizontal_tile_20_8_to_tile_20_9_3),
		.out_wire_0_0(horizontal_tile_20_9_to_tile_20_10_0),
		.out_wire_0_1(horizontal_tile_20_9_to_tile_20_10_1),
		.out_wire_0_2(horizontal_tile_20_9_to_tile_20_10_2),
		.out_wire_0_3(horizontal_tile_20_9_to_tile_20_10_3),
		.in_wire_0_0(horizontal_tile_20_10_to_tile_20_9_0),
		.in_wire_0_1(horizontal_tile_20_10_to_tile_20_9_1),
		.in_wire_0_2(horizontal_tile_20_10_to_tile_20_9_2),
		.in_wire_0_3(horizontal_tile_20_10_to_tile_20_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(650)
	);

	pe_tile pe_tile_20_10(
		.out_wire_3_0(vertical_tile_20_10_to_tile_19_10_0),
		.out_wire_3_1(vertical_tile_20_10_to_tile_19_10_1),
		.out_wire_3_2(vertical_tile_20_10_to_tile_19_10_2),
		.out_wire_3_3(vertical_tile_20_10_to_tile_19_10_3),
		.in_wire_3_0(vertical_tile_19_10_to_tile_20_10_0),
		.in_wire_3_1(vertical_tile_19_10_to_tile_20_10_1),
		.in_wire_3_2(vertical_tile_19_10_to_tile_20_10_2),
		.in_wire_3_3(vertical_tile_19_10_to_tile_20_10_3),
		.out_wire_1_0(vertical_tile_20_10_to_tile_21_10_0),
		.out_wire_1_1(vertical_tile_20_10_to_tile_21_10_1),
		.out_wire_1_2(vertical_tile_20_10_to_tile_21_10_2),
		.out_wire_1_3(vertical_tile_20_10_to_tile_21_10_3),
		.in_wire_1_0(vertical_tile_21_10_to_tile_20_10_0),
		.in_wire_1_1(vertical_tile_21_10_to_tile_20_10_1),
		.in_wire_1_2(vertical_tile_21_10_to_tile_20_10_2),
		.in_wire_1_3(vertical_tile_21_10_to_tile_20_10_3),
		.out_wire_2_0(horizontal_tile_20_10_to_tile_20_9_0),
		.out_wire_2_1(horizontal_tile_20_10_to_tile_20_9_1),
		.out_wire_2_2(horizontal_tile_20_10_to_tile_20_9_2),
		.out_wire_2_3(horizontal_tile_20_10_to_tile_20_9_3),
		.in_wire_2_0(horizontal_tile_20_9_to_tile_20_10_0),
		.in_wire_2_1(horizontal_tile_20_9_to_tile_20_10_1),
		.in_wire_2_2(horizontal_tile_20_9_to_tile_20_10_2),
		.in_wire_2_3(horizontal_tile_20_9_to_tile_20_10_3),
		.out_wire_0_0(horizontal_tile_20_10_to_tile_20_11_0),
		.out_wire_0_1(horizontal_tile_20_10_to_tile_20_11_1),
		.out_wire_0_2(horizontal_tile_20_10_to_tile_20_11_2),
		.out_wire_0_3(horizontal_tile_20_10_to_tile_20_11_3),
		.in_wire_0_0(horizontal_tile_20_11_to_tile_20_10_0),
		.in_wire_0_1(horizontal_tile_20_11_to_tile_20_10_1),
		.in_wire_0_2(horizontal_tile_20_11_to_tile_20_10_2),
		.in_wire_0_3(horizontal_tile_20_11_to_tile_20_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(651)
	);

	pe_tile pe_tile_20_11(
		.out_wire_3_0(vertical_tile_20_11_to_tile_19_11_0),
		.out_wire_3_1(vertical_tile_20_11_to_tile_19_11_1),
		.out_wire_3_2(vertical_tile_20_11_to_tile_19_11_2),
		.out_wire_3_3(vertical_tile_20_11_to_tile_19_11_3),
		.in_wire_3_0(vertical_tile_19_11_to_tile_20_11_0),
		.in_wire_3_1(vertical_tile_19_11_to_tile_20_11_1),
		.in_wire_3_2(vertical_tile_19_11_to_tile_20_11_2),
		.in_wire_3_3(vertical_tile_19_11_to_tile_20_11_3),
		.out_wire_1_0(vertical_tile_20_11_to_tile_21_11_0),
		.out_wire_1_1(vertical_tile_20_11_to_tile_21_11_1),
		.out_wire_1_2(vertical_tile_20_11_to_tile_21_11_2),
		.out_wire_1_3(vertical_tile_20_11_to_tile_21_11_3),
		.in_wire_1_0(vertical_tile_21_11_to_tile_20_11_0),
		.in_wire_1_1(vertical_tile_21_11_to_tile_20_11_1),
		.in_wire_1_2(vertical_tile_21_11_to_tile_20_11_2),
		.in_wire_1_3(vertical_tile_21_11_to_tile_20_11_3),
		.out_wire_2_0(horizontal_tile_20_11_to_tile_20_10_0),
		.out_wire_2_1(horizontal_tile_20_11_to_tile_20_10_1),
		.out_wire_2_2(horizontal_tile_20_11_to_tile_20_10_2),
		.out_wire_2_3(horizontal_tile_20_11_to_tile_20_10_3),
		.in_wire_2_0(horizontal_tile_20_10_to_tile_20_11_0),
		.in_wire_2_1(horizontal_tile_20_10_to_tile_20_11_1),
		.in_wire_2_2(horizontal_tile_20_10_to_tile_20_11_2),
		.in_wire_2_3(horizontal_tile_20_10_to_tile_20_11_3),
		.out_wire_0_0(horizontal_tile_20_11_to_tile_20_12_0),
		.out_wire_0_1(horizontal_tile_20_11_to_tile_20_12_1),
		.out_wire_0_2(horizontal_tile_20_11_to_tile_20_12_2),
		.out_wire_0_3(horizontal_tile_20_11_to_tile_20_12_3),
		.in_wire_0_0(horizontal_tile_20_12_to_tile_20_11_0),
		.in_wire_0_1(horizontal_tile_20_12_to_tile_20_11_1),
		.in_wire_0_2(horizontal_tile_20_12_to_tile_20_11_2),
		.in_wire_0_3(horizontal_tile_20_12_to_tile_20_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(652)
	);

	pe_tile pe_tile_20_12(
		.out_wire_3_0(vertical_tile_20_12_to_tile_19_12_0),
		.out_wire_3_1(vertical_tile_20_12_to_tile_19_12_1),
		.out_wire_3_2(vertical_tile_20_12_to_tile_19_12_2),
		.out_wire_3_3(vertical_tile_20_12_to_tile_19_12_3),
		.in_wire_3_0(vertical_tile_19_12_to_tile_20_12_0),
		.in_wire_3_1(vertical_tile_19_12_to_tile_20_12_1),
		.in_wire_3_2(vertical_tile_19_12_to_tile_20_12_2),
		.in_wire_3_3(vertical_tile_19_12_to_tile_20_12_3),
		.out_wire_1_0(vertical_tile_20_12_to_tile_21_12_0),
		.out_wire_1_1(vertical_tile_20_12_to_tile_21_12_1),
		.out_wire_1_2(vertical_tile_20_12_to_tile_21_12_2),
		.out_wire_1_3(vertical_tile_20_12_to_tile_21_12_3),
		.in_wire_1_0(vertical_tile_21_12_to_tile_20_12_0),
		.in_wire_1_1(vertical_tile_21_12_to_tile_20_12_1),
		.in_wire_1_2(vertical_tile_21_12_to_tile_20_12_2),
		.in_wire_1_3(vertical_tile_21_12_to_tile_20_12_3),
		.out_wire_2_0(horizontal_tile_20_12_to_tile_20_11_0),
		.out_wire_2_1(horizontal_tile_20_12_to_tile_20_11_1),
		.out_wire_2_2(horizontal_tile_20_12_to_tile_20_11_2),
		.out_wire_2_3(horizontal_tile_20_12_to_tile_20_11_3),
		.in_wire_2_0(horizontal_tile_20_11_to_tile_20_12_0),
		.in_wire_2_1(horizontal_tile_20_11_to_tile_20_12_1),
		.in_wire_2_2(horizontal_tile_20_11_to_tile_20_12_2),
		.in_wire_2_3(horizontal_tile_20_11_to_tile_20_12_3),
		.out_wire_0_0(horizontal_tile_20_12_to_tile_20_13_0),
		.out_wire_0_1(horizontal_tile_20_12_to_tile_20_13_1),
		.out_wire_0_2(horizontal_tile_20_12_to_tile_20_13_2),
		.out_wire_0_3(horizontal_tile_20_12_to_tile_20_13_3),
		.in_wire_0_0(horizontal_tile_20_13_to_tile_20_12_0),
		.in_wire_0_1(horizontal_tile_20_13_to_tile_20_12_1),
		.in_wire_0_2(horizontal_tile_20_13_to_tile_20_12_2),
		.in_wire_0_3(horizontal_tile_20_13_to_tile_20_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(653)
	);

	pe_tile pe_tile_20_13(
		.out_wire_3_0(vertical_tile_20_13_to_tile_19_13_0),
		.out_wire_3_1(vertical_tile_20_13_to_tile_19_13_1),
		.out_wire_3_2(vertical_tile_20_13_to_tile_19_13_2),
		.out_wire_3_3(vertical_tile_20_13_to_tile_19_13_3),
		.in_wire_3_0(vertical_tile_19_13_to_tile_20_13_0),
		.in_wire_3_1(vertical_tile_19_13_to_tile_20_13_1),
		.in_wire_3_2(vertical_tile_19_13_to_tile_20_13_2),
		.in_wire_3_3(vertical_tile_19_13_to_tile_20_13_3),
		.out_wire_1_0(vertical_tile_20_13_to_tile_21_13_0),
		.out_wire_1_1(vertical_tile_20_13_to_tile_21_13_1),
		.out_wire_1_2(vertical_tile_20_13_to_tile_21_13_2),
		.out_wire_1_3(vertical_tile_20_13_to_tile_21_13_3),
		.in_wire_1_0(vertical_tile_21_13_to_tile_20_13_0),
		.in_wire_1_1(vertical_tile_21_13_to_tile_20_13_1),
		.in_wire_1_2(vertical_tile_21_13_to_tile_20_13_2),
		.in_wire_1_3(vertical_tile_21_13_to_tile_20_13_3),
		.out_wire_2_0(horizontal_tile_20_13_to_tile_20_12_0),
		.out_wire_2_1(horizontal_tile_20_13_to_tile_20_12_1),
		.out_wire_2_2(horizontal_tile_20_13_to_tile_20_12_2),
		.out_wire_2_3(horizontal_tile_20_13_to_tile_20_12_3),
		.in_wire_2_0(horizontal_tile_20_12_to_tile_20_13_0),
		.in_wire_2_1(horizontal_tile_20_12_to_tile_20_13_1),
		.in_wire_2_2(horizontal_tile_20_12_to_tile_20_13_2),
		.in_wire_2_3(horizontal_tile_20_12_to_tile_20_13_3),
		.out_wire_0_0(horizontal_tile_20_13_to_tile_20_14_0),
		.out_wire_0_1(horizontal_tile_20_13_to_tile_20_14_1),
		.out_wire_0_2(horizontal_tile_20_13_to_tile_20_14_2),
		.out_wire_0_3(horizontal_tile_20_13_to_tile_20_14_3),
		.in_wire_0_0(horizontal_tile_20_14_to_tile_20_13_0),
		.in_wire_0_1(horizontal_tile_20_14_to_tile_20_13_1),
		.in_wire_0_2(horizontal_tile_20_14_to_tile_20_13_2),
		.in_wire_0_3(horizontal_tile_20_14_to_tile_20_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(654)
	);

	pe_tile pe_tile_20_14(
		.out_wire_3_0(vertical_tile_20_14_to_tile_19_14_0),
		.out_wire_3_1(vertical_tile_20_14_to_tile_19_14_1),
		.out_wire_3_2(vertical_tile_20_14_to_tile_19_14_2),
		.out_wire_3_3(vertical_tile_20_14_to_tile_19_14_3),
		.in_wire_3_0(vertical_tile_19_14_to_tile_20_14_0),
		.in_wire_3_1(vertical_tile_19_14_to_tile_20_14_1),
		.in_wire_3_2(vertical_tile_19_14_to_tile_20_14_2),
		.in_wire_3_3(vertical_tile_19_14_to_tile_20_14_3),
		.out_wire_1_0(vertical_tile_20_14_to_tile_21_14_0),
		.out_wire_1_1(vertical_tile_20_14_to_tile_21_14_1),
		.out_wire_1_2(vertical_tile_20_14_to_tile_21_14_2),
		.out_wire_1_3(vertical_tile_20_14_to_tile_21_14_3),
		.in_wire_1_0(vertical_tile_21_14_to_tile_20_14_0),
		.in_wire_1_1(vertical_tile_21_14_to_tile_20_14_1),
		.in_wire_1_2(vertical_tile_21_14_to_tile_20_14_2),
		.in_wire_1_3(vertical_tile_21_14_to_tile_20_14_3),
		.out_wire_2_0(horizontal_tile_20_14_to_tile_20_13_0),
		.out_wire_2_1(horizontal_tile_20_14_to_tile_20_13_1),
		.out_wire_2_2(horizontal_tile_20_14_to_tile_20_13_2),
		.out_wire_2_3(horizontal_tile_20_14_to_tile_20_13_3),
		.in_wire_2_0(horizontal_tile_20_13_to_tile_20_14_0),
		.in_wire_2_1(horizontal_tile_20_13_to_tile_20_14_1),
		.in_wire_2_2(horizontal_tile_20_13_to_tile_20_14_2),
		.in_wire_2_3(horizontal_tile_20_13_to_tile_20_14_3),
		.out_wire_0_0(horizontal_tile_20_14_to_tile_20_15_0),
		.out_wire_0_1(horizontal_tile_20_14_to_tile_20_15_1),
		.out_wire_0_2(horizontal_tile_20_14_to_tile_20_15_2),
		.out_wire_0_3(horizontal_tile_20_14_to_tile_20_15_3),
		.in_wire_0_0(horizontal_tile_20_15_to_tile_20_14_0),
		.in_wire_0_1(horizontal_tile_20_15_to_tile_20_14_1),
		.in_wire_0_2(horizontal_tile_20_15_to_tile_20_14_2),
		.in_wire_0_3(horizontal_tile_20_15_to_tile_20_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(655)
	);

	pe_tile pe_tile_20_15(
		.out_wire_3_0(vertical_tile_20_15_to_tile_19_15_0),
		.out_wire_3_1(vertical_tile_20_15_to_tile_19_15_1),
		.out_wire_3_2(vertical_tile_20_15_to_tile_19_15_2),
		.out_wire_3_3(vertical_tile_20_15_to_tile_19_15_3),
		.in_wire_3_0(vertical_tile_19_15_to_tile_20_15_0),
		.in_wire_3_1(vertical_tile_19_15_to_tile_20_15_1),
		.in_wire_3_2(vertical_tile_19_15_to_tile_20_15_2),
		.in_wire_3_3(vertical_tile_19_15_to_tile_20_15_3),
		.out_wire_1_0(vertical_tile_20_15_to_tile_21_15_0),
		.out_wire_1_1(vertical_tile_20_15_to_tile_21_15_1),
		.out_wire_1_2(vertical_tile_20_15_to_tile_21_15_2),
		.out_wire_1_3(vertical_tile_20_15_to_tile_21_15_3),
		.in_wire_1_0(vertical_tile_21_15_to_tile_20_15_0),
		.in_wire_1_1(vertical_tile_21_15_to_tile_20_15_1),
		.in_wire_1_2(vertical_tile_21_15_to_tile_20_15_2),
		.in_wire_1_3(vertical_tile_21_15_to_tile_20_15_3),
		.out_wire_2_0(horizontal_tile_20_15_to_tile_20_14_0),
		.out_wire_2_1(horizontal_tile_20_15_to_tile_20_14_1),
		.out_wire_2_2(horizontal_tile_20_15_to_tile_20_14_2),
		.out_wire_2_3(horizontal_tile_20_15_to_tile_20_14_3),
		.in_wire_2_0(horizontal_tile_20_14_to_tile_20_15_0),
		.in_wire_2_1(horizontal_tile_20_14_to_tile_20_15_1),
		.in_wire_2_2(horizontal_tile_20_14_to_tile_20_15_2),
		.in_wire_2_3(horizontal_tile_20_14_to_tile_20_15_3),
		.out_wire_0_0(horizontal_tile_20_15_to_tile_20_16_0),
		.out_wire_0_1(horizontal_tile_20_15_to_tile_20_16_1),
		.out_wire_0_2(horizontal_tile_20_15_to_tile_20_16_2),
		.out_wire_0_3(horizontal_tile_20_15_to_tile_20_16_3),
		.in_wire_0_0(horizontal_tile_20_16_to_tile_20_15_0),
		.in_wire_0_1(horizontal_tile_20_16_to_tile_20_15_1),
		.in_wire_0_2(horizontal_tile_20_16_to_tile_20_15_2),
		.in_wire_0_3(horizontal_tile_20_16_to_tile_20_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(656)
	);

	pe_tile pe_tile_20_16(
		.out_wire_3_0(vertical_tile_20_16_to_tile_19_16_0),
		.out_wire_3_1(vertical_tile_20_16_to_tile_19_16_1),
		.out_wire_3_2(vertical_tile_20_16_to_tile_19_16_2),
		.out_wire_3_3(vertical_tile_20_16_to_tile_19_16_3),
		.in_wire_3_0(vertical_tile_19_16_to_tile_20_16_0),
		.in_wire_3_1(vertical_tile_19_16_to_tile_20_16_1),
		.in_wire_3_2(vertical_tile_19_16_to_tile_20_16_2),
		.in_wire_3_3(vertical_tile_19_16_to_tile_20_16_3),
		.out_wire_1_0(vertical_tile_20_16_to_tile_21_16_0),
		.out_wire_1_1(vertical_tile_20_16_to_tile_21_16_1),
		.out_wire_1_2(vertical_tile_20_16_to_tile_21_16_2),
		.out_wire_1_3(vertical_tile_20_16_to_tile_21_16_3),
		.in_wire_1_0(vertical_tile_21_16_to_tile_20_16_0),
		.in_wire_1_1(vertical_tile_21_16_to_tile_20_16_1),
		.in_wire_1_2(vertical_tile_21_16_to_tile_20_16_2),
		.in_wire_1_3(vertical_tile_21_16_to_tile_20_16_3),
		.out_wire_2_0(horizontal_tile_20_16_to_tile_20_15_0),
		.out_wire_2_1(horizontal_tile_20_16_to_tile_20_15_1),
		.out_wire_2_2(horizontal_tile_20_16_to_tile_20_15_2),
		.out_wire_2_3(horizontal_tile_20_16_to_tile_20_15_3),
		.in_wire_2_0(horizontal_tile_20_15_to_tile_20_16_0),
		.in_wire_2_1(horizontal_tile_20_15_to_tile_20_16_1),
		.in_wire_2_2(horizontal_tile_20_15_to_tile_20_16_2),
		.in_wire_2_3(horizontal_tile_20_15_to_tile_20_16_3),
		.out_wire_0_0(horizontal_tile_20_16_to_tile_20_17_0),
		.out_wire_0_1(horizontal_tile_20_16_to_tile_20_17_1),
		.out_wire_0_2(horizontal_tile_20_16_to_tile_20_17_2),
		.out_wire_0_3(horizontal_tile_20_16_to_tile_20_17_3),
		.in_wire_0_0(horizontal_tile_20_17_to_tile_20_16_0),
		.in_wire_0_1(horizontal_tile_20_17_to_tile_20_16_1),
		.in_wire_0_2(horizontal_tile_20_17_to_tile_20_16_2),
		.in_wire_0_3(horizontal_tile_20_17_to_tile_20_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(657)
	);

	pe_tile pe_tile_20_17(
		.out_wire_3_0(vertical_tile_20_17_to_tile_19_17_0),
		.out_wire_3_1(vertical_tile_20_17_to_tile_19_17_1),
		.out_wire_3_2(vertical_tile_20_17_to_tile_19_17_2),
		.out_wire_3_3(vertical_tile_20_17_to_tile_19_17_3),
		.in_wire_3_0(vertical_tile_19_17_to_tile_20_17_0),
		.in_wire_3_1(vertical_tile_19_17_to_tile_20_17_1),
		.in_wire_3_2(vertical_tile_19_17_to_tile_20_17_2),
		.in_wire_3_3(vertical_tile_19_17_to_tile_20_17_3),
		.out_wire_1_0(vertical_tile_20_17_to_tile_21_17_0),
		.out_wire_1_1(vertical_tile_20_17_to_tile_21_17_1),
		.out_wire_1_2(vertical_tile_20_17_to_tile_21_17_2),
		.out_wire_1_3(vertical_tile_20_17_to_tile_21_17_3),
		.in_wire_1_0(vertical_tile_21_17_to_tile_20_17_0),
		.in_wire_1_1(vertical_tile_21_17_to_tile_20_17_1),
		.in_wire_1_2(vertical_tile_21_17_to_tile_20_17_2),
		.in_wire_1_3(vertical_tile_21_17_to_tile_20_17_3),
		.out_wire_2_0(horizontal_tile_20_17_to_tile_20_16_0),
		.out_wire_2_1(horizontal_tile_20_17_to_tile_20_16_1),
		.out_wire_2_2(horizontal_tile_20_17_to_tile_20_16_2),
		.out_wire_2_3(horizontal_tile_20_17_to_tile_20_16_3),
		.in_wire_2_0(horizontal_tile_20_16_to_tile_20_17_0),
		.in_wire_2_1(horizontal_tile_20_16_to_tile_20_17_1),
		.in_wire_2_2(horizontal_tile_20_16_to_tile_20_17_2),
		.in_wire_2_3(horizontal_tile_20_16_to_tile_20_17_3),
		.out_wire_0_0(horizontal_tile_20_17_to_tile_20_18_0),
		.out_wire_0_1(horizontal_tile_20_17_to_tile_20_18_1),
		.out_wire_0_2(horizontal_tile_20_17_to_tile_20_18_2),
		.out_wire_0_3(horizontal_tile_20_17_to_tile_20_18_3),
		.in_wire_0_0(horizontal_tile_20_18_to_tile_20_17_0),
		.in_wire_0_1(horizontal_tile_20_18_to_tile_20_17_1),
		.in_wire_0_2(horizontal_tile_20_18_to_tile_20_17_2),
		.in_wire_0_3(horizontal_tile_20_18_to_tile_20_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(658)
	);

	pe_tile pe_tile_20_18(
		.out_wire_3_0(vertical_tile_20_18_to_tile_19_18_0),
		.out_wire_3_1(vertical_tile_20_18_to_tile_19_18_1),
		.out_wire_3_2(vertical_tile_20_18_to_tile_19_18_2),
		.out_wire_3_3(vertical_tile_20_18_to_tile_19_18_3),
		.in_wire_3_0(vertical_tile_19_18_to_tile_20_18_0),
		.in_wire_3_1(vertical_tile_19_18_to_tile_20_18_1),
		.in_wire_3_2(vertical_tile_19_18_to_tile_20_18_2),
		.in_wire_3_3(vertical_tile_19_18_to_tile_20_18_3),
		.out_wire_1_0(vertical_tile_20_18_to_tile_21_18_0),
		.out_wire_1_1(vertical_tile_20_18_to_tile_21_18_1),
		.out_wire_1_2(vertical_tile_20_18_to_tile_21_18_2),
		.out_wire_1_3(vertical_tile_20_18_to_tile_21_18_3),
		.in_wire_1_0(vertical_tile_21_18_to_tile_20_18_0),
		.in_wire_1_1(vertical_tile_21_18_to_tile_20_18_1),
		.in_wire_1_2(vertical_tile_21_18_to_tile_20_18_2),
		.in_wire_1_3(vertical_tile_21_18_to_tile_20_18_3),
		.out_wire_2_0(horizontal_tile_20_18_to_tile_20_17_0),
		.out_wire_2_1(horizontal_tile_20_18_to_tile_20_17_1),
		.out_wire_2_2(horizontal_tile_20_18_to_tile_20_17_2),
		.out_wire_2_3(horizontal_tile_20_18_to_tile_20_17_3),
		.in_wire_2_0(horizontal_tile_20_17_to_tile_20_18_0),
		.in_wire_2_1(horizontal_tile_20_17_to_tile_20_18_1),
		.in_wire_2_2(horizontal_tile_20_17_to_tile_20_18_2),
		.in_wire_2_3(horizontal_tile_20_17_to_tile_20_18_3),
		.out_wire_0_0(horizontal_tile_20_18_to_tile_20_19_0),
		.out_wire_0_1(horizontal_tile_20_18_to_tile_20_19_1),
		.out_wire_0_2(horizontal_tile_20_18_to_tile_20_19_2),
		.out_wire_0_3(horizontal_tile_20_18_to_tile_20_19_3),
		.in_wire_0_0(horizontal_tile_20_19_to_tile_20_18_0),
		.in_wire_0_1(horizontal_tile_20_19_to_tile_20_18_1),
		.in_wire_0_2(horizontal_tile_20_19_to_tile_20_18_2),
		.in_wire_0_3(horizontal_tile_20_19_to_tile_20_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(659)
	);

	pe_tile pe_tile_20_19(
		.out_wire_3_0(vertical_tile_20_19_to_tile_19_19_0),
		.out_wire_3_1(vertical_tile_20_19_to_tile_19_19_1),
		.out_wire_3_2(vertical_tile_20_19_to_tile_19_19_2),
		.out_wire_3_3(vertical_tile_20_19_to_tile_19_19_3),
		.in_wire_3_0(vertical_tile_19_19_to_tile_20_19_0),
		.in_wire_3_1(vertical_tile_19_19_to_tile_20_19_1),
		.in_wire_3_2(vertical_tile_19_19_to_tile_20_19_2),
		.in_wire_3_3(vertical_tile_19_19_to_tile_20_19_3),
		.out_wire_1_0(vertical_tile_20_19_to_tile_21_19_0),
		.out_wire_1_1(vertical_tile_20_19_to_tile_21_19_1),
		.out_wire_1_2(vertical_tile_20_19_to_tile_21_19_2),
		.out_wire_1_3(vertical_tile_20_19_to_tile_21_19_3),
		.in_wire_1_0(vertical_tile_21_19_to_tile_20_19_0),
		.in_wire_1_1(vertical_tile_21_19_to_tile_20_19_1),
		.in_wire_1_2(vertical_tile_21_19_to_tile_20_19_2),
		.in_wire_1_3(vertical_tile_21_19_to_tile_20_19_3),
		.out_wire_2_0(horizontal_tile_20_19_to_tile_20_18_0),
		.out_wire_2_1(horizontal_tile_20_19_to_tile_20_18_1),
		.out_wire_2_2(horizontal_tile_20_19_to_tile_20_18_2),
		.out_wire_2_3(horizontal_tile_20_19_to_tile_20_18_3),
		.in_wire_2_0(horizontal_tile_20_18_to_tile_20_19_0),
		.in_wire_2_1(horizontal_tile_20_18_to_tile_20_19_1),
		.in_wire_2_2(horizontal_tile_20_18_to_tile_20_19_2),
		.in_wire_2_3(horizontal_tile_20_18_to_tile_20_19_3),
		.out_wire_0_0(horizontal_tile_20_19_to_tile_20_20_0),
		.out_wire_0_1(horizontal_tile_20_19_to_tile_20_20_1),
		.out_wire_0_2(horizontal_tile_20_19_to_tile_20_20_2),
		.out_wire_0_3(horizontal_tile_20_19_to_tile_20_20_3),
		.in_wire_0_0(horizontal_tile_20_20_to_tile_20_19_0),
		.in_wire_0_1(horizontal_tile_20_20_to_tile_20_19_1),
		.in_wire_0_2(horizontal_tile_20_20_to_tile_20_19_2),
		.in_wire_0_3(horizontal_tile_20_20_to_tile_20_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(660)
	);

	pe_tile pe_tile_20_20(
		.out_wire_3_0(vertical_tile_20_20_to_tile_19_20_0),
		.out_wire_3_1(vertical_tile_20_20_to_tile_19_20_1),
		.out_wire_3_2(vertical_tile_20_20_to_tile_19_20_2),
		.out_wire_3_3(vertical_tile_20_20_to_tile_19_20_3),
		.in_wire_3_0(vertical_tile_19_20_to_tile_20_20_0),
		.in_wire_3_1(vertical_tile_19_20_to_tile_20_20_1),
		.in_wire_3_2(vertical_tile_19_20_to_tile_20_20_2),
		.in_wire_3_3(vertical_tile_19_20_to_tile_20_20_3),
		.out_wire_1_0(vertical_tile_20_20_to_tile_21_20_0),
		.out_wire_1_1(vertical_tile_20_20_to_tile_21_20_1),
		.out_wire_1_2(vertical_tile_20_20_to_tile_21_20_2),
		.out_wire_1_3(vertical_tile_20_20_to_tile_21_20_3),
		.in_wire_1_0(vertical_tile_21_20_to_tile_20_20_0),
		.in_wire_1_1(vertical_tile_21_20_to_tile_20_20_1),
		.in_wire_1_2(vertical_tile_21_20_to_tile_20_20_2),
		.in_wire_1_3(vertical_tile_21_20_to_tile_20_20_3),
		.out_wire_2_0(horizontal_tile_20_20_to_tile_20_19_0),
		.out_wire_2_1(horizontal_tile_20_20_to_tile_20_19_1),
		.out_wire_2_2(horizontal_tile_20_20_to_tile_20_19_2),
		.out_wire_2_3(horizontal_tile_20_20_to_tile_20_19_3),
		.in_wire_2_0(horizontal_tile_20_19_to_tile_20_20_0),
		.in_wire_2_1(horizontal_tile_20_19_to_tile_20_20_1),
		.in_wire_2_2(horizontal_tile_20_19_to_tile_20_20_2),
		.in_wire_2_3(horizontal_tile_20_19_to_tile_20_20_3),
		.out_wire_0_0(horizontal_tile_20_20_to_tile_20_21_0),
		.out_wire_0_1(horizontal_tile_20_20_to_tile_20_21_1),
		.out_wire_0_2(horizontal_tile_20_20_to_tile_20_21_2),
		.out_wire_0_3(horizontal_tile_20_20_to_tile_20_21_3),
		.in_wire_0_0(horizontal_tile_20_21_to_tile_20_20_0),
		.in_wire_0_1(horizontal_tile_20_21_to_tile_20_20_1),
		.in_wire_0_2(horizontal_tile_20_21_to_tile_20_20_2),
		.in_wire_0_3(horizontal_tile_20_21_to_tile_20_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(661)
	);

	pe_tile pe_tile_20_21(
		.out_wire_3_0(vertical_tile_20_21_to_tile_19_21_0),
		.out_wire_3_1(vertical_tile_20_21_to_tile_19_21_1),
		.out_wire_3_2(vertical_tile_20_21_to_tile_19_21_2),
		.out_wire_3_3(vertical_tile_20_21_to_tile_19_21_3),
		.in_wire_3_0(vertical_tile_19_21_to_tile_20_21_0),
		.in_wire_3_1(vertical_tile_19_21_to_tile_20_21_1),
		.in_wire_3_2(vertical_tile_19_21_to_tile_20_21_2),
		.in_wire_3_3(vertical_tile_19_21_to_tile_20_21_3),
		.out_wire_1_0(vertical_tile_20_21_to_tile_21_21_0),
		.out_wire_1_1(vertical_tile_20_21_to_tile_21_21_1),
		.out_wire_1_2(vertical_tile_20_21_to_tile_21_21_2),
		.out_wire_1_3(vertical_tile_20_21_to_tile_21_21_3),
		.in_wire_1_0(vertical_tile_21_21_to_tile_20_21_0),
		.in_wire_1_1(vertical_tile_21_21_to_tile_20_21_1),
		.in_wire_1_2(vertical_tile_21_21_to_tile_20_21_2),
		.in_wire_1_3(vertical_tile_21_21_to_tile_20_21_3),
		.out_wire_2_0(horizontal_tile_20_21_to_tile_20_20_0),
		.out_wire_2_1(horizontal_tile_20_21_to_tile_20_20_1),
		.out_wire_2_2(horizontal_tile_20_21_to_tile_20_20_2),
		.out_wire_2_3(horizontal_tile_20_21_to_tile_20_20_3),
		.in_wire_2_0(horizontal_tile_20_20_to_tile_20_21_0),
		.in_wire_2_1(horizontal_tile_20_20_to_tile_20_21_1),
		.in_wire_2_2(horizontal_tile_20_20_to_tile_20_21_2),
		.in_wire_2_3(horizontal_tile_20_20_to_tile_20_21_3),
		.out_wire_0_0(horizontal_tile_20_21_to_tile_20_22_0),
		.out_wire_0_1(horizontal_tile_20_21_to_tile_20_22_1),
		.out_wire_0_2(horizontal_tile_20_21_to_tile_20_22_2),
		.out_wire_0_3(horizontal_tile_20_21_to_tile_20_22_3),
		.in_wire_0_0(horizontal_tile_20_22_to_tile_20_21_0),
		.in_wire_0_1(horizontal_tile_20_22_to_tile_20_21_1),
		.in_wire_0_2(horizontal_tile_20_22_to_tile_20_21_2),
		.in_wire_0_3(horizontal_tile_20_22_to_tile_20_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(662)
	);

	pe_tile pe_tile_20_22(
		.out_wire_3_0(vertical_tile_20_22_to_tile_19_22_0),
		.out_wire_3_1(vertical_tile_20_22_to_tile_19_22_1),
		.out_wire_3_2(vertical_tile_20_22_to_tile_19_22_2),
		.out_wire_3_3(vertical_tile_20_22_to_tile_19_22_3),
		.in_wire_3_0(vertical_tile_19_22_to_tile_20_22_0),
		.in_wire_3_1(vertical_tile_19_22_to_tile_20_22_1),
		.in_wire_3_2(vertical_tile_19_22_to_tile_20_22_2),
		.in_wire_3_3(vertical_tile_19_22_to_tile_20_22_3),
		.out_wire_1_0(vertical_tile_20_22_to_tile_21_22_0),
		.out_wire_1_1(vertical_tile_20_22_to_tile_21_22_1),
		.out_wire_1_2(vertical_tile_20_22_to_tile_21_22_2),
		.out_wire_1_3(vertical_tile_20_22_to_tile_21_22_3),
		.in_wire_1_0(vertical_tile_21_22_to_tile_20_22_0),
		.in_wire_1_1(vertical_tile_21_22_to_tile_20_22_1),
		.in_wire_1_2(vertical_tile_21_22_to_tile_20_22_2),
		.in_wire_1_3(vertical_tile_21_22_to_tile_20_22_3),
		.out_wire_2_0(horizontal_tile_20_22_to_tile_20_21_0),
		.out_wire_2_1(horizontal_tile_20_22_to_tile_20_21_1),
		.out_wire_2_2(horizontal_tile_20_22_to_tile_20_21_2),
		.out_wire_2_3(horizontal_tile_20_22_to_tile_20_21_3),
		.in_wire_2_0(horizontal_tile_20_21_to_tile_20_22_0),
		.in_wire_2_1(horizontal_tile_20_21_to_tile_20_22_1),
		.in_wire_2_2(horizontal_tile_20_21_to_tile_20_22_2),
		.in_wire_2_3(horizontal_tile_20_21_to_tile_20_22_3),
		.out_wire_0_0(horizontal_tile_20_22_to_tile_20_23_0),
		.out_wire_0_1(horizontal_tile_20_22_to_tile_20_23_1),
		.out_wire_0_2(horizontal_tile_20_22_to_tile_20_23_2),
		.out_wire_0_3(horizontal_tile_20_22_to_tile_20_23_3),
		.in_wire_0_0(horizontal_tile_20_23_to_tile_20_22_0),
		.in_wire_0_1(horizontal_tile_20_23_to_tile_20_22_1),
		.in_wire_0_2(horizontal_tile_20_23_to_tile_20_22_2),
		.in_wire_0_3(horizontal_tile_20_23_to_tile_20_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(663)
	);

	pe_tile pe_tile_20_23(
		.out_wire_3_0(vertical_tile_20_23_to_tile_19_23_0),
		.out_wire_3_1(vertical_tile_20_23_to_tile_19_23_1),
		.out_wire_3_2(vertical_tile_20_23_to_tile_19_23_2),
		.out_wire_3_3(vertical_tile_20_23_to_tile_19_23_3),
		.in_wire_3_0(vertical_tile_19_23_to_tile_20_23_0),
		.in_wire_3_1(vertical_tile_19_23_to_tile_20_23_1),
		.in_wire_3_2(vertical_tile_19_23_to_tile_20_23_2),
		.in_wire_3_3(vertical_tile_19_23_to_tile_20_23_3),
		.out_wire_1_0(vertical_tile_20_23_to_tile_21_23_0),
		.out_wire_1_1(vertical_tile_20_23_to_tile_21_23_1),
		.out_wire_1_2(vertical_tile_20_23_to_tile_21_23_2),
		.out_wire_1_3(vertical_tile_20_23_to_tile_21_23_3),
		.in_wire_1_0(vertical_tile_21_23_to_tile_20_23_0),
		.in_wire_1_1(vertical_tile_21_23_to_tile_20_23_1),
		.in_wire_1_2(vertical_tile_21_23_to_tile_20_23_2),
		.in_wire_1_3(vertical_tile_21_23_to_tile_20_23_3),
		.out_wire_2_0(horizontal_tile_20_23_to_tile_20_22_0),
		.out_wire_2_1(horizontal_tile_20_23_to_tile_20_22_1),
		.out_wire_2_2(horizontal_tile_20_23_to_tile_20_22_2),
		.out_wire_2_3(horizontal_tile_20_23_to_tile_20_22_3),
		.in_wire_2_0(horizontal_tile_20_22_to_tile_20_23_0),
		.in_wire_2_1(horizontal_tile_20_22_to_tile_20_23_1),
		.in_wire_2_2(horizontal_tile_20_22_to_tile_20_23_2),
		.in_wire_2_3(horizontal_tile_20_22_to_tile_20_23_3),
		.out_wire_0_0(horizontal_tile_20_23_to_tile_20_24_0),
		.out_wire_0_1(horizontal_tile_20_23_to_tile_20_24_1),
		.out_wire_0_2(horizontal_tile_20_23_to_tile_20_24_2),
		.out_wire_0_3(horizontal_tile_20_23_to_tile_20_24_3),
		.in_wire_0_0(horizontal_tile_20_24_to_tile_20_23_0),
		.in_wire_0_1(horizontal_tile_20_24_to_tile_20_23_1),
		.in_wire_0_2(horizontal_tile_20_24_to_tile_20_23_2),
		.in_wire_0_3(horizontal_tile_20_24_to_tile_20_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(664)
	);

	pe_tile pe_tile_20_24(
		.out_wire_3_0(vertical_tile_20_24_to_tile_19_24_0),
		.out_wire_3_1(vertical_tile_20_24_to_tile_19_24_1),
		.out_wire_3_2(vertical_tile_20_24_to_tile_19_24_2),
		.out_wire_3_3(vertical_tile_20_24_to_tile_19_24_3),
		.in_wire_3_0(vertical_tile_19_24_to_tile_20_24_0),
		.in_wire_3_1(vertical_tile_19_24_to_tile_20_24_1),
		.in_wire_3_2(vertical_tile_19_24_to_tile_20_24_2),
		.in_wire_3_3(vertical_tile_19_24_to_tile_20_24_3),
		.out_wire_1_0(vertical_tile_20_24_to_tile_21_24_0),
		.out_wire_1_1(vertical_tile_20_24_to_tile_21_24_1),
		.out_wire_1_2(vertical_tile_20_24_to_tile_21_24_2),
		.out_wire_1_3(vertical_tile_20_24_to_tile_21_24_3),
		.in_wire_1_0(vertical_tile_21_24_to_tile_20_24_0),
		.in_wire_1_1(vertical_tile_21_24_to_tile_20_24_1),
		.in_wire_1_2(vertical_tile_21_24_to_tile_20_24_2),
		.in_wire_1_3(vertical_tile_21_24_to_tile_20_24_3),
		.out_wire_2_0(horizontal_tile_20_24_to_tile_20_23_0),
		.out_wire_2_1(horizontal_tile_20_24_to_tile_20_23_1),
		.out_wire_2_2(horizontal_tile_20_24_to_tile_20_23_2),
		.out_wire_2_3(horizontal_tile_20_24_to_tile_20_23_3),
		.in_wire_2_0(horizontal_tile_20_23_to_tile_20_24_0),
		.in_wire_2_1(horizontal_tile_20_23_to_tile_20_24_1),
		.in_wire_2_2(horizontal_tile_20_23_to_tile_20_24_2),
		.in_wire_2_3(horizontal_tile_20_23_to_tile_20_24_3),
		.out_wire_0_0(horizontal_tile_20_24_to_tile_20_25_0),
		.out_wire_0_1(horizontal_tile_20_24_to_tile_20_25_1),
		.out_wire_0_2(horizontal_tile_20_24_to_tile_20_25_2),
		.out_wire_0_3(horizontal_tile_20_24_to_tile_20_25_3),
		.in_wire_0_0(horizontal_tile_20_25_to_tile_20_24_0),
		.in_wire_0_1(horizontal_tile_20_25_to_tile_20_24_1),
		.in_wire_0_2(horizontal_tile_20_25_to_tile_20_24_2),
		.in_wire_0_3(horizontal_tile_20_25_to_tile_20_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(665)
	);

	pe_tile pe_tile_20_25(
		.out_wire_3_0(vertical_tile_20_25_to_tile_19_25_0),
		.out_wire_3_1(vertical_tile_20_25_to_tile_19_25_1),
		.out_wire_3_2(vertical_tile_20_25_to_tile_19_25_2),
		.out_wire_3_3(vertical_tile_20_25_to_tile_19_25_3),
		.in_wire_3_0(vertical_tile_19_25_to_tile_20_25_0),
		.in_wire_3_1(vertical_tile_19_25_to_tile_20_25_1),
		.in_wire_3_2(vertical_tile_19_25_to_tile_20_25_2),
		.in_wire_3_3(vertical_tile_19_25_to_tile_20_25_3),
		.out_wire_1_0(vertical_tile_20_25_to_tile_21_25_0),
		.out_wire_1_1(vertical_tile_20_25_to_tile_21_25_1),
		.out_wire_1_2(vertical_tile_20_25_to_tile_21_25_2),
		.out_wire_1_3(vertical_tile_20_25_to_tile_21_25_3),
		.in_wire_1_0(vertical_tile_21_25_to_tile_20_25_0),
		.in_wire_1_1(vertical_tile_21_25_to_tile_20_25_1),
		.in_wire_1_2(vertical_tile_21_25_to_tile_20_25_2),
		.in_wire_1_3(vertical_tile_21_25_to_tile_20_25_3),
		.out_wire_2_0(horizontal_tile_20_25_to_tile_20_24_0),
		.out_wire_2_1(horizontal_tile_20_25_to_tile_20_24_1),
		.out_wire_2_2(horizontal_tile_20_25_to_tile_20_24_2),
		.out_wire_2_3(horizontal_tile_20_25_to_tile_20_24_3),
		.in_wire_2_0(horizontal_tile_20_24_to_tile_20_25_0),
		.in_wire_2_1(horizontal_tile_20_24_to_tile_20_25_1),
		.in_wire_2_2(horizontal_tile_20_24_to_tile_20_25_2),
		.in_wire_2_3(horizontal_tile_20_24_to_tile_20_25_3),
		.out_wire_0_0(horizontal_tile_20_25_to_tile_20_26_0),
		.out_wire_0_1(horizontal_tile_20_25_to_tile_20_26_1),
		.out_wire_0_2(horizontal_tile_20_25_to_tile_20_26_2),
		.out_wire_0_3(horizontal_tile_20_25_to_tile_20_26_3),
		.in_wire_0_0(horizontal_tile_20_26_to_tile_20_25_0),
		.in_wire_0_1(horizontal_tile_20_26_to_tile_20_25_1),
		.in_wire_0_2(horizontal_tile_20_26_to_tile_20_25_2),
		.in_wire_0_3(horizontal_tile_20_26_to_tile_20_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(666)
	);

	pe_tile pe_tile_20_26(
		.out_wire_3_0(vertical_tile_20_26_to_tile_19_26_0),
		.out_wire_3_1(vertical_tile_20_26_to_tile_19_26_1),
		.out_wire_3_2(vertical_tile_20_26_to_tile_19_26_2),
		.out_wire_3_3(vertical_tile_20_26_to_tile_19_26_3),
		.in_wire_3_0(vertical_tile_19_26_to_tile_20_26_0),
		.in_wire_3_1(vertical_tile_19_26_to_tile_20_26_1),
		.in_wire_3_2(vertical_tile_19_26_to_tile_20_26_2),
		.in_wire_3_3(vertical_tile_19_26_to_tile_20_26_3),
		.out_wire_1_0(vertical_tile_20_26_to_tile_21_26_0),
		.out_wire_1_1(vertical_tile_20_26_to_tile_21_26_1),
		.out_wire_1_2(vertical_tile_20_26_to_tile_21_26_2),
		.out_wire_1_3(vertical_tile_20_26_to_tile_21_26_3),
		.in_wire_1_0(vertical_tile_21_26_to_tile_20_26_0),
		.in_wire_1_1(vertical_tile_21_26_to_tile_20_26_1),
		.in_wire_1_2(vertical_tile_21_26_to_tile_20_26_2),
		.in_wire_1_3(vertical_tile_21_26_to_tile_20_26_3),
		.out_wire_2_0(horizontal_tile_20_26_to_tile_20_25_0),
		.out_wire_2_1(horizontal_tile_20_26_to_tile_20_25_1),
		.out_wire_2_2(horizontal_tile_20_26_to_tile_20_25_2),
		.out_wire_2_3(horizontal_tile_20_26_to_tile_20_25_3),
		.in_wire_2_0(horizontal_tile_20_25_to_tile_20_26_0),
		.in_wire_2_1(horizontal_tile_20_25_to_tile_20_26_1),
		.in_wire_2_2(horizontal_tile_20_25_to_tile_20_26_2),
		.in_wire_2_3(horizontal_tile_20_25_to_tile_20_26_3),
		.out_wire_0_0(horizontal_tile_20_26_to_tile_20_27_0),
		.out_wire_0_1(horizontal_tile_20_26_to_tile_20_27_1),
		.out_wire_0_2(horizontal_tile_20_26_to_tile_20_27_2),
		.out_wire_0_3(horizontal_tile_20_26_to_tile_20_27_3),
		.in_wire_0_0(horizontal_tile_20_27_to_tile_20_26_0),
		.in_wire_0_1(horizontal_tile_20_27_to_tile_20_26_1),
		.in_wire_0_2(horizontal_tile_20_27_to_tile_20_26_2),
		.in_wire_0_3(horizontal_tile_20_27_to_tile_20_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(667)
	);

	pe_tile pe_tile_20_27(
		.out_wire_3_0(vertical_tile_20_27_to_tile_19_27_0),
		.out_wire_3_1(vertical_tile_20_27_to_tile_19_27_1),
		.out_wire_3_2(vertical_tile_20_27_to_tile_19_27_2),
		.out_wire_3_3(vertical_tile_20_27_to_tile_19_27_3),
		.in_wire_3_0(vertical_tile_19_27_to_tile_20_27_0),
		.in_wire_3_1(vertical_tile_19_27_to_tile_20_27_1),
		.in_wire_3_2(vertical_tile_19_27_to_tile_20_27_2),
		.in_wire_3_3(vertical_tile_19_27_to_tile_20_27_3),
		.out_wire_1_0(vertical_tile_20_27_to_tile_21_27_0),
		.out_wire_1_1(vertical_tile_20_27_to_tile_21_27_1),
		.out_wire_1_2(vertical_tile_20_27_to_tile_21_27_2),
		.out_wire_1_3(vertical_tile_20_27_to_tile_21_27_3),
		.in_wire_1_0(vertical_tile_21_27_to_tile_20_27_0),
		.in_wire_1_1(vertical_tile_21_27_to_tile_20_27_1),
		.in_wire_1_2(vertical_tile_21_27_to_tile_20_27_2),
		.in_wire_1_3(vertical_tile_21_27_to_tile_20_27_3),
		.out_wire_2_0(horizontal_tile_20_27_to_tile_20_26_0),
		.out_wire_2_1(horizontal_tile_20_27_to_tile_20_26_1),
		.out_wire_2_2(horizontal_tile_20_27_to_tile_20_26_2),
		.out_wire_2_3(horizontal_tile_20_27_to_tile_20_26_3),
		.in_wire_2_0(horizontal_tile_20_26_to_tile_20_27_0),
		.in_wire_2_1(horizontal_tile_20_26_to_tile_20_27_1),
		.in_wire_2_2(horizontal_tile_20_26_to_tile_20_27_2),
		.in_wire_2_3(horizontal_tile_20_26_to_tile_20_27_3),
		.out_wire_0_0(horizontal_tile_20_27_to_tile_20_28_0),
		.out_wire_0_1(horizontal_tile_20_27_to_tile_20_28_1),
		.out_wire_0_2(horizontal_tile_20_27_to_tile_20_28_2),
		.out_wire_0_3(horizontal_tile_20_27_to_tile_20_28_3),
		.in_wire_0_0(horizontal_tile_20_28_to_tile_20_27_0),
		.in_wire_0_1(horizontal_tile_20_28_to_tile_20_27_1),
		.in_wire_0_2(horizontal_tile_20_28_to_tile_20_27_2),
		.in_wire_0_3(horizontal_tile_20_28_to_tile_20_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(668)
	);

	pe_tile pe_tile_20_28(
		.out_wire_3_0(vertical_tile_20_28_to_tile_19_28_0),
		.out_wire_3_1(vertical_tile_20_28_to_tile_19_28_1),
		.out_wire_3_2(vertical_tile_20_28_to_tile_19_28_2),
		.out_wire_3_3(vertical_tile_20_28_to_tile_19_28_3),
		.in_wire_3_0(vertical_tile_19_28_to_tile_20_28_0),
		.in_wire_3_1(vertical_tile_19_28_to_tile_20_28_1),
		.in_wire_3_2(vertical_tile_19_28_to_tile_20_28_2),
		.in_wire_3_3(vertical_tile_19_28_to_tile_20_28_3),
		.out_wire_1_0(vertical_tile_20_28_to_tile_21_28_0),
		.out_wire_1_1(vertical_tile_20_28_to_tile_21_28_1),
		.out_wire_1_2(vertical_tile_20_28_to_tile_21_28_2),
		.out_wire_1_3(vertical_tile_20_28_to_tile_21_28_3),
		.in_wire_1_0(vertical_tile_21_28_to_tile_20_28_0),
		.in_wire_1_1(vertical_tile_21_28_to_tile_20_28_1),
		.in_wire_1_2(vertical_tile_21_28_to_tile_20_28_2),
		.in_wire_1_3(vertical_tile_21_28_to_tile_20_28_3),
		.out_wire_2_0(horizontal_tile_20_28_to_tile_20_27_0),
		.out_wire_2_1(horizontal_tile_20_28_to_tile_20_27_1),
		.out_wire_2_2(horizontal_tile_20_28_to_tile_20_27_2),
		.out_wire_2_3(horizontal_tile_20_28_to_tile_20_27_3),
		.in_wire_2_0(horizontal_tile_20_27_to_tile_20_28_0),
		.in_wire_2_1(horizontal_tile_20_27_to_tile_20_28_1),
		.in_wire_2_2(horizontal_tile_20_27_to_tile_20_28_2),
		.in_wire_2_3(horizontal_tile_20_27_to_tile_20_28_3),
		.out_wire_0_0(horizontal_tile_20_28_to_tile_20_29_0),
		.out_wire_0_1(horizontal_tile_20_28_to_tile_20_29_1),
		.out_wire_0_2(horizontal_tile_20_28_to_tile_20_29_2),
		.out_wire_0_3(horizontal_tile_20_28_to_tile_20_29_3),
		.in_wire_0_0(horizontal_tile_20_29_to_tile_20_28_0),
		.in_wire_0_1(horizontal_tile_20_29_to_tile_20_28_1),
		.in_wire_0_2(horizontal_tile_20_29_to_tile_20_28_2),
		.in_wire_0_3(horizontal_tile_20_29_to_tile_20_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(669)
	);

	pe_tile pe_tile_20_29(
		.out_wire_3_0(vertical_tile_20_29_to_tile_19_29_0),
		.out_wire_3_1(vertical_tile_20_29_to_tile_19_29_1),
		.out_wire_3_2(vertical_tile_20_29_to_tile_19_29_2),
		.out_wire_3_3(vertical_tile_20_29_to_tile_19_29_3),
		.in_wire_3_0(vertical_tile_19_29_to_tile_20_29_0),
		.in_wire_3_1(vertical_tile_19_29_to_tile_20_29_1),
		.in_wire_3_2(vertical_tile_19_29_to_tile_20_29_2),
		.in_wire_3_3(vertical_tile_19_29_to_tile_20_29_3),
		.out_wire_1_0(vertical_tile_20_29_to_tile_21_29_0),
		.out_wire_1_1(vertical_tile_20_29_to_tile_21_29_1),
		.out_wire_1_2(vertical_tile_20_29_to_tile_21_29_2),
		.out_wire_1_3(vertical_tile_20_29_to_tile_21_29_3),
		.in_wire_1_0(vertical_tile_21_29_to_tile_20_29_0),
		.in_wire_1_1(vertical_tile_21_29_to_tile_20_29_1),
		.in_wire_1_2(vertical_tile_21_29_to_tile_20_29_2),
		.in_wire_1_3(vertical_tile_21_29_to_tile_20_29_3),
		.out_wire_2_0(horizontal_tile_20_29_to_tile_20_28_0),
		.out_wire_2_1(horizontal_tile_20_29_to_tile_20_28_1),
		.out_wire_2_2(horizontal_tile_20_29_to_tile_20_28_2),
		.out_wire_2_3(horizontal_tile_20_29_to_tile_20_28_3),
		.in_wire_2_0(horizontal_tile_20_28_to_tile_20_29_0),
		.in_wire_2_1(horizontal_tile_20_28_to_tile_20_29_1),
		.in_wire_2_2(horizontal_tile_20_28_to_tile_20_29_2),
		.in_wire_2_3(horizontal_tile_20_28_to_tile_20_29_3),
		.out_wire_0_0(horizontal_tile_20_29_to_tile_20_30_0),
		.out_wire_0_1(horizontal_tile_20_29_to_tile_20_30_1),
		.out_wire_0_2(horizontal_tile_20_29_to_tile_20_30_2),
		.out_wire_0_3(horizontal_tile_20_29_to_tile_20_30_3),
		.in_wire_0_0(horizontal_tile_20_30_to_tile_20_29_0),
		.in_wire_0_1(horizontal_tile_20_30_to_tile_20_29_1),
		.in_wire_0_2(horizontal_tile_20_30_to_tile_20_29_2),
		.in_wire_0_3(horizontal_tile_20_30_to_tile_20_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(670)
	);

	pe_tile pe_tile_20_30(
		.out_wire_3_0(vertical_tile_20_30_to_tile_19_30_0),
		.out_wire_3_1(vertical_tile_20_30_to_tile_19_30_1),
		.out_wire_3_2(vertical_tile_20_30_to_tile_19_30_2),
		.out_wire_3_3(vertical_tile_20_30_to_tile_19_30_3),
		.in_wire_3_0(vertical_tile_19_30_to_tile_20_30_0),
		.in_wire_3_1(vertical_tile_19_30_to_tile_20_30_1),
		.in_wire_3_2(vertical_tile_19_30_to_tile_20_30_2),
		.in_wire_3_3(vertical_tile_19_30_to_tile_20_30_3),
		.out_wire_1_0(vertical_tile_20_30_to_tile_21_30_0),
		.out_wire_1_1(vertical_tile_20_30_to_tile_21_30_1),
		.out_wire_1_2(vertical_tile_20_30_to_tile_21_30_2),
		.out_wire_1_3(vertical_tile_20_30_to_tile_21_30_3),
		.in_wire_1_0(vertical_tile_21_30_to_tile_20_30_0),
		.in_wire_1_1(vertical_tile_21_30_to_tile_20_30_1),
		.in_wire_1_2(vertical_tile_21_30_to_tile_20_30_2),
		.in_wire_1_3(vertical_tile_21_30_to_tile_20_30_3),
		.out_wire_2_0(horizontal_tile_20_30_to_tile_20_29_0),
		.out_wire_2_1(horizontal_tile_20_30_to_tile_20_29_1),
		.out_wire_2_2(horizontal_tile_20_30_to_tile_20_29_2),
		.out_wire_2_3(horizontal_tile_20_30_to_tile_20_29_3),
		.in_wire_2_0(horizontal_tile_20_29_to_tile_20_30_0),
		.in_wire_2_1(horizontal_tile_20_29_to_tile_20_30_1),
		.in_wire_2_2(horizontal_tile_20_29_to_tile_20_30_2),
		.in_wire_2_3(horizontal_tile_20_29_to_tile_20_30_3),
		.out_wire_0_0(horizontal_tile_20_30_to_tile_20_31_0),
		.out_wire_0_1(horizontal_tile_20_30_to_tile_20_31_1),
		.out_wire_0_2(horizontal_tile_20_30_to_tile_20_31_2),
		.out_wire_0_3(horizontal_tile_20_30_to_tile_20_31_3),
		.in_wire_0_0(horizontal_tile_20_31_to_tile_20_30_0),
		.in_wire_0_1(horizontal_tile_20_31_to_tile_20_30_1),
		.in_wire_0_2(horizontal_tile_20_31_to_tile_20_30_2),
		.in_wire_0_3(horizontal_tile_20_31_to_tile_20_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(671)
	);

	pe_tile_right pe_tile_20_31(
		.out_wire_3_0(vertical_tile_20_31_to_tile_19_31_0),
		.out_wire_3_1(vertical_tile_20_31_to_tile_19_31_1),
		.out_wire_3_2(vertical_tile_20_31_to_tile_19_31_2),
		.out_wire_3_3(vertical_tile_20_31_to_tile_19_31_3),
		.in_wire_3_0(vertical_tile_19_31_to_tile_20_31_0),
		.in_wire_3_1(vertical_tile_19_31_to_tile_20_31_1),
		.in_wire_3_2(vertical_tile_19_31_to_tile_20_31_2),
		.in_wire_3_3(vertical_tile_19_31_to_tile_20_31_3),
		.out_wire_1_0(vertical_tile_20_31_to_tile_21_31_0),
		.out_wire_1_1(vertical_tile_20_31_to_tile_21_31_1),
		.out_wire_1_2(vertical_tile_20_31_to_tile_21_31_2),
		.out_wire_1_3(vertical_tile_20_31_to_tile_21_31_3),
		.in_wire_1_0(vertical_tile_21_31_to_tile_20_31_0),
		.in_wire_1_1(vertical_tile_21_31_to_tile_20_31_1),
		.in_wire_1_2(vertical_tile_21_31_to_tile_20_31_2),
		.in_wire_1_3(vertical_tile_21_31_to_tile_20_31_3),
		.out_wire_2_0(horizontal_tile_20_31_to_tile_20_30_0),
		.out_wire_2_1(horizontal_tile_20_31_to_tile_20_30_1),
		.out_wire_2_2(horizontal_tile_20_31_to_tile_20_30_2),
		.out_wire_2_3(horizontal_tile_20_31_to_tile_20_30_3),
		.in_wire_2_0(horizontal_tile_20_30_to_tile_20_31_0),
		.in_wire_2_1(horizontal_tile_20_30_to_tile_20_31_1),
		.in_wire_2_2(horizontal_tile_20_30_to_tile_20_31_2),
		.in_wire_2_3(horizontal_tile_20_30_to_tile_20_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(672)
	);

	pe_tile_left pe_tile_21_0(
		.out_wire_3_0(vertical_tile_21_0_to_tile_20_0_0),
		.out_wire_3_1(vertical_tile_21_0_to_tile_20_0_1),
		.out_wire_3_2(vertical_tile_21_0_to_tile_20_0_2),
		.out_wire_3_3(vertical_tile_21_0_to_tile_20_0_3),
		.in_wire_3_0(vertical_tile_20_0_to_tile_21_0_0),
		.in_wire_3_1(vertical_tile_20_0_to_tile_21_0_1),
		.in_wire_3_2(vertical_tile_20_0_to_tile_21_0_2),
		.in_wire_3_3(vertical_tile_20_0_to_tile_21_0_3),
		.out_wire_1_0(vertical_tile_21_0_to_tile_22_0_0),
		.out_wire_1_1(vertical_tile_21_0_to_tile_22_0_1),
		.out_wire_1_2(vertical_tile_21_0_to_tile_22_0_2),
		.out_wire_1_3(vertical_tile_21_0_to_tile_22_0_3),
		.in_wire_1_0(vertical_tile_22_0_to_tile_21_0_0),
		.in_wire_1_1(vertical_tile_22_0_to_tile_21_0_1),
		.in_wire_1_2(vertical_tile_22_0_to_tile_21_0_2),
		.in_wire_1_3(vertical_tile_22_0_to_tile_21_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_21_0_to_tile_21_1_0),
		.out_wire_0_1(horizontal_tile_21_0_to_tile_21_1_1),
		.out_wire_0_2(horizontal_tile_21_0_to_tile_21_1_2),
		.out_wire_0_3(horizontal_tile_21_0_to_tile_21_1_3),
		.in_wire_0_0(horizontal_tile_21_1_to_tile_21_0_0),
		.in_wire_0_1(horizontal_tile_21_1_to_tile_21_0_1),
		.in_wire_0_2(horizontal_tile_21_1_to_tile_21_0_2),
		.in_wire_0_3(horizontal_tile_21_1_to_tile_21_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(673)
	);

	pe_tile pe_tile_21_1(
		.out_wire_3_0(vertical_tile_21_1_to_tile_20_1_0),
		.out_wire_3_1(vertical_tile_21_1_to_tile_20_1_1),
		.out_wire_3_2(vertical_tile_21_1_to_tile_20_1_2),
		.out_wire_3_3(vertical_tile_21_1_to_tile_20_1_3),
		.in_wire_3_0(vertical_tile_20_1_to_tile_21_1_0),
		.in_wire_3_1(vertical_tile_20_1_to_tile_21_1_1),
		.in_wire_3_2(vertical_tile_20_1_to_tile_21_1_2),
		.in_wire_3_3(vertical_tile_20_1_to_tile_21_1_3),
		.out_wire_1_0(vertical_tile_21_1_to_tile_22_1_0),
		.out_wire_1_1(vertical_tile_21_1_to_tile_22_1_1),
		.out_wire_1_2(vertical_tile_21_1_to_tile_22_1_2),
		.out_wire_1_3(vertical_tile_21_1_to_tile_22_1_3),
		.in_wire_1_0(vertical_tile_22_1_to_tile_21_1_0),
		.in_wire_1_1(vertical_tile_22_1_to_tile_21_1_1),
		.in_wire_1_2(vertical_tile_22_1_to_tile_21_1_2),
		.in_wire_1_3(vertical_tile_22_1_to_tile_21_1_3),
		.out_wire_2_0(horizontal_tile_21_1_to_tile_21_0_0),
		.out_wire_2_1(horizontal_tile_21_1_to_tile_21_0_1),
		.out_wire_2_2(horizontal_tile_21_1_to_tile_21_0_2),
		.out_wire_2_3(horizontal_tile_21_1_to_tile_21_0_3),
		.in_wire_2_0(horizontal_tile_21_0_to_tile_21_1_0),
		.in_wire_2_1(horizontal_tile_21_0_to_tile_21_1_1),
		.in_wire_2_2(horizontal_tile_21_0_to_tile_21_1_2),
		.in_wire_2_3(horizontal_tile_21_0_to_tile_21_1_3),
		.out_wire_0_0(horizontal_tile_21_1_to_tile_21_2_0),
		.out_wire_0_1(horizontal_tile_21_1_to_tile_21_2_1),
		.out_wire_0_2(horizontal_tile_21_1_to_tile_21_2_2),
		.out_wire_0_3(horizontal_tile_21_1_to_tile_21_2_3),
		.in_wire_0_0(horizontal_tile_21_2_to_tile_21_1_0),
		.in_wire_0_1(horizontal_tile_21_2_to_tile_21_1_1),
		.in_wire_0_2(horizontal_tile_21_2_to_tile_21_1_2),
		.in_wire_0_3(horizontal_tile_21_2_to_tile_21_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(674)
	);

	pe_tile pe_tile_21_2(
		.out_wire_3_0(vertical_tile_21_2_to_tile_20_2_0),
		.out_wire_3_1(vertical_tile_21_2_to_tile_20_2_1),
		.out_wire_3_2(vertical_tile_21_2_to_tile_20_2_2),
		.out_wire_3_3(vertical_tile_21_2_to_tile_20_2_3),
		.in_wire_3_0(vertical_tile_20_2_to_tile_21_2_0),
		.in_wire_3_1(vertical_tile_20_2_to_tile_21_2_1),
		.in_wire_3_2(vertical_tile_20_2_to_tile_21_2_2),
		.in_wire_3_3(vertical_tile_20_2_to_tile_21_2_3),
		.out_wire_1_0(vertical_tile_21_2_to_tile_22_2_0),
		.out_wire_1_1(vertical_tile_21_2_to_tile_22_2_1),
		.out_wire_1_2(vertical_tile_21_2_to_tile_22_2_2),
		.out_wire_1_3(vertical_tile_21_2_to_tile_22_2_3),
		.in_wire_1_0(vertical_tile_22_2_to_tile_21_2_0),
		.in_wire_1_1(vertical_tile_22_2_to_tile_21_2_1),
		.in_wire_1_2(vertical_tile_22_2_to_tile_21_2_2),
		.in_wire_1_3(vertical_tile_22_2_to_tile_21_2_3),
		.out_wire_2_0(horizontal_tile_21_2_to_tile_21_1_0),
		.out_wire_2_1(horizontal_tile_21_2_to_tile_21_1_1),
		.out_wire_2_2(horizontal_tile_21_2_to_tile_21_1_2),
		.out_wire_2_3(horizontal_tile_21_2_to_tile_21_1_3),
		.in_wire_2_0(horizontal_tile_21_1_to_tile_21_2_0),
		.in_wire_2_1(horizontal_tile_21_1_to_tile_21_2_1),
		.in_wire_2_2(horizontal_tile_21_1_to_tile_21_2_2),
		.in_wire_2_3(horizontal_tile_21_1_to_tile_21_2_3),
		.out_wire_0_0(horizontal_tile_21_2_to_tile_21_3_0),
		.out_wire_0_1(horizontal_tile_21_2_to_tile_21_3_1),
		.out_wire_0_2(horizontal_tile_21_2_to_tile_21_3_2),
		.out_wire_0_3(horizontal_tile_21_2_to_tile_21_3_3),
		.in_wire_0_0(horizontal_tile_21_3_to_tile_21_2_0),
		.in_wire_0_1(horizontal_tile_21_3_to_tile_21_2_1),
		.in_wire_0_2(horizontal_tile_21_3_to_tile_21_2_2),
		.in_wire_0_3(horizontal_tile_21_3_to_tile_21_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(675)
	);

	pe_tile pe_tile_21_3(
		.out_wire_3_0(vertical_tile_21_3_to_tile_20_3_0),
		.out_wire_3_1(vertical_tile_21_3_to_tile_20_3_1),
		.out_wire_3_2(vertical_tile_21_3_to_tile_20_3_2),
		.out_wire_3_3(vertical_tile_21_3_to_tile_20_3_3),
		.in_wire_3_0(vertical_tile_20_3_to_tile_21_3_0),
		.in_wire_3_1(vertical_tile_20_3_to_tile_21_3_1),
		.in_wire_3_2(vertical_tile_20_3_to_tile_21_3_2),
		.in_wire_3_3(vertical_tile_20_3_to_tile_21_3_3),
		.out_wire_1_0(vertical_tile_21_3_to_tile_22_3_0),
		.out_wire_1_1(vertical_tile_21_3_to_tile_22_3_1),
		.out_wire_1_2(vertical_tile_21_3_to_tile_22_3_2),
		.out_wire_1_3(vertical_tile_21_3_to_tile_22_3_3),
		.in_wire_1_0(vertical_tile_22_3_to_tile_21_3_0),
		.in_wire_1_1(vertical_tile_22_3_to_tile_21_3_1),
		.in_wire_1_2(vertical_tile_22_3_to_tile_21_3_2),
		.in_wire_1_3(vertical_tile_22_3_to_tile_21_3_3),
		.out_wire_2_0(horizontal_tile_21_3_to_tile_21_2_0),
		.out_wire_2_1(horizontal_tile_21_3_to_tile_21_2_1),
		.out_wire_2_2(horizontal_tile_21_3_to_tile_21_2_2),
		.out_wire_2_3(horizontal_tile_21_3_to_tile_21_2_3),
		.in_wire_2_0(horizontal_tile_21_2_to_tile_21_3_0),
		.in_wire_2_1(horizontal_tile_21_2_to_tile_21_3_1),
		.in_wire_2_2(horizontal_tile_21_2_to_tile_21_3_2),
		.in_wire_2_3(horizontal_tile_21_2_to_tile_21_3_3),
		.out_wire_0_0(horizontal_tile_21_3_to_tile_21_4_0),
		.out_wire_0_1(horizontal_tile_21_3_to_tile_21_4_1),
		.out_wire_0_2(horizontal_tile_21_3_to_tile_21_4_2),
		.out_wire_0_3(horizontal_tile_21_3_to_tile_21_4_3),
		.in_wire_0_0(horizontal_tile_21_4_to_tile_21_3_0),
		.in_wire_0_1(horizontal_tile_21_4_to_tile_21_3_1),
		.in_wire_0_2(horizontal_tile_21_4_to_tile_21_3_2),
		.in_wire_0_3(horizontal_tile_21_4_to_tile_21_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(676)
	);

	pe_tile pe_tile_21_4(
		.out_wire_3_0(vertical_tile_21_4_to_tile_20_4_0),
		.out_wire_3_1(vertical_tile_21_4_to_tile_20_4_1),
		.out_wire_3_2(vertical_tile_21_4_to_tile_20_4_2),
		.out_wire_3_3(vertical_tile_21_4_to_tile_20_4_3),
		.in_wire_3_0(vertical_tile_20_4_to_tile_21_4_0),
		.in_wire_3_1(vertical_tile_20_4_to_tile_21_4_1),
		.in_wire_3_2(vertical_tile_20_4_to_tile_21_4_2),
		.in_wire_3_3(vertical_tile_20_4_to_tile_21_4_3),
		.out_wire_1_0(vertical_tile_21_4_to_tile_22_4_0),
		.out_wire_1_1(vertical_tile_21_4_to_tile_22_4_1),
		.out_wire_1_2(vertical_tile_21_4_to_tile_22_4_2),
		.out_wire_1_3(vertical_tile_21_4_to_tile_22_4_3),
		.in_wire_1_0(vertical_tile_22_4_to_tile_21_4_0),
		.in_wire_1_1(vertical_tile_22_4_to_tile_21_4_1),
		.in_wire_1_2(vertical_tile_22_4_to_tile_21_4_2),
		.in_wire_1_3(vertical_tile_22_4_to_tile_21_4_3),
		.out_wire_2_0(horizontal_tile_21_4_to_tile_21_3_0),
		.out_wire_2_1(horizontal_tile_21_4_to_tile_21_3_1),
		.out_wire_2_2(horizontal_tile_21_4_to_tile_21_3_2),
		.out_wire_2_3(horizontal_tile_21_4_to_tile_21_3_3),
		.in_wire_2_0(horizontal_tile_21_3_to_tile_21_4_0),
		.in_wire_2_1(horizontal_tile_21_3_to_tile_21_4_1),
		.in_wire_2_2(horizontal_tile_21_3_to_tile_21_4_2),
		.in_wire_2_3(horizontal_tile_21_3_to_tile_21_4_3),
		.out_wire_0_0(horizontal_tile_21_4_to_tile_21_5_0),
		.out_wire_0_1(horizontal_tile_21_4_to_tile_21_5_1),
		.out_wire_0_2(horizontal_tile_21_4_to_tile_21_5_2),
		.out_wire_0_3(horizontal_tile_21_4_to_tile_21_5_3),
		.in_wire_0_0(horizontal_tile_21_5_to_tile_21_4_0),
		.in_wire_0_1(horizontal_tile_21_5_to_tile_21_4_1),
		.in_wire_0_2(horizontal_tile_21_5_to_tile_21_4_2),
		.in_wire_0_3(horizontal_tile_21_5_to_tile_21_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(677)
	);

	pe_tile pe_tile_21_5(
		.out_wire_3_0(vertical_tile_21_5_to_tile_20_5_0),
		.out_wire_3_1(vertical_tile_21_5_to_tile_20_5_1),
		.out_wire_3_2(vertical_tile_21_5_to_tile_20_5_2),
		.out_wire_3_3(vertical_tile_21_5_to_tile_20_5_3),
		.in_wire_3_0(vertical_tile_20_5_to_tile_21_5_0),
		.in_wire_3_1(vertical_tile_20_5_to_tile_21_5_1),
		.in_wire_3_2(vertical_tile_20_5_to_tile_21_5_2),
		.in_wire_3_3(vertical_tile_20_5_to_tile_21_5_3),
		.out_wire_1_0(vertical_tile_21_5_to_tile_22_5_0),
		.out_wire_1_1(vertical_tile_21_5_to_tile_22_5_1),
		.out_wire_1_2(vertical_tile_21_5_to_tile_22_5_2),
		.out_wire_1_3(vertical_tile_21_5_to_tile_22_5_3),
		.in_wire_1_0(vertical_tile_22_5_to_tile_21_5_0),
		.in_wire_1_1(vertical_tile_22_5_to_tile_21_5_1),
		.in_wire_1_2(vertical_tile_22_5_to_tile_21_5_2),
		.in_wire_1_3(vertical_tile_22_5_to_tile_21_5_3),
		.out_wire_2_0(horizontal_tile_21_5_to_tile_21_4_0),
		.out_wire_2_1(horizontal_tile_21_5_to_tile_21_4_1),
		.out_wire_2_2(horizontal_tile_21_5_to_tile_21_4_2),
		.out_wire_2_3(horizontal_tile_21_5_to_tile_21_4_3),
		.in_wire_2_0(horizontal_tile_21_4_to_tile_21_5_0),
		.in_wire_2_1(horizontal_tile_21_4_to_tile_21_5_1),
		.in_wire_2_2(horizontal_tile_21_4_to_tile_21_5_2),
		.in_wire_2_3(horizontal_tile_21_4_to_tile_21_5_3),
		.out_wire_0_0(horizontal_tile_21_5_to_tile_21_6_0),
		.out_wire_0_1(horizontal_tile_21_5_to_tile_21_6_1),
		.out_wire_0_2(horizontal_tile_21_5_to_tile_21_6_2),
		.out_wire_0_3(horizontal_tile_21_5_to_tile_21_6_3),
		.in_wire_0_0(horizontal_tile_21_6_to_tile_21_5_0),
		.in_wire_0_1(horizontal_tile_21_6_to_tile_21_5_1),
		.in_wire_0_2(horizontal_tile_21_6_to_tile_21_5_2),
		.in_wire_0_3(horizontal_tile_21_6_to_tile_21_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(678)
	);

	pe_tile pe_tile_21_6(
		.out_wire_3_0(vertical_tile_21_6_to_tile_20_6_0),
		.out_wire_3_1(vertical_tile_21_6_to_tile_20_6_1),
		.out_wire_3_2(vertical_tile_21_6_to_tile_20_6_2),
		.out_wire_3_3(vertical_tile_21_6_to_tile_20_6_3),
		.in_wire_3_0(vertical_tile_20_6_to_tile_21_6_0),
		.in_wire_3_1(vertical_tile_20_6_to_tile_21_6_1),
		.in_wire_3_2(vertical_tile_20_6_to_tile_21_6_2),
		.in_wire_3_3(vertical_tile_20_6_to_tile_21_6_3),
		.out_wire_1_0(vertical_tile_21_6_to_tile_22_6_0),
		.out_wire_1_1(vertical_tile_21_6_to_tile_22_6_1),
		.out_wire_1_2(vertical_tile_21_6_to_tile_22_6_2),
		.out_wire_1_3(vertical_tile_21_6_to_tile_22_6_3),
		.in_wire_1_0(vertical_tile_22_6_to_tile_21_6_0),
		.in_wire_1_1(vertical_tile_22_6_to_tile_21_6_1),
		.in_wire_1_2(vertical_tile_22_6_to_tile_21_6_2),
		.in_wire_1_3(vertical_tile_22_6_to_tile_21_6_3),
		.out_wire_2_0(horizontal_tile_21_6_to_tile_21_5_0),
		.out_wire_2_1(horizontal_tile_21_6_to_tile_21_5_1),
		.out_wire_2_2(horizontal_tile_21_6_to_tile_21_5_2),
		.out_wire_2_3(horizontal_tile_21_6_to_tile_21_5_3),
		.in_wire_2_0(horizontal_tile_21_5_to_tile_21_6_0),
		.in_wire_2_1(horizontal_tile_21_5_to_tile_21_6_1),
		.in_wire_2_2(horizontal_tile_21_5_to_tile_21_6_2),
		.in_wire_2_3(horizontal_tile_21_5_to_tile_21_6_3),
		.out_wire_0_0(horizontal_tile_21_6_to_tile_21_7_0),
		.out_wire_0_1(horizontal_tile_21_6_to_tile_21_7_1),
		.out_wire_0_2(horizontal_tile_21_6_to_tile_21_7_2),
		.out_wire_0_3(horizontal_tile_21_6_to_tile_21_7_3),
		.in_wire_0_0(horizontal_tile_21_7_to_tile_21_6_0),
		.in_wire_0_1(horizontal_tile_21_7_to_tile_21_6_1),
		.in_wire_0_2(horizontal_tile_21_7_to_tile_21_6_2),
		.in_wire_0_3(horizontal_tile_21_7_to_tile_21_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(679)
	);

	pe_tile pe_tile_21_7(
		.out_wire_3_0(vertical_tile_21_7_to_tile_20_7_0),
		.out_wire_3_1(vertical_tile_21_7_to_tile_20_7_1),
		.out_wire_3_2(vertical_tile_21_7_to_tile_20_7_2),
		.out_wire_3_3(vertical_tile_21_7_to_tile_20_7_3),
		.in_wire_3_0(vertical_tile_20_7_to_tile_21_7_0),
		.in_wire_3_1(vertical_tile_20_7_to_tile_21_7_1),
		.in_wire_3_2(vertical_tile_20_7_to_tile_21_7_2),
		.in_wire_3_3(vertical_tile_20_7_to_tile_21_7_3),
		.out_wire_1_0(vertical_tile_21_7_to_tile_22_7_0),
		.out_wire_1_1(vertical_tile_21_7_to_tile_22_7_1),
		.out_wire_1_2(vertical_tile_21_7_to_tile_22_7_2),
		.out_wire_1_3(vertical_tile_21_7_to_tile_22_7_3),
		.in_wire_1_0(vertical_tile_22_7_to_tile_21_7_0),
		.in_wire_1_1(vertical_tile_22_7_to_tile_21_7_1),
		.in_wire_1_2(vertical_tile_22_7_to_tile_21_7_2),
		.in_wire_1_3(vertical_tile_22_7_to_tile_21_7_3),
		.out_wire_2_0(horizontal_tile_21_7_to_tile_21_6_0),
		.out_wire_2_1(horizontal_tile_21_7_to_tile_21_6_1),
		.out_wire_2_2(horizontal_tile_21_7_to_tile_21_6_2),
		.out_wire_2_3(horizontal_tile_21_7_to_tile_21_6_3),
		.in_wire_2_0(horizontal_tile_21_6_to_tile_21_7_0),
		.in_wire_2_1(horizontal_tile_21_6_to_tile_21_7_1),
		.in_wire_2_2(horizontal_tile_21_6_to_tile_21_7_2),
		.in_wire_2_3(horizontal_tile_21_6_to_tile_21_7_3),
		.out_wire_0_0(horizontal_tile_21_7_to_tile_21_8_0),
		.out_wire_0_1(horizontal_tile_21_7_to_tile_21_8_1),
		.out_wire_0_2(horizontal_tile_21_7_to_tile_21_8_2),
		.out_wire_0_3(horizontal_tile_21_7_to_tile_21_8_3),
		.in_wire_0_0(horizontal_tile_21_8_to_tile_21_7_0),
		.in_wire_0_1(horizontal_tile_21_8_to_tile_21_7_1),
		.in_wire_0_2(horizontal_tile_21_8_to_tile_21_7_2),
		.in_wire_0_3(horizontal_tile_21_8_to_tile_21_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(680)
	);

	pe_tile pe_tile_21_8(
		.out_wire_3_0(vertical_tile_21_8_to_tile_20_8_0),
		.out_wire_3_1(vertical_tile_21_8_to_tile_20_8_1),
		.out_wire_3_2(vertical_tile_21_8_to_tile_20_8_2),
		.out_wire_3_3(vertical_tile_21_8_to_tile_20_8_3),
		.in_wire_3_0(vertical_tile_20_8_to_tile_21_8_0),
		.in_wire_3_1(vertical_tile_20_8_to_tile_21_8_1),
		.in_wire_3_2(vertical_tile_20_8_to_tile_21_8_2),
		.in_wire_3_3(vertical_tile_20_8_to_tile_21_8_3),
		.out_wire_1_0(vertical_tile_21_8_to_tile_22_8_0),
		.out_wire_1_1(vertical_tile_21_8_to_tile_22_8_1),
		.out_wire_1_2(vertical_tile_21_8_to_tile_22_8_2),
		.out_wire_1_3(vertical_tile_21_8_to_tile_22_8_3),
		.in_wire_1_0(vertical_tile_22_8_to_tile_21_8_0),
		.in_wire_1_1(vertical_tile_22_8_to_tile_21_8_1),
		.in_wire_1_2(vertical_tile_22_8_to_tile_21_8_2),
		.in_wire_1_3(vertical_tile_22_8_to_tile_21_8_3),
		.out_wire_2_0(horizontal_tile_21_8_to_tile_21_7_0),
		.out_wire_2_1(horizontal_tile_21_8_to_tile_21_7_1),
		.out_wire_2_2(horizontal_tile_21_8_to_tile_21_7_2),
		.out_wire_2_3(horizontal_tile_21_8_to_tile_21_7_3),
		.in_wire_2_0(horizontal_tile_21_7_to_tile_21_8_0),
		.in_wire_2_1(horizontal_tile_21_7_to_tile_21_8_1),
		.in_wire_2_2(horizontal_tile_21_7_to_tile_21_8_2),
		.in_wire_2_3(horizontal_tile_21_7_to_tile_21_8_3),
		.out_wire_0_0(horizontal_tile_21_8_to_tile_21_9_0),
		.out_wire_0_1(horizontal_tile_21_8_to_tile_21_9_1),
		.out_wire_0_2(horizontal_tile_21_8_to_tile_21_9_2),
		.out_wire_0_3(horizontal_tile_21_8_to_tile_21_9_3),
		.in_wire_0_0(horizontal_tile_21_9_to_tile_21_8_0),
		.in_wire_0_1(horizontal_tile_21_9_to_tile_21_8_1),
		.in_wire_0_2(horizontal_tile_21_9_to_tile_21_8_2),
		.in_wire_0_3(horizontal_tile_21_9_to_tile_21_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(681)
	);

	pe_tile pe_tile_21_9(
		.out_wire_3_0(vertical_tile_21_9_to_tile_20_9_0),
		.out_wire_3_1(vertical_tile_21_9_to_tile_20_9_1),
		.out_wire_3_2(vertical_tile_21_9_to_tile_20_9_2),
		.out_wire_3_3(vertical_tile_21_9_to_tile_20_9_3),
		.in_wire_3_0(vertical_tile_20_9_to_tile_21_9_0),
		.in_wire_3_1(vertical_tile_20_9_to_tile_21_9_1),
		.in_wire_3_2(vertical_tile_20_9_to_tile_21_9_2),
		.in_wire_3_3(vertical_tile_20_9_to_tile_21_9_3),
		.out_wire_1_0(vertical_tile_21_9_to_tile_22_9_0),
		.out_wire_1_1(vertical_tile_21_9_to_tile_22_9_1),
		.out_wire_1_2(vertical_tile_21_9_to_tile_22_9_2),
		.out_wire_1_3(vertical_tile_21_9_to_tile_22_9_3),
		.in_wire_1_0(vertical_tile_22_9_to_tile_21_9_0),
		.in_wire_1_1(vertical_tile_22_9_to_tile_21_9_1),
		.in_wire_1_2(vertical_tile_22_9_to_tile_21_9_2),
		.in_wire_1_3(vertical_tile_22_9_to_tile_21_9_3),
		.out_wire_2_0(horizontal_tile_21_9_to_tile_21_8_0),
		.out_wire_2_1(horizontal_tile_21_9_to_tile_21_8_1),
		.out_wire_2_2(horizontal_tile_21_9_to_tile_21_8_2),
		.out_wire_2_3(horizontal_tile_21_9_to_tile_21_8_3),
		.in_wire_2_0(horizontal_tile_21_8_to_tile_21_9_0),
		.in_wire_2_1(horizontal_tile_21_8_to_tile_21_9_1),
		.in_wire_2_2(horizontal_tile_21_8_to_tile_21_9_2),
		.in_wire_2_3(horizontal_tile_21_8_to_tile_21_9_3),
		.out_wire_0_0(horizontal_tile_21_9_to_tile_21_10_0),
		.out_wire_0_1(horizontal_tile_21_9_to_tile_21_10_1),
		.out_wire_0_2(horizontal_tile_21_9_to_tile_21_10_2),
		.out_wire_0_3(horizontal_tile_21_9_to_tile_21_10_3),
		.in_wire_0_0(horizontal_tile_21_10_to_tile_21_9_0),
		.in_wire_0_1(horizontal_tile_21_10_to_tile_21_9_1),
		.in_wire_0_2(horizontal_tile_21_10_to_tile_21_9_2),
		.in_wire_0_3(horizontal_tile_21_10_to_tile_21_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(682)
	);

	pe_tile pe_tile_21_10(
		.out_wire_3_0(vertical_tile_21_10_to_tile_20_10_0),
		.out_wire_3_1(vertical_tile_21_10_to_tile_20_10_1),
		.out_wire_3_2(vertical_tile_21_10_to_tile_20_10_2),
		.out_wire_3_3(vertical_tile_21_10_to_tile_20_10_3),
		.in_wire_3_0(vertical_tile_20_10_to_tile_21_10_0),
		.in_wire_3_1(vertical_tile_20_10_to_tile_21_10_1),
		.in_wire_3_2(vertical_tile_20_10_to_tile_21_10_2),
		.in_wire_3_3(vertical_tile_20_10_to_tile_21_10_3),
		.out_wire_1_0(vertical_tile_21_10_to_tile_22_10_0),
		.out_wire_1_1(vertical_tile_21_10_to_tile_22_10_1),
		.out_wire_1_2(vertical_tile_21_10_to_tile_22_10_2),
		.out_wire_1_3(vertical_tile_21_10_to_tile_22_10_3),
		.in_wire_1_0(vertical_tile_22_10_to_tile_21_10_0),
		.in_wire_1_1(vertical_tile_22_10_to_tile_21_10_1),
		.in_wire_1_2(vertical_tile_22_10_to_tile_21_10_2),
		.in_wire_1_3(vertical_tile_22_10_to_tile_21_10_3),
		.out_wire_2_0(horizontal_tile_21_10_to_tile_21_9_0),
		.out_wire_2_1(horizontal_tile_21_10_to_tile_21_9_1),
		.out_wire_2_2(horizontal_tile_21_10_to_tile_21_9_2),
		.out_wire_2_3(horizontal_tile_21_10_to_tile_21_9_3),
		.in_wire_2_0(horizontal_tile_21_9_to_tile_21_10_0),
		.in_wire_2_1(horizontal_tile_21_9_to_tile_21_10_1),
		.in_wire_2_2(horizontal_tile_21_9_to_tile_21_10_2),
		.in_wire_2_3(horizontal_tile_21_9_to_tile_21_10_3),
		.out_wire_0_0(horizontal_tile_21_10_to_tile_21_11_0),
		.out_wire_0_1(horizontal_tile_21_10_to_tile_21_11_1),
		.out_wire_0_2(horizontal_tile_21_10_to_tile_21_11_2),
		.out_wire_0_3(horizontal_tile_21_10_to_tile_21_11_3),
		.in_wire_0_0(horizontal_tile_21_11_to_tile_21_10_0),
		.in_wire_0_1(horizontal_tile_21_11_to_tile_21_10_1),
		.in_wire_0_2(horizontal_tile_21_11_to_tile_21_10_2),
		.in_wire_0_3(horizontal_tile_21_11_to_tile_21_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(683)
	);

	pe_tile pe_tile_21_11(
		.out_wire_3_0(vertical_tile_21_11_to_tile_20_11_0),
		.out_wire_3_1(vertical_tile_21_11_to_tile_20_11_1),
		.out_wire_3_2(vertical_tile_21_11_to_tile_20_11_2),
		.out_wire_3_3(vertical_tile_21_11_to_tile_20_11_3),
		.in_wire_3_0(vertical_tile_20_11_to_tile_21_11_0),
		.in_wire_3_1(vertical_tile_20_11_to_tile_21_11_1),
		.in_wire_3_2(vertical_tile_20_11_to_tile_21_11_2),
		.in_wire_3_3(vertical_tile_20_11_to_tile_21_11_3),
		.out_wire_1_0(vertical_tile_21_11_to_tile_22_11_0),
		.out_wire_1_1(vertical_tile_21_11_to_tile_22_11_1),
		.out_wire_1_2(vertical_tile_21_11_to_tile_22_11_2),
		.out_wire_1_3(vertical_tile_21_11_to_tile_22_11_3),
		.in_wire_1_0(vertical_tile_22_11_to_tile_21_11_0),
		.in_wire_1_1(vertical_tile_22_11_to_tile_21_11_1),
		.in_wire_1_2(vertical_tile_22_11_to_tile_21_11_2),
		.in_wire_1_3(vertical_tile_22_11_to_tile_21_11_3),
		.out_wire_2_0(horizontal_tile_21_11_to_tile_21_10_0),
		.out_wire_2_1(horizontal_tile_21_11_to_tile_21_10_1),
		.out_wire_2_2(horizontal_tile_21_11_to_tile_21_10_2),
		.out_wire_2_3(horizontal_tile_21_11_to_tile_21_10_3),
		.in_wire_2_0(horizontal_tile_21_10_to_tile_21_11_0),
		.in_wire_2_1(horizontal_tile_21_10_to_tile_21_11_1),
		.in_wire_2_2(horizontal_tile_21_10_to_tile_21_11_2),
		.in_wire_2_3(horizontal_tile_21_10_to_tile_21_11_3),
		.out_wire_0_0(horizontal_tile_21_11_to_tile_21_12_0),
		.out_wire_0_1(horizontal_tile_21_11_to_tile_21_12_1),
		.out_wire_0_2(horizontal_tile_21_11_to_tile_21_12_2),
		.out_wire_0_3(horizontal_tile_21_11_to_tile_21_12_3),
		.in_wire_0_0(horizontal_tile_21_12_to_tile_21_11_0),
		.in_wire_0_1(horizontal_tile_21_12_to_tile_21_11_1),
		.in_wire_0_2(horizontal_tile_21_12_to_tile_21_11_2),
		.in_wire_0_3(horizontal_tile_21_12_to_tile_21_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(684)
	);

	pe_tile pe_tile_21_12(
		.out_wire_3_0(vertical_tile_21_12_to_tile_20_12_0),
		.out_wire_3_1(vertical_tile_21_12_to_tile_20_12_1),
		.out_wire_3_2(vertical_tile_21_12_to_tile_20_12_2),
		.out_wire_3_3(vertical_tile_21_12_to_tile_20_12_3),
		.in_wire_3_0(vertical_tile_20_12_to_tile_21_12_0),
		.in_wire_3_1(vertical_tile_20_12_to_tile_21_12_1),
		.in_wire_3_2(vertical_tile_20_12_to_tile_21_12_2),
		.in_wire_3_3(vertical_tile_20_12_to_tile_21_12_3),
		.out_wire_1_0(vertical_tile_21_12_to_tile_22_12_0),
		.out_wire_1_1(vertical_tile_21_12_to_tile_22_12_1),
		.out_wire_1_2(vertical_tile_21_12_to_tile_22_12_2),
		.out_wire_1_3(vertical_tile_21_12_to_tile_22_12_3),
		.in_wire_1_0(vertical_tile_22_12_to_tile_21_12_0),
		.in_wire_1_1(vertical_tile_22_12_to_tile_21_12_1),
		.in_wire_1_2(vertical_tile_22_12_to_tile_21_12_2),
		.in_wire_1_3(vertical_tile_22_12_to_tile_21_12_3),
		.out_wire_2_0(horizontal_tile_21_12_to_tile_21_11_0),
		.out_wire_2_1(horizontal_tile_21_12_to_tile_21_11_1),
		.out_wire_2_2(horizontal_tile_21_12_to_tile_21_11_2),
		.out_wire_2_3(horizontal_tile_21_12_to_tile_21_11_3),
		.in_wire_2_0(horizontal_tile_21_11_to_tile_21_12_0),
		.in_wire_2_1(horizontal_tile_21_11_to_tile_21_12_1),
		.in_wire_2_2(horizontal_tile_21_11_to_tile_21_12_2),
		.in_wire_2_3(horizontal_tile_21_11_to_tile_21_12_3),
		.out_wire_0_0(horizontal_tile_21_12_to_tile_21_13_0),
		.out_wire_0_1(horizontal_tile_21_12_to_tile_21_13_1),
		.out_wire_0_2(horizontal_tile_21_12_to_tile_21_13_2),
		.out_wire_0_3(horizontal_tile_21_12_to_tile_21_13_3),
		.in_wire_0_0(horizontal_tile_21_13_to_tile_21_12_0),
		.in_wire_0_1(horizontal_tile_21_13_to_tile_21_12_1),
		.in_wire_0_2(horizontal_tile_21_13_to_tile_21_12_2),
		.in_wire_0_3(horizontal_tile_21_13_to_tile_21_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(685)
	);

	pe_tile pe_tile_21_13(
		.out_wire_3_0(vertical_tile_21_13_to_tile_20_13_0),
		.out_wire_3_1(vertical_tile_21_13_to_tile_20_13_1),
		.out_wire_3_2(vertical_tile_21_13_to_tile_20_13_2),
		.out_wire_3_3(vertical_tile_21_13_to_tile_20_13_3),
		.in_wire_3_0(vertical_tile_20_13_to_tile_21_13_0),
		.in_wire_3_1(vertical_tile_20_13_to_tile_21_13_1),
		.in_wire_3_2(vertical_tile_20_13_to_tile_21_13_2),
		.in_wire_3_3(vertical_tile_20_13_to_tile_21_13_3),
		.out_wire_1_0(vertical_tile_21_13_to_tile_22_13_0),
		.out_wire_1_1(vertical_tile_21_13_to_tile_22_13_1),
		.out_wire_1_2(vertical_tile_21_13_to_tile_22_13_2),
		.out_wire_1_3(vertical_tile_21_13_to_tile_22_13_3),
		.in_wire_1_0(vertical_tile_22_13_to_tile_21_13_0),
		.in_wire_1_1(vertical_tile_22_13_to_tile_21_13_1),
		.in_wire_1_2(vertical_tile_22_13_to_tile_21_13_2),
		.in_wire_1_3(vertical_tile_22_13_to_tile_21_13_3),
		.out_wire_2_0(horizontal_tile_21_13_to_tile_21_12_0),
		.out_wire_2_1(horizontal_tile_21_13_to_tile_21_12_1),
		.out_wire_2_2(horizontal_tile_21_13_to_tile_21_12_2),
		.out_wire_2_3(horizontal_tile_21_13_to_tile_21_12_3),
		.in_wire_2_0(horizontal_tile_21_12_to_tile_21_13_0),
		.in_wire_2_1(horizontal_tile_21_12_to_tile_21_13_1),
		.in_wire_2_2(horizontal_tile_21_12_to_tile_21_13_2),
		.in_wire_2_3(horizontal_tile_21_12_to_tile_21_13_3),
		.out_wire_0_0(horizontal_tile_21_13_to_tile_21_14_0),
		.out_wire_0_1(horizontal_tile_21_13_to_tile_21_14_1),
		.out_wire_0_2(horizontal_tile_21_13_to_tile_21_14_2),
		.out_wire_0_3(horizontal_tile_21_13_to_tile_21_14_3),
		.in_wire_0_0(horizontal_tile_21_14_to_tile_21_13_0),
		.in_wire_0_1(horizontal_tile_21_14_to_tile_21_13_1),
		.in_wire_0_2(horizontal_tile_21_14_to_tile_21_13_2),
		.in_wire_0_3(horizontal_tile_21_14_to_tile_21_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(686)
	);

	pe_tile pe_tile_21_14(
		.out_wire_3_0(vertical_tile_21_14_to_tile_20_14_0),
		.out_wire_3_1(vertical_tile_21_14_to_tile_20_14_1),
		.out_wire_3_2(vertical_tile_21_14_to_tile_20_14_2),
		.out_wire_3_3(vertical_tile_21_14_to_tile_20_14_3),
		.in_wire_3_0(vertical_tile_20_14_to_tile_21_14_0),
		.in_wire_3_1(vertical_tile_20_14_to_tile_21_14_1),
		.in_wire_3_2(vertical_tile_20_14_to_tile_21_14_2),
		.in_wire_3_3(vertical_tile_20_14_to_tile_21_14_3),
		.out_wire_1_0(vertical_tile_21_14_to_tile_22_14_0),
		.out_wire_1_1(vertical_tile_21_14_to_tile_22_14_1),
		.out_wire_1_2(vertical_tile_21_14_to_tile_22_14_2),
		.out_wire_1_3(vertical_tile_21_14_to_tile_22_14_3),
		.in_wire_1_0(vertical_tile_22_14_to_tile_21_14_0),
		.in_wire_1_1(vertical_tile_22_14_to_tile_21_14_1),
		.in_wire_1_2(vertical_tile_22_14_to_tile_21_14_2),
		.in_wire_1_3(vertical_tile_22_14_to_tile_21_14_3),
		.out_wire_2_0(horizontal_tile_21_14_to_tile_21_13_0),
		.out_wire_2_1(horizontal_tile_21_14_to_tile_21_13_1),
		.out_wire_2_2(horizontal_tile_21_14_to_tile_21_13_2),
		.out_wire_2_3(horizontal_tile_21_14_to_tile_21_13_3),
		.in_wire_2_0(horizontal_tile_21_13_to_tile_21_14_0),
		.in_wire_2_1(horizontal_tile_21_13_to_tile_21_14_1),
		.in_wire_2_2(horizontal_tile_21_13_to_tile_21_14_2),
		.in_wire_2_3(horizontal_tile_21_13_to_tile_21_14_3),
		.out_wire_0_0(horizontal_tile_21_14_to_tile_21_15_0),
		.out_wire_0_1(horizontal_tile_21_14_to_tile_21_15_1),
		.out_wire_0_2(horizontal_tile_21_14_to_tile_21_15_2),
		.out_wire_0_3(horizontal_tile_21_14_to_tile_21_15_3),
		.in_wire_0_0(horizontal_tile_21_15_to_tile_21_14_0),
		.in_wire_0_1(horizontal_tile_21_15_to_tile_21_14_1),
		.in_wire_0_2(horizontal_tile_21_15_to_tile_21_14_2),
		.in_wire_0_3(horizontal_tile_21_15_to_tile_21_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(687)
	);

	pe_tile pe_tile_21_15(
		.out_wire_3_0(vertical_tile_21_15_to_tile_20_15_0),
		.out_wire_3_1(vertical_tile_21_15_to_tile_20_15_1),
		.out_wire_3_2(vertical_tile_21_15_to_tile_20_15_2),
		.out_wire_3_3(vertical_tile_21_15_to_tile_20_15_3),
		.in_wire_3_0(vertical_tile_20_15_to_tile_21_15_0),
		.in_wire_3_1(vertical_tile_20_15_to_tile_21_15_1),
		.in_wire_3_2(vertical_tile_20_15_to_tile_21_15_2),
		.in_wire_3_3(vertical_tile_20_15_to_tile_21_15_3),
		.out_wire_1_0(vertical_tile_21_15_to_tile_22_15_0),
		.out_wire_1_1(vertical_tile_21_15_to_tile_22_15_1),
		.out_wire_1_2(vertical_tile_21_15_to_tile_22_15_2),
		.out_wire_1_3(vertical_tile_21_15_to_tile_22_15_3),
		.in_wire_1_0(vertical_tile_22_15_to_tile_21_15_0),
		.in_wire_1_1(vertical_tile_22_15_to_tile_21_15_1),
		.in_wire_1_2(vertical_tile_22_15_to_tile_21_15_2),
		.in_wire_1_3(vertical_tile_22_15_to_tile_21_15_3),
		.out_wire_2_0(horizontal_tile_21_15_to_tile_21_14_0),
		.out_wire_2_1(horizontal_tile_21_15_to_tile_21_14_1),
		.out_wire_2_2(horizontal_tile_21_15_to_tile_21_14_2),
		.out_wire_2_3(horizontal_tile_21_15_to_tile_21_14_3),
		.in_wire_2_0(horizontal_tile_21_14_to_tile_21_15_0),
		.in_wire_2_1(horizontal_tile_21_14_to_tile_21_15_1),
		.in_wire_2_2(horizontal_tile_21_14_to_tile_21_15_2),
		.in_wire_2_3(horizontal_tile_21_14_to_tile_21_15_3),
		.out_wire_0_0(horizontal_tile_21_15_to_tile_21_16_0),
		.out_wire_0_1(horizontal_tile_21_15_to_tile_21_16_1),
		.out_wire_0_2(horizontal_tile_21_15_to_tile_21_16_2),
		.out_wire_0_3(horizontal_tile_21_15_to_tile_21_16_3),
		.in_wire_0_0(horizontal_tile_21_16_to_tile_21_15_0),
		.in_wire_0_1(horizontal_tile_21_16_to_tile_21_15_1),
		.in_wire_0_2(horizontal_tile_21_16_to_tile_21_15_2),
		.in_wire_0_3(horizontal_tile_21_16_to_tile_21_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(688)
	);

	pe_tile pe_tile_21_16(
		.out_wire_3_0(vertical_tile_21_16_to_tile_20_16_0),
		.out_wire_3_1(vertical_tile_21_16_to_tile_20_16_1),
		.out_wire_3_2(vertical_tile_21_16_to_tile_20_16_2),
		.out_wire_3_3(vertical_tile_21_16_to_tile_20_16_3),
		.in_wire_3_0(vertical_tile_20_16_to_tile_21_16_0),
		.in_wire_3_1(vertical_tile_20_16_to_tile_21_16_1),
		.in_wire_3_2(vertical_tile_20_16_to_tile_21_16_2),
		.in_wire_3_3(vertical_tile_20_16_to_tile_21_16_3),
		.out_wire_1_0(vertical_tile_21_16_to_tile_22_16_0),
		.out_wire_1_1(vertical_tile_21_16_to_tile_22_16_1),
		.out_wire_1_2(vertical_tile_21_16_to_tile_22_16_2),
		.out_wire_1_3(vertical_tile_21_16_to_tile_22_16_3),
		.in_wire_1_0(vertical_tile_22_16_to_tile_21_16_0),
		.in_wire_1_1(vertical_tile_22_16_to_tile_21_16_1),
		.in_wire_1_2(vertical_tile_22_16_to_tile_21_16_2),
		.in_wire_1_3(vertical_tile_22_16_to_tile_21_16_3),
		.out_wire_2_0(horizontal_tile_21_16_to_tile_21_15_0),
		.out_wire_2_1(horizontal_tile_21_16_to_tile_21_15_1),
		.out_wire_2_2(horizontal_tile_21_16_to_tile_21_15_2),
		.out_wire_2_3(horizontal_tile_21_16_to_tile_21_15_3),
		.in_wire_2_0(horizontal_tile_21_15_to_tile_21_16_0),
		.in_wire_2_1(horizontal_tile_21_15_to_tile_21_16_1),
		.in_wire_2_2(horizontal_tile_21_15_to_tile_21_16_2),
		.in_wire_2_3(horizontal_tile_21_15_to_tile_21_16_3),
		.out_wire_0_0(horizontal_tile_21_16_to_tile_21_17_0),
		.out_wire_0_1(horizontal_tile_21_16_to_tile_21_17_1),
		.out_wire_0_2(horizontal_tile_21_16_to_tile_21_17_2),
		.out_wire_0_3(horizontal_tile_21_16_to_tile_21_17_3),
		.in_wire_0_0(horizontal_tile_21_17_to_tile_21_16_0),
		.in_wire_0_1(horizontal_tile_21_17_to_tile_21_16_1),
		.in_wire_0_2(horizontal_tile_21_17_to_tile_21_16_2),
		.in_wire_0_3(horizontal_tile_21_17_to_tile_21_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(689)
	);

	pe_tile pe_tile_21_17(
		.out_wire_3_0(vertical_tile_21_17_to_tile_20_17_0),
		.out_wire_3_1(vertical_tile_21_17_to_tile_20_17_1),
		.out_wire_3_2(vertical_tile_21_17_to_tile_20_17_2),
		.out_wire_3_3(vertical_tile_21_17_to_tile_20_17_3),
		.in_wire_3_0(vertical_tile_20_17_to_tile_21_17_0),
		.in_wire_3_1(vertical_tile_20_17_to_tile_21_17_1),
		.in_wire_3_2(vertical_tile_20_17_to_tile_21_17_2),
		.in_wire_3_3(vertical_tile_20_17_to_tile_21_17_3),
		.out_wire_1_0(vertical_tile_21_17_to_tile_22_17_0),
		.out_wire_1_1(vertical_tile_21_17_to_tile_22_17_1),
		.out_wire_1_2(vertical_tile_21_17_to_tile_22_17_2),
		.out_wire_1_3(vertical_tile_21_17_to_tile_22_17_3),
		.in_wire_1_0(vertical_tile_22_17_to_tile_21_17_0),
		.in_wire_1_1(vertical_tile_22_17_to_tile_21_17_1),
		.in_wire_1_2(vertical_tile_22_17_to_tile_21_17_2),
		.in_wire_1_3(vertical_tile_22_17_to_tile_21_17_3),
		.out_wire_2_0(horizontal_tile_21_17_to_tile_21_16_0),
		.out_wire_2_1(horizontal_tile_21_17_to_tile_21_16_1),
		.out_wire_2_2(horizontal_tile_21_17_to_tile_21_16_2),
		.out_wire_2_3(horizontal_tile_21_17_to_tile_21_16_3),
		.in_wire_2_0(horizontal_tile_21_16_to_tile_21_17_0),
		.in_wire_2_1(horizontal_tile_21_16_to_tile_21_17_1),
		.in_wire_2_2(horizontal_tile_21_16_to_tile_21_17_2),
		.in_wire_2_3(horizontal_tile_21_16_to_tile_21_17_3),
		.out_wire_0_0(horizontal_tile_21_17_to_tile_21_18_0),
		.out_wire_0_1(horizontal_tile_21_17_to_tile_21_18_1),
		.out_wire_0_2(horizontal_tile_21_17_to_tile_21_18_2),
		.out_wire_0_3(horizontal_tile_21_17_to_tile_21_18_3),
		.in_wire_0_0(horizontal_tile_21_18_to_tile_21_17_0),
		.in_wire_0_1(horizontal_tile_21_18_to_tile_21_17_1),
		.in_wire_0_2(horizontal_tile_21_18_to_tile_21_17_2),
		.in_wire_0_3(horizontal_tile_21_18_to_tile_21_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(690)
	);

	pe_tile pe_tile_21_18(
		.out_wire_3_0(vertical_tile_21_18_to_tile_20_18_0),
		.out_wire_3_1(vertical_tile_21_18_to_tile_20_18_1),
		.out_wire_3_2(vertical_tile_21_18_to_tile_20_18_2),
		.out_wire_3_3(vertical_tile_21_18_to_tile_20_18_3),
		.in_wire_3_0(vertical_tile_20_18_to_tile_21_18_0),
		.in_wire_3_1(vertical_tile_20_18_to_tile_21_18_1),
		.in_wire_3_2(vertical_tile_20_18_to_tile_21_18_2),
		.in_wire_3_3(vertical_tile_20_18_to_tile_21_18_3),
		.out_wire_1_0(vertical_tile_21_18_to_tile_22_18_0),
		.out_wire_1_1(vertical_tile_21_18_to_tile_22_18_1),
		.out_wire_1_2(vertical_tile_21_18_to_tile_22_18_2),
		.out_wire_1_3(vertical_tile_21_18_to_tile_22_18_3),
		.in_wire_1_0(vertical_tile_22_18_to_tile_21_18_0),
		.in_wire_1_1(vertical_tile_22_18_to_tile_21_18_1),
		.in_wire_1_2(vertical_tile_22_18_to_tile_21_18_2),
		.in_wire_1_3(vertical_tile_22_18_to_tile_21_18_3),
		.out_wire_2_0(horizontal_tile_21_18_to_tile_21_17_0),
		.out_wire_2_1(horizontal_tile_21_18_to_tile_21_17_1),
		.out_wire_2_2(horizontal_tile_21_18_to_tile_21_17_2),
		.out_wire_2_3(horizontal_tile_21_18_to_tile_21_17_3),
		.in_wire_2_0(horizontal_tile_21_17_to_tile_21_18_0),
		.in_wire_2_1(horizontal_tile_21_17_to_tile_21_18_1),
		.in_wire_2_2(horizontal_tile_21_17_to_tile_21_18_2),
		.in_wire_2_3(horizontal_tile_21_17_to_tile_21_18_3),
		.out_wire_0_0(horizontal_tile_21_18_to_tile_21_19_0),
		.out_wire_0_1(horizontal_tile_21_18_to_tile_21_19_1),
		.out_wire_0_2(horizontal_tile_21_18_to_tile_21_19_2),
		.out_wire_0_3(horizontal_tile_21_18_to_tile_21_19_3),
		.in_wire_0_0(horizontal_tile_21_19_to_tile_21_18_0),
		.in_wire_0_1(horizontal_tile_21_19_to_tile_21_18_1),
		.in_wire_0_2(horizontal_tile_21_19_to_tile_21_18_2),
		.in_wire_0_3(horizontal_tile_21_19_to_tile_21_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(691)
	);

	pe_tile pe_tile_21_19(
		.out_wire_3_0(vertical_tile_21_19_to_tile_20_19_0),
		.out_wire_3_1(vertical_tile_21_19_to_tile_20_19_1),
		.out_wire_3_2(vertical_tile_21_19_to_tile_20_19_2),
		.out_wire_3_3(vertical_tile_21_19_to_tile_20_19_3),
		.in_wire_3_0(vertical_tile_20_19_to_tile_21_19_0),
		.in_wire_3_1(vertical_tile_20_19_to_tile_21_19_1),
		.in_wire_3_2(vertical_tile_20_19_to_tile_21_19_2),
		.in_wire_3_3(vertical_tile_20_19_to_tile_21_19_3),
		.out_wire_1_0(vertical_tile_21_19_to_tile_22_19_0),
		.out_wire_1_1(vertical_tile_21_19_to_tile_22_19_1),
		.out_wire_1_2(vertical_tile_21_19_to_tile_22_19_2),
		.out_wire_1_3(vertical_tile_21_19_to_tile_22_19_3),
		.in_wire_1_0(vertical_tile_22_19_to_tile_21_19_0),
		.in_wire_1_1(vertical_tile_22_19_to_tile_21_19_1),
		.in_wire_1_2(vertical_tile_22_19_to_tile_21_19_2),
		.in_wire_1_3(vertical_tile_22_19_to_tile_21_19_3),
		.out_wire_2_0(horizontal_tile_21_19_to_tile_21_18_0),
		.out_wire_2_1(horizontal_tile_21_19_to_tile_21_18_1),
		.out_wire_2_2(horizontal_tile_21_19_to_tile_21_18_2),
		.out_wire_2_3(horizontal_tile_21_19_to_tile_21_18_3),
		.in_wire_2_0(horizontal_tile_21_18_to_tile_21_19_0),
		.in_wire_2_1(horizontal_tile_21_18_to_tile_21_19_1),
		.in_wire_2_2(horizontal_tile_21_18_to_tile_21_19_2),
		.in_wire_2_3(horizontal_tile_21_18_to_tile_21_19_3),
		.out_wire_0_0(horizontal_tile_21_19_to_tile_21_20_0),
		.out_wire_0_1(horizontal_tile_21_19_to_tile_21_20_1),
		.out_wire_0_2(horizontal_tile_21_19_to_tile_21_20_2),
		.out_wire_0_3(horizontal_tile_21_19_to_tile_21_20_3),
		.in_wire_0_0(horizontal_tile_21_20_to_tile_21_19_0),
		.in_wire_0_1(horizontal_tile_21_20_to_tile_21_19_1),
		.in_wire_0_2(horizontal_tile_21_20_to_tile_21_19_2),
		.in_wire_0_3(horizontal_tile_21_20_to_tile_21_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(692)
	);

	pe_tile pe_tile_21_20(
		.out_wire_3_0(vertical_tile_21_20_to_tile_20_20_0),
		.out_wire_3_1(vertical_tile_21_20_to_tile_20_20_1),
		.out_wire_3_2(vertical_tile_21_20_to_tile_20_20_2),
		.out_wire_3_3(vertical_tile_21_20_to_tile_20_20_3),
		.in_wire_3_0(vertical_tile_20_20_to_tile_21_20_0),
		.in_wire_3_1(vertical_tile_20_20_to_tile_21_20_1),
		.in_wire_3_2(vertical_tile_20_20_to_tile_21_20_2),
		.in_wire_3_3(vertical_tile_20_20_to_tile_21_20_3),
		.out_wire_1_0(vertical_tile_21_20_to_tile_22_20_0),
		.out_wire_1_1(vertical_tile_21_20_to_tile_22_20_1),
		.out_wire_1_2(vertical_tile_21_20_to_tile_22_20_2),
		.out_wire_1_3(vertical_tile_21_20_to_tile_22_20_3),
		.in_wire_1_0(vertical_tile_22_20_to_tile_21_20_0),
		.in_wire_1_1(vertical_tile_22_20_to_tile_21_20_1),
		.in_wire_1_2(vertical_tile_22_20_to_tile_21_20_2),
		.in_wire_1_3(vertical_tile_22_20_to_tile_21_20_3),
		.out_wire_2_0(horizontal_tile_21_20_to_tile_21_19_0),
		.out_wire_2_1(horizontal_tile_21_20_to_tile_21_19_1),
		.out_wire_2_2(horizontal_tile_21_20_to_tile_21_19_2),
		.out_wire_2_3(horizontal_tile_21_20_to_tile_21_19_3),
		.in_wire_2_0(horizontal_tile_21_19_to_tile_21_20_0),
		.in_wire_2_1(horizontal_tile_21_19_to_tile_21_20_1),
		.in_wire_2_2(horizontal_tile_21_19_to_tile_21_20_2),
		.in_wire_2_3(horizontal_tile_21_19_to_tile_21_20_3),
		.out_wire_0_0(horizontal_tile_21_20_to_tile_21_21_0),
		.out_wire_0_1(horizontal_tile_21_20_to_tile_21_21_1),
		.out_wire_0_2(horizontal_tile_21_20_to_tile_21_21_2),
		.out_wire_0_3(horizontal_tile_21_20_to_tile_21_21_3),
		.in_wire_0_0(horizontal_tile_21_21_to_tile_21_20_0),
		.in_wire_0_1(horizontal_tile_21_21_to_tile_21_20_1),
		.in_wire_0_2(horizontal_tile_21_21_to_tile_21_20_2),
		.in_wire_0_3(horizontal_tile_21_21_to_tile_21_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(693)
	);

	pe_tile pe_tile_21_21(
		.out_wire_3_0(vertical_tile_21_21_to_tile_20_21_0),
		.out_wire_3_1(vertical_tile_21_21_to_tile_20_21_1),
		.out_wire_3_2(vertical_tile_21_21_to_tile_20_21_2),
		.out_wire_3_3(vertical_tile_21_21_to_tile_20_21_3),
		.in_wire_3_0(vertical_tile_20_21_to_tile_21_21_0),
		.in_wire_3_1(vertical_tile_20_21_to_tile_21_21_1),
		.in_wire_3_2(vertical_tile_20_21_to_tile_21_21_2),
		.in_wire_3_3(vertical_tile_20_21_to_tile_21_21_3),
		.out_wire_1_0(vertical_tile_21_21_to_tile_22_21_0),
		.out_wire_1_1(vertical_tile_21_21_to_tile_22_21_1),
		.out_wire_1_2(vertical_tile_21_21_to_tile_22_21_2),
		.out_wire_1_3(vertical_tile_21_21_to_tile_22_21_3),
		.in_wire_1_0(vertical_tile_22_21_to_tile_21_21_0),
		.in_wire_1_1(vertical_tile_22_21_to_tile_21_21_1),
		.in_wire_1_2(vertical_tile_22_21_to_tile_21_21_2),
		.in_wire_1_3(vertical_tile_22_21_to_tile_21_21_3),
		.out_wire_2_0(horizontal_tile_21_21_to_tile_21_20_0),
		.out_wire_2_1(horizontal_tile_21_21_to_tile_21_20_1),
		.out_wire_2_2(horizontal_tile_21_21_to_tile_21_20_2),
		.out_wire_2_3(horizontal_tile_21_21_to_tile_21_20_3),
		.in_wire_2_0(horizontal_tile_21_20_to_tile_21_21_0),
		.in_wire_2_1(horizontal_tile_21_20_to_tile_21_21_1),
		.in_wire_2_2(horizontal_tile_21_20_to_tile_21_21_2),
		.in_wire_2_3(horizontal_tile_21_20_to_tile_21_21_3),
		.out_wire_0_0(horizontal_tile_21_21_to_tile_21_22_0),
		.out_wire_0_1(horizontal_tile_21_21_to_tile_21_22_1),
		.out_wire_0_2(horizontal_tile_21_21_to_tile_21_22_2),
		.out_wire_0_3(horizontal_tile_21_21_to_tile_21_22_3),
		.in_wire_0_0(horizontal_tile_21_22_to_tile_21_21_0),
		.in_wire_0_1(horizontal_tile_21_22_to_tile_21_21_1),
		.in_wire_0_2(horizontal_tile_21_22_to_tile_21_21_2),
		.in_wire_0_3(horizontal_tile_21_22_to_tile_21_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(694)
	);

	pe_tile pe_tile_21_22(
		.out_wire_3_0(vertical_tile_21_22_to_tile_20_22_0),
		.out_wire_3_1(vertical_tile_21_22_to_tile_20_22_1),
		.out_wire_3_2(vertical_tile_21_22_to_tile_20_22_2),
		.out_wire_3_3(vertical_tile_21_22_to_tile_20_22_3),
		.in_wire_3_0(vertical_tile_20_22_to_tile_21_22_0),
		.in_wire_3_1(vertical_tile_20_22_to_tile_21_22_1),
		.in_wire_3_2(vertical_tile_20_22_to_tile_21_22_2),
		.in_wire_3_3(vertical_tile_20_22_to_tile_21_22_3),
		.out_wire_1_0(vertical_tile_21_22_to_tile_22_22_0),
		.out_wire_1_1(vertical_tile_21_22_to_tile_22_22_1),
		.out_wire_1_2(vertical_tile_21_22_to_tile_22_22_2),
		.out_wire_1_3(vertical_tile_21_22_to_tile_22_22_3),
		.in_wire_1_0(vertical_tile_22_22_to_tile_21_22_0),
		.in_wire_1_1(vertical_tile_22_22_to_tile_21_22_1),
		.in_wire_1_2(vertical_tile_22_22_to_tile_21_22_2),
		.in_wire_1_3(vertical_tile_22_22_to_tile_21_22_3),
		.out_wire_2_0(horizontal_tile_21_22_to_tile_21_21_0),
		.out_wire_2_1(horizontal_tile_21_22_to_tile_21_21_1),
		.out_wire_2_2(horizontal_tile_21_22_to_tile_21_21_2),
		.out_wire_2_3(horizontal_tile_21_22_to_tile_21_21_3),
		.in_wire_2_0(horizontal_tile_21_21_to_tile_21_22_0),
		.in_wire_2_1(horizontal_tile_21_21_to_tile_21_22_1),
		.in_wire_2_2(horizontal_tile_21_21_to_tile_21_22_2),
		.in_wire_2_3(horizontal_tile_21_21_to_tile_21_22_3),
		.out_wire_0_0(horizontal_tile_21_22_to_tile_21_23_0),
		.out_wire_0_1(horizontal_tile_21_22_to_tile_21_23_1),
		.out_wire_0_2(horizontal_tile_21_22_to_tile_21_23_2),
		.out_wire_0_3(horizontal_tile_21_22_to_tile_21_23_3),
		.in_wire_0_0(horizontal_tile_21_23_to_tile_21_22_0),
		.in_wire_0_1(horizontal_tile_21_23_to_tile_21_22_1),
		.in_wire_0_2(horizontal_tile_21_23_to_tile_21_22_2),
		.in_wire_0_3(horizontal_tile_21_23_to_tile_21_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(695)
	);

	pe_tile pe_tile_21_23(
		.out_wire_3_0(vertical_tile_21_23_to_tile_20_23_0),
		.out_wire_3_1(vertical_tile_21_23_to_tile_20_23_1),
		.out_wire_3_2(vertical_tile_21_23_to_tile_20_23_2),
		.out_wire_3_3(vertical_tile_21_23_to_tile_20_23_3),
		.in_wire_3_0(vertical_tile_20_23_to_tile_21_23_0),
		.in_wire_3_1(vertical_tile_20_23_to_tile_21_23_1),
		.in_wire_3_2(vertical_tile_20_23_to_tile_21_23_2),
		.in_wire_3_3(vertical_tile_20_23_to_tile_21_23_3),
		.out_wire_1_0(vertical_tile_21_23_to_tile_22_23_0),
		.out_wire_1_1(vertical_tile_21_23_to_tile_22_23_1),
		.out_wire_1_2(vertical_tile_21_23_to_tile_22_23_2),
		.out_wire_1_3(vertical_tile_21_23_to_tile_22_23_3),
		.in_wire_1_0(vertical_tile_22_23_to_tile_21_23_0),
		.in_wire_1_1(vertical_tile_22_23_to_tile_21_23_1),
		.in_wire_1_2(vertical_tile_22_23_to_tile_21_23_2),
		.in_wire_1_3(vertical_tile_22_23_to_tile_21_23_3),
		.out_wire_2_0(horizontal_tile_21_23_to_tile_21_22_0),
		.out_wire_2_1(horizontal_tile_21_23_to_tile_21_22_1),
		.out_wire_2_2(horizontal_tile_21_23_to_tile_21_22_2),
		.out_wire_2_3(horizontal_tile_21_23_to_tile_21_22_3),
		.in_wire_2_0(horizontal_tile_21_22_to_tile_21_23_0),
		.in_wire_2_1(horizontal_tile_21_22_to_tile_21_23_1),
		.in_wire_2_2(horizontal_tile_21_22_to_tile_21_23_2),
		.in_wire_2_3(horizontal_tile_21_22_to_tile_21_23_3),
		.out_wire_0_0(horizontal_tile_21_23_to_tile_21_24_0),
		.out_wire_0_1(horizontal_tile_21_23_to_tile_21_24_1),
		.out_wire_0_2(horizontal_tile_21_23_to_tile_21_24_2),
		.out_wire_0_3(horizontal_tile_21_23_to_tile_21_24_3),
		.in_wire_0_0(horizontal_tile_21_24_to_tile_21_23_0),
		.in_wire_0_1(horizontal_tile_21_24_to_tile_21_23_1),
		.in_wire_0_2(horizontal_tile_21_24_to_tile_21_23_2),
		.in_wire_0_3(horizontal_tile_21_24_to_tile_21_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(696)
	);

	pe_tile pe_tile_21_24(
		.out_wire_3_0(vertical_tile_21_24_to_tile_20_24_0),
		.out_wire_3_1(vertical_tile_21_24_to_tile_20_24_1),
		.out_wire_3_2(vertical_tile_21_24_to_tile_20_24_2),
		.out_wire_3_3(vertical_tile_21_24_to_tile_20_24_3),
		.in_wire_3_0(vertical_tile_20_24_to_tile_21_24_0),
		.in_wire_3_1(vertical_tile_20_24_to_tile_21_24_1),
		.in_wire_3_2(vertical_tile_20_24_to_tile_21_24_2),
		.in_wire_3_3(vertical_tile_20_24_to_tile_21_24_3),
		.out_wire_1_0(vertical_tile_21_24_to_tile_22_24_0),
		.out_wire_1_1(vertical_tile_21_24_to_tile_22_24_1),
		.out_wire_1_2(vertical_tile_21_24_to_tile_22_24_2),
		.out_wire_1_3(vertical_tile_21_24_to_tile_22_24_3),
		.in_wire_1_0(vertical_tile_22_24_to_tile_21_24_0),
		.in_wire_1_1(vertical_tile_22_24_to_tile_21_24_1),
		.in_wire_1_2(vertical_tile_22_24_to_tile_21_24_2),
		.in_wire_1_3(vertical_tile_22_24_to_tile_21_24_3),
		.out_wire_2_0(horizontal_tile_21_24_to_tile_21_23_0),
		.out_wire_2_1(horizontal_tile_21_24_to_tile_21_23_1),
		.out_wire_2_2(horizontal_tile_21_24_to_tile_21_23_2),
		.out_wire_2_3(horizontal_tile_21_24_to_tile_21_23_3),
		.in_wire_2_0(horizontal_tile_21_23_to_tile_21_24_0),
		.in_wire_2_1(horizontal_tile_21_23_to_tile_21_24_1),
		.in_wire_2_2(horizontal_tile_21_23_to_tile_21_24_2),
		.in_wire_2_3(horizontal_tile_21_23_to_tile_21_24_3),
		.out_wire_0_0(horizontal_tile_21_24_to_tile_21_25_0),
		.out_wire_0_1(horizontal_tile_21_24_to_tile_21_25_1),
		.out_wire_0_2(horizontal_tile_21_24_to_tile_21_25_2),
		.out_wire_0_3(horizontal_tile_21_24_to_tile_21_25_3),
		.in_wire_0_0(horizontal_tile_21_25_to_tile_21_24_0),
		.in_wire_0_1(horizontal_tile_21_25_to_tile_21_24_1),
		.in_wire_0_2(horizontal_tile_21_25_to_tile_21_24_2),
		.in_wire_0_3(horizontal_tile_21_25_to_tile_21_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(697)
	);

	pe_tile pe_tile_21_25(
		.out_wire_3_0(vertical_tile_21_25_to_tile_20_25_0),
		.out_wire_3_1(vertical_tile_21_25_to_tile_20_25_1),
		.out_wire_3_2(vertical_tile_21_25_to_tile_20_25_2),
		.out_wire_3_3(vertical_tile_21_25_to_tile_20_25_3),
		.in_wire_3_0(vertical_tile_20_25_to_tile_21_25_0),
		.in_wire_3_1(vertical_tile_20_25_to_tile_21_25_1),
		.in_wire_3_2(vertical_tile_20_25_to_tile_21_25_2),
		.in_wire_3_3(vertical_tile_20_25_to_tile_21_25_3),
		.out_wire_1_0(vertical_tile_21_25_to_tile_22_25_0),
		.out_wire_1_1(vertical_tile_21_25_to_tile_22_25_1),
		.out_wire_1_2(vertical_tile_21_25_to_tile_22_25_2),
		.out_wire_1_3(vertical_tile_21_25_to_tile_22_25_3),
		.in_wire_1_0(vertical_tile_22_25_to_tile_21_25_0),
		.in_wire_1_1(vertical_tile_22_25_to_tile_21_25_1),
		.in_wire_1_2(vertical_tile_22_25_to_tile_21_25_2),
		.in_wire_1_3(vertical_tile_22_25_to_tile_21_25_3),
		.out_wire_2_0(horizontal_tile_21_25_to_tile_21_24_0),
		.out_wire_2_1(horizontal_tile_21_25_to_tile_21_24_1),
		.out_wire_2_2(horizontal_tile_21_25_to_tile_21_24_2),
		.out_wire_2_3(horizontal_tile_21_25_to_tile_21_24_3),
		.in_wire_2_0(horizontal_tile_21_24_to_tile_21_25_0),
		.in_wire_2_1(horizontal_tile_21_24_to_tile_21_25_1),
		.in_wire_2_2(horizontal_tile_21_24_to_tile_21_25_2),
		.in_wire_2_3(horizontal_tile_21_24_to_tile_21_25_3),
		.out_wire_0_0(horizontal_tile_21_25_to_tile_21_26_0),
		.out_wire_0_1(horizontal_tile_21_25_to_tile_21_26_1),
		.out_wire_0_2(horizontal_tile_21_25_to_tile_21_26_2),
		.out_wire_0_3(horizontal_tile_21_25_to_tile_21_26_3),
		.in_wire_0_0(horizontal_tile_21_26_to_tile_21_25_0),
		.in_wire_0_1(horizontal_tile_21_26_to_tile_21_25_1),
		.in_wire_0_2(horizontal_tile_21_26_to_tile_21_25_2),
		.in_wire_0_3(horizontal_tile_21_26_to_tile_21_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(698)
	);

	pe_tile pe_tile_21_26(
		.out_wire_3_0(vertical_tile_21_26_to_tile_20_26_0),
		.out_wire_3_1(vertical_tile_21_26_to_tile_20_26_1),
		.out_wire_3_2(vertical_tile_21_26_to_tile_20_26_2),
		.out_wire_3_3(vertical_tile_21_26_to_tile_20_26_3),
		.in_wire_3_0(vertical_tile_20_26_to_tile_21_26_0),
		.in_wire_3_1(vertical_tile_20_26_to_tile_21_26_1),
		.in_wire_3_2(vertical_tile_20_26_to_tile_21_26_2),
		.in_wire_3_3(vertical_tile_20_26_to_tile_21_26_3),
		.out_wire_1_0(vertical_tile_21_26_to_tile_22_26_0),
		.out_wire_1_1(vertical_tile_21_26_to_tile_22_26_1),
		.out_wire_1_2(vertical_tile_21_26_to_tile_22_26_2),
		.out_wire_1_3(vertical_tile_21_26_to_tile_22_26_3),
		.in_wire_1_0(vertical_tile_22_26_to_tile_21_26_0),
		.in_wire_1_1(vertical_tile_22_26_to_tile_21_26_1),
		.in_wire_1_2(vertical_tile_22_26_to_tile_21_26_2),
		.in_wire_1_3(vertical_tile_22_26_to_tile_21_26_3),
		.out_wire_2_0(horizontal_tile_21_26_to_tile_21_25_0),
		.out_wire_2_1(horizontal_tile_21_26_to_tile_21_25_1),
		.out_wire_2_2(horizontal_tile_21_26_to_tile_21_25_2),
		.out_wire_2_3(horizontal_tile_21_26_to_tile_21_25_3),
		.in_wire_2_0(horizontal_tile_21_25_to_tile_21_26_0),
		.in_wire_2_1(horizontal_tile_21_25_to_tile_21_26_1),
		.in_wire_2_2(horizontal_tile_21_25_to_tile_21_26_2),
		.in_wire_2_3(horizontal_tile_21_25_to_tile_21_26_3),
		.out_wire_0_0(horizontal_tile_21_26_to_tile_21_27_0),
		.out_wire_0_1(horizontal_tile_21_26_to_tile_21_27_1),
		.out_wire_0_2(horizontal_tile_21_26_to_tile_21_27_2),
		.out_wire_0_3(horizontal_tile_21_26_to_tile_21_27_3),
		.in_wire_0_0(horizontal_tile_21_27_to_tile_21_26_0),
		.in_wire_0_1(horizontal_tile_21_27_to_tile_21_26_1),
		.in_wire_0_2(horizontal_tile_21_27_to_tile_21_26_2),
		.in_wire_0_3(horizontal_tile_21_27_to_tile_21_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(699)
	);

	pe_tile pe_tile_21_27(
		.out_wire_3_0(vertical_tile_21_27_to_tile_20_27_0),
		.out_wire_3_1(vertical_tile_21_27_to_tile_20_27_1),
		.out_wire_3_2(vertical_tile_21_27_to_tile_20_27_2),
		.out_wire_3_3(vertical_tile_21_27_to_tile_20_27_3),
		.in_wire_3_0(vertical_tile_20_27_to_tile_21_27_0),
		.in_wire_3_1(vertical_tile_20_27_to_tile_21_27_1),
		.in_wire_3_2(vertical_tile_20_27_to_tile_21_27_2),
		.in_wire_3_3(vertical_tile_20_27_to_tile_21_27_3),
		.out_wire_1_0(vertical_tile_21_27_to_tile_22_27_0),
		.out_wire_1_1(vertical_tile_21_27_to_tile_22_27_1),
		.out_wire_1_2(vertical_tile_21_27_to_tile_22_27_2),
		.out_wire_1_3(vertical_tile_21_27_to_tile_22_27_3),
		.in_wire_1_0(vertical_tile_22_27_to_tile_21_27_0),
		.in_wire_1_1(vertical_tile_22_27_to_tile_21_27_1),
		.in_wire_1_2(vertical_tile_22_27_to_tile_21_27_2),
		.in_wire_1_3(vertical_tile_22_27_to_tile_21_27_3),
		.out_wire_2_0(horizontal_tile_21_27_to_tile_21_26_0),
		.out_wire_2_1(horizontal_tile_21_27_to_tile_21_26_1),
		.out_wire_2_2(horizontal_tile_21_27_to_tile_21_26_2),
		.out_wire_2_3(horizontal_tile_21_27_to_tile_21_26_3),
		.in_wire_2_0(horizontal_tile_21_26_to_tile_21_27_0),
		.in_wire_2_1(horizontal_tile_21_26_to_tile_21_27_1),
		.in_wire_2_2(horizontal_tile_21_26_to_tile_21_27_2),
		.in_wire_2_3(horizontal_tile_21_26_to_tile_21_27_3),
		.out_wire_0_0(horizontal_tile_21_27_to_tile_21_28_0),
		.out_wire_0_1(horizontal_tile_21_27_to_tile_21_28_1),
		.out_wire_0_2(horizontal_tile_21_27_to_tile_21_28_2),
		.out_wire_0_3(horizontal_tile_21_27_to_tile_21_28_3),
		.in_wire_0_0(horizontal_tile_21_28_to_tile_21_27_0),
		.in_wire_0_1(horizontal_tile_21_28_to_tile_21_27_1),
		.in_wire_0_2(horizontal_tile_21_28_to_tile_21_27_2),
		.in_wire_0_3(horizontal_tile_21_28_to_tile_21_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(700)
	);

	pe_tile pe_tile_21_28(
		.out_wire_3_0(vertical_tile_21_28_to_tile_20_28_0),
		.out_wire_3_1(vertical_tile_21_28_to_tile_20_28_1),
		.out_wire_3_2(vertical_tile_21_28_to_tile_20_28_2),
		.out_wire_3_3(vertical_tile_21_28_to_tile_20_28_3),
		.in_wire_3_0(vertical_tile_20_28_to_tile_21_28_0),
		.in_wire_3_1(vertical_tile_20_28_to_tile_21_28_1),
		.in_wire_3_2(vertical_tile_20_28_to_tile_21_28_2),
		.in_wire_3_3(vertical_tile_20_28_to_tile_21_28_3),
		.out_wire_1_0(vertical_tile_21_28_to_tile_22_28_0),
		.out_wire_1_1(vertical_tile_21_28_to_tile_22_28_1),
		.out_wire_1_2(vertical_tile_21_28_to_tile_22_28_2),
		.out_wire_1_3(vertical_tile_21_28_to_tile_22_28_3),
		.in_wire_1_0(vertical_tile_22_28_to_tile_21_28_0),
		.in_wire_1_1(vertical_tile_22_28_to_tile_21_28_1),
		.in_wire_1_2(vertical_tile_22_28_to_tile_21_28_2),
		.in_wire_1_3(vertical_tile_22_28_to_tile_21_28_3),
		.out_wire_2_0(horizontal_tile_21_28_to_tile_21_27_0),
		.out_wire_2_1(horizontal_tile_21_28_to_tile_21_27_1),
		.out_wire_2_2(horizontal_tile_21_28_to_tile_21_27_2),
		.out_wire_2_3(horizontal_tile_21_28_to_tile_21_27_3),
		.in_wire_2_0(horizontal_tile_21_27_to_tile_21_28_0),
		.in_wire_2_1(horizontal_tile_21_27_to_tile_21_28_1),
		.in_wire_2_2(horizontal_tile_21_27_to_tile_21_28_2),
		.in_wire_2_3(horizontal_tile_21_27_to_tile_21_28_3),
		.out_wire_0_0(horizontal_tile_21_28_to_tile_21_29_0),
		.out_wire_0_1(horizontal_tile_21_28_to_tile_21_29_1),
		.out_wire_0_2(horizontal_tile_21_28_to_tile_21_29_2),
		.out_wire_0_3(horizontal_tile_21_28_to_tile_21_29_3),
		.in_wire_0_0(horizontal_tile_21_29_to_tile_21_28_0),
		.in_wire_0_1(horizontal_tile_21_29_to_tile_21_28_1),
		.in_wire_0_2(horizontal_tile_21_29_to_tile_21_28_2),
		.in_wire_0_3(horizontal_tile_21_29_to_tile_21_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(701)
	);

	pe_tile pe_tile_21_29(
		.out_wire_3_0(vertical_tile_21_29_to_tile_20_29_0),
		.out_wire_3_1(vertical_tile_21_29_to_tile_20_29_1),
		.out_wire_3_2(vertical_tile_21_29_to_tile_20_29_2),
		.out_wire_3_3(vertical_tile_21_29_to_tile_20_29_3),
		.in_wire_3_0(vertical_tile_20_29_to_tile_21_29_0),
		.in_wire_3_1(vertical_tile_20_29_to_tile_21_29_1),
		.in_wire_3_2(vertical_tile_20_29_to_tile_21_29_2),
		.in_wire_3_3(vertical_tile_20_29_to_tile_21_29_3),
		.out_wire_1_0(vertical_tile_21_29_to_tile_22_29_0),
		.out_wire_1_1(vertical_tile_21_29_to_tile_22_29_1),
		.out_wire_1_2(vertical_tile_21_29_to_tile_22_29_2),
		.out_wire_1_3(vertical_tile_21_29_to_tile_22_29_3),
		.in_wire_1_0(vertical_tile_22_29_to_tile_21_29_0),
		.in_wire_1_1(vertical_tile_22_29_to_tile_21_29_1),
		.in_wire_1_2(vertical_tile_22_29_to_tile_21_29_2),
		.in_wire_1_3(vertical_tile_22_29_to_tile_21_29_3),
		.out_wire_2_0(horizontal_tile_21_29_to_tile_21_28_0),
		.out_wire_2_1(horizontal_tile_21_29_to_tile_21_28_1),
		.out_wire_2_2(horizontal_tile_21_29_to_tile_21_28_2),
		.out_wire_2_3(horizontal_tile_21_29_to_tile_21_28_3),
		.in_wire_2_0(horizontal_tile_21_28_to_tile_21_29_0),
		.in_wire_2_1(horizontal_tile_21_28_to_tile_21_29_1),
		.in_wire_2_2(horizontal_tile_21_28_to_tile_21_29_2),
		.in_wire_2_3(horizontal_tile_21_28_to_tile_21_29_3),
		.out_wire_0_0(horizontal_tile_21_29_to_tile_21_30_0),
		.out_wire_0_1(horizontal_tile_21_29_to_tile_21_30_1),
		.out_wire_0_2(horizontal_tile_21_29_to_tile_21_30_2),
		.out_wire_0_3(horizontal_tile_21_29_to_tile_21_30_3),
		.in_wire_0_0(horizontal_tile_21_30_to_tile_21_29_0),
		.in_wire_0_1(horizontal_tile_21_30_to_tile_21_29_1),
		.in_wire_0_2(horizontal_tile_21_30_to_tile_21_29_2),
		.in_wire_0_3(horizontal_tile_21_30_to_tile_21_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(702)
	);

	pe_tile pe_tile_21_30(
		.out_wire_3_0(vertical_tile_21_30_to_tile_20_30_0),
		.out_wire_3_1(vertical_tile_21_30_to_tile_20_30_1),
		.out_wire_3_2(vertical_tile_21_30_to_tile_20_30_2),
		.out_wire_3_3(vertical_tile_21_30_to_tile_20_30_3),
		.in_wire_3_0(vertical_tile_20_30_to_tile_21_30_0),
		.in_wire_3_1(vertical_tile_20_30_to_tile_21_30_1),
		.in_wire_3_2(vertical_tile_20_30_to_tile_21_30_2),
		.in_wire_3_3(vertical_tile_20_30_to_tile_21_30_3),
		.out_wire_1_0(vertical_tile_21_30_to_tile_22_30_0),
		.out_wire_1_1(vertical_tile_21_30_to_tile_22_30_1),
		.out_wire_1_2(vertical_tile_21_30_to_tile_22_30_2),
		.out_wire_1_3(vertical_tile_21_30_to_tile_22_30_3),
		.in_wire_1_0(vertical_tile_22_30_to_tile_21_30_0),
		.in_wire_1_1(vertical_tile_22_30_to_tile_21_30_1),
		.in_wire_1_2(vertical_tile_22_30_to_tile_21_30_2),
		.in_wire_1_3(vertical_tile_22_30_to_tile_21_30_3),
		.out_wire_2_0(horizontal_tile_21_30_to_tile_21_29_0),
		.out_wire_2_1(horizontal_tile_21_30_to_tile_21_29_1),
		.out_wire_2_2(horizontal_tile_21_30_to_tile_21_29_2),
		.out_wire_2_3(horizontal_tile_21_30_to_tile_21_29_3),
		.in_wire_2_0(horizontal_tile_21_29_to_tile_21_30_0),
		.in_wire_2_1(horizontal_tile_21_29_to_tile_21_30_1),
		.in_wire_2_2(horizontal_tile_21_29_to_tile_21_30_2),
		.in_wire_2_3(horizontal_tile_21_29_to_tile_21_30_3),
		.out_wire_0_0(horizontal_tile_21_30_to_tile_21_31_0),
		.out_wire_0_1(horizontal_tile_21_30_to_tile_21_31_1),
		.out_wire_0_2(horizontal_tile_21_30_to_tile_21_31_2),
		.out_wire_0_3(horizontal_tile_21_30_to_tile_21_31_3),
		.in_wire_0_0(horizontal_tile_21_31_to_tile_21_30_0),
		.in_wire_0_1(horizontal_tile_21_31_to_tile_21_30_1),
		.in_wire_0_2(horizontal_tile_21_31_to_tile_21_30_2),
		.in_wire_0_3(horizontal_tile_21_31_to_tile_21_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(703)
	);

	pe_tile_right pe_tile_21_31(
		.out_wire_3_0(vertical_tile_21_31_to_tile_20_31_0),
		.out_wire_3_1(vertical_tile_21_31_to_tile_20_31_1),
		.out_wire_3_2(vertical_tile_21_31_to_tile_20_31_2),
		.out_wire_3_3(vertical_tile_21_31_to_tile_20_31_3),
		.in_wire_3_0(vertical_tile_20_31_to_tile_21_31_0),
		.in_wire_3_1(vertical_tile_20_31_to_tile_21_31_1),
		.in_wire_3_2(vertical_tile_20_31_to_tile_21_31_2),
		.in_wire_3_3(vertical_tile_20_31_to_tile_21_31_3),
		.out_wire_1_0(vertical_tile_21_31_to_tile_22_31_0),
		.out_wire_1_1(vertical_tile_21_31_to_tile_22_31_1),
		.out_wire_1_2(vertical_tile_21_31_to_tile_22_31_2),
		.out_wire_1_3(vertical_tile_21_31_to_tile_22_31_3),
		.in_wire_1_0(vertical_tile_22_31_to_tile_21_31_0),
		.in_wire_1_1(vertical_tile_22_31_to_tile_21_31_1),
		.in_wire_1_2(vertical_tile_22_31_to_tile_21_31_2),
		.in_wire_1_3(vertical_tile_22_31_to_tile_21_31_3),
		.out_wire_2_0(horizontal_tile_21_31_to_tile_21_30_0),
		.out_wire_2_1(horizontal_tile_21_31_to_tile_21_30_1),
		.out_wire_2_2(horizontal_tile_21_31_to_tile_21_30_2),
		.out_wire_2_3(horizontal_tile_21_31_to_tile_21_30_3),
		.in_wire_2_0(horizontal_tile_21_30_to_tile_21_31_0),
		.in_wire_2_1(horizontal_tile_21_30_to_tile_21_31_1),
		.in_wire_2_2(horizontal_tile_21_30_to_tile_21_31_2),
		.in_wire_2_3(horizontal_tile_21_30_to_tile_21_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(704)
	);

	pe_tile_left pe_tile_22_0(
		.out_wire_3_0(vertical_tile_22_0_to_tile_21_0_0),
		.out_wire_3_1(vertical_tile_22_0_to_tile_21_0_1),
		.out_wire_3_2(vertical_tile_22_0_to_tile_21_0_2),
		.out_wire_3_3(vertical_tile_22_0_to_tile_21_0_3),
		.in_wire_3_0(vertical_tile_21_0_to_tile_22_0_0),
		.in_wire_3_1(vertical_tile_21_0_to_tile_22_0_1),
		.in_wire_3_2(vertical_tile_21_0_to_tile_22_0_2),
		.in_wire_3_3(vertical_tile_21_0_to_tile_22_0_3),
		.out_wire_1_0(vertical_tile_22_0_to_tile_23_0_0),
		.out_wire_1_1(vertical_tile_22_0_to_tile_23_0_1),
		.out_wire_1_2(vertical_tile_22_0_to_tile_23_0_2),
		.out_wire_1_3(vertical_tile_22_0_to_tile_23_0_3),
		.in_wire_1_0(vertical_tile_23_0_to_tile_22_0_0),
		.in_wire_1_1(vertical_tile_23_0_to_tile_22_0_1),
		.in_wire_1_2(vertical_tile_23_0_to_tile_22_0_2),
		.in_wire_1_3(vertical_tile_23_0_to_tile_22_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_22_0_to_tile_22_1_0),
		.out_wire_0_1(horizontal_tile_22_0_to_tile_22_1_1),
		.out_wire_0_2(horizontal_tile_22_0_to_tile_22_1_2),
		.out_wire_0_3(horizontal_tile_22_0_to_tile_22_1_3),
		.in_wire_0_0(horizontal_tile_22_1_to_tile_22_0_0),
		.in_wire_0_1(horizontal_tile_22_1_to_tile_22_0_1),
		.in_wire_0_2(horizontal_tile_22_1_to_tile_22_0_2),
		.in_wire_0_3(horizontal_tile_22_1_to_tile_22_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(705)
	);

	pe_tile pe_tile_22_1(
		.out_wire_3_0(vertical_tile_22_1_to_tile_21_1_0),
		.out_wire_3_1(vertical_tile_22_1_to_tile_21_1_1),
		.out_wire_3_2(vertical_tile_22_1_to_tile_21_1_2),
		.out_wire_3_3(vertical_tile_22_1_to_tile_21_1_3),
		.in_wire_3_0(vertical_tile_21_1_to_tile_22_1_0),
		.in_wire_3_1(vertical_tile_21_1_to_tile_22_1_1),
		.in_wire_3_2(vertical_tile_21_1_to_tile_22_1_2),
		.in_wire_3_3(vertical_tile_21_1_to_tile_22_1_3),
		.out_wire_1_0(vertical_tile_22_1_to_tile_23_1_0),
		.out_wire_1_1(vertical_tile_22_1_to_tile_23_1_1),
		.out_wire_1_2(vertical_tile_22_1_to_tile_23_1_2),
		.out_wire_1_3(vertical_tile_22_1_to_tile_23_1_3),
		.in_wire_1_0(vertical_tile_23_1_to_tile_22_1_0),
		.in_wire_1_1(vertical_tile_23_1_to_tile_22_1_1),
		.in_wire_1_2(vertical_tile_23_1_to_tile_22_1_2),
		.in_wire_1_3(vertical_tile_23_1_to_tile_22_1_3),
		.out_wire_2_0(horizontal_tile_22_1_to_tile_22_0_0),
		.out_wire_2_1(horizontal_tile_22_1_to_tile_22_0_1),
		.out_wire_2_2(horizontal_tile_22_1_to_tile_22_0_2),
		.out_wire_2_3(horizontal_tile_22_1_to_tile_22_0_3),
		.in_wire_2_0(horizontal_tile_22_0_to_tile_22_1_0),
		.in_wire_2_1(horizontal_tile_22_0_to_tile_22_1_1),
		.in_wire_2_2(horizontal_tile_22_0_to_tile_22_1_2),
		.in_wire_2_3(horizontal_tile_22_0_to_tile_22_1_3),
		.out_wire_0_0(horizontal_tile_22_1_to_tile_22_2_0),
		.out_wire_0_1(horizontal_tile_22_1_to_tile_22_2_1),
		.out_wire_0_2(horizontal_tile_22_1_to_tile_22_2_2),
		.out_wire_0_3(horizontal_tile_22_1_to_tile_22_2_3),
		.in_wire_0_0(horizontal_tile_22_2_to_tile_22_1_0),
		.in_wire_0_1(horizontal_tile_22_2_to_tile_22_1_1),
		.in_wire_0_2(horizontal_tile_22_2_to_tile_22_1_2),
		.in_wire_0_3(horizontal_tile_22_2_to_tile_22_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(706)
	);

	pe_tile pe_tile_22_2(
		.out_wire_3_0(vertical_tile_22_2_to_tile_21_2_0),
		.out_wire_3_1(vertical_tile_22_2_to_tile_21_2_1),
		.out_wire_3_2(vertical_tile_22_2_to_tile_21_2_2),
		.out_wire_3_3(vertical_tile_22_2_to_tile_21_2_3),
		.in_wire_3_0(vertical_tile_21_2_to_tile_22_2_0),
		.in_wire_3_1(vertical_tile_21_2_to_tile_22_2_1),
		.in_wire_3_2(vertical_tile_21_2_to_tile_22_2_2),
		.in_wire_3_3(vertical_tile_21_2_to_tile_22_2_3),
		.out_wire_1_0(vertical_tile_22_2_to_tile_23_2_0),
		.out_wire_1_1(vertical_tile_22_2_to_tile_23_2_1),
		.out_wire_1_2(vertical_tile_22_2_to_tile_23_2_2),
		.out_wire_1_3(vertical_tile_22_2_to_tile_23_2_3),
		.in_wire_1_0(vertical_tile_23_2_to_tile_22_2_0),
		.in_wire_1_1(vertical_tile_23_2_to_tile_22_2_1),
		.in_wire_1_2(vertical_tile_23_2_to_tile_22_2_2),
		.in_wire_1_3(vertical_tile_23_2_to_tile_22_2_3),
		.out_wire_2_0(horizontal_tile_22_2_to_tile_22_1_0),
		.out_wire_2_1(horizontal_tile_22_2_to_tile_22_1_1),
		.out_wire_2_2(horizontal_tile_22_2_to_tile_22_1_2),
		.out_wire_2_3(horizontal_tile_22_2_to_tile_22_1_3),
		.in_wire_2_0(horizontal_tile_22_1_to_tile_22_2_0),
		.in_wire_2_1(horizontal_tile_22_1_to_tile_22_2_1),
		.in_wire_2_2(horizontal_tile_22_1_to_tile_22_2_2),
		.in_wire_2_3(horizontal_tile_22_1_to_tile_22_2_3),
		.out_wire_0_0(horizontal_tile_22_2_to_tile_22_3_0),
		.out_wire_0_1(horizontal_tile_22_2_to_tile_22_3_1),
		.out_wire_0_2(horizontal_tile_22_2_to_tile_22_3_2),
		.out_wire_0_3(horizontal_tile_22_2_to_tile_22_3_3),
		.in_wire_0_0(horizontal_tile_22_3_to_tile_22_2_0),
		.in_wire_0_1(horizontal_tile_22_3_to_tile_22_2_1),
		.in_wire_0_2(horizontal_tile_22_3_to_tile_22_2_2),
		.in_wire_0_3(horizontal_tile_22_3_to_tile_22_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(707)
	);

	pe_tile pe_tile_22_3(
		.out_wire_3_0(vertical_tile_22_3_to_tile_21_3_0),
		.out_wire_3_1(vertical_tile_22_3_to_tile_21_3_1),
		.out_wire_3_2(vertical_tile_22_3_to_tile_21_3_2),
		.out_wire_3_3(vertical_tile_22_3_to_tile_21_3_3),
		.in_wire_3_0(vertical_tile_21_3_to_tile_22_3_0),
		.in_wire_3_1(vertical_tile_21_3_to_tile_22_3_1),
		.in_wire_3_2(vertical_tile_21_3_to_tile_22_3_2),
		.in_wire_3_3(vertical_tile_21_3_to_tile_22_3_3),
		.out_wire_1_0(vertical_tile_22_3_to_tile_23_3_0),
		.out_wire_1_1(vertical_tile_22_3_to_tile_23_3_1),
		.out_wire_1_2(vertical_tile_22_3_to_tile_23_3_2),
		.out_wire_1_3(vertical_tile_22_3_to_tile_23_3_3),
		.in_wire_1_0(vertical_tile_23_3_to_tile_22_3_0),
		.in_wire_1_1(vertical_tile_23_3_to_tile_22_3_1),
		.in_wire_1_2(vertical_tile_23_3_to_tile_22_3_2),
		.in_wire_1_3(vertical_tile_23_3_to_tile_22_3_3),
		.out_wire_2_0(horizontal_tile_22_3_to_tile_22_2_0),
		.out_wire_2_1(horizontal_tile_22_3_to_tile_22_2_1),
		.out_wire_2_2(horizontal_tile_22_3_to_tile_22_2_2),
		.out_wire_2_3(horizontal_tile_22_3_to_tile_22_2_3),
		.in_wire_2_0(horizontal_tile_22_2_to_tile_22_3_0),
		.in_wire_2_1(horizontal_tile_22_2_to_tile_22_3_1),
		.in_wire_2_2(horizontal_tile_22_2_to_tile_22_3_2),
		.in_wire_2_3(horizontal_tile_22_2_to_tile_22_3_3),
		.out_wire_0_0(horizontal_tile_22_3_to_tile_22_4_0),
		.out_wire_0_1(horizontal_tile_22_3_to_tile_22_4_1),
		.out_wire_0_2(horizontal_tile_22_3_to_tile_22_4_2),
		.out_wire_0_3(horizontal_tile_22_3_to_tile_22_4_3),
		.in_wire_0_0(horizontal_tile_22_4_to_tile_22_3_0),
		.in_wire_0_1(horizontal_tile_22_4_to_tile_22_3_1),
		.in_wire_0_2(horizontal_tile_22_4_to_tile_22_3_2),
		.in_wire_0_3(horizontal_tile_22_4_to_tile_22_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(708)
	);

	pe_tile pe_tile_22_4(
		.out_wire_3_0(vertical_tile_22_4_to_tile_21_4_0),
		.out_wire_3_1(vertical_tile_22_4_to_tile_21_4_1),
		.out_wire_3_2(vertical_tile_22_4_to_tile_21_4_2),
		.out_wire_3_3(vertical_tile_22_4_to_tile_21_4_3),
		.in_wire_3_0(vertical_tile_21_4_to_tile_22_4_0),
		.in_wire_3_1(vertical_tile_21_4_to_tile_22_4_1),
		.in_wire_3_2(vertical_tile_21_4_to_tile_22_4_2),
		.in_wire_3_3(vertical_tile_21_4_to_tile_22_4_3),
		.out_wire_1_0(vertical_tile_22_4_to_tile_23_4_0),
		.out_wire_1_1(vertical_tile_22_4_to_tile_23_4_1),
		.out_wire_1_2(vertical_tile_22_4_to_tile_23_4_2),
		.out_wire_1_3(vertical_tile_22_4_to_tile_23_4_3),
		.in_wire_1_0(vertical_tile_23_4_to_tile_22_4_0),
		.in_wire_1_1(vertical_tile_23_4_to_tile_22_4_1),
		.in_wire_1_2(vertical_tile_23_4_to_tile_22_4_2),
		.in_wire_1_3(vertical_tile_23_4_to_tile_22_4_3),
		.out_wire_2_0(horizontal_tile_22_4_to_tile_22_3_0),
		.out_wire_2_1(horizontal_tile_22_4_to_tile_22_3_1),
		.out_wire_2_2(horizontal_tile_22_4_to_tile_22_3_2),
		.out_wire_2_3(horizontal_tile_22_4_to_tile_22_3_3),
		.in_wire_2_0(horizontal_tile_22_3_to_tile_22_4_0),
		.in_wire_2_1(horizontal_tile_22_3_to_tile_22_4_1),
		.in_wire_2_2(horizontal_tile_22_3_to_tile_22_4_2),
		.in_wire_2_3(horizontal_tile_22_3_to_tile_22_4_3),
		.out_wire_0_0(horizontal_tile_22_4_to_tile_22_5_0),
		.out_wire_0_1(horizontal_tile_22_4_to_tile_22_5_1),
		.out_wire_0_2(horizontal_tile_22_4_to_tile_22_5_2),
		.out_wire_0_3(horizontal_tile_22_4_to_tile_22_5_3),
		.in_wire_0_0(horizontal_tile_22_5_to_tile_22_4_0),
		.in_wire_0_1(horizontal_tile_22_5_to_tile_22_4_1),
		.in_wire_0_2(horizontal_tile_22_5_to_tile_22_4_2),
		.in_wire_0_3(horizontal_tile_22_5_to_tile_22_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(709)
	);

	pe_tile pe_tile_22_5(
		.out_wire_3_0(vertical_tile_22_5_to_tile_21_5_0),
		.out_wire_3_1(vertical_tile_22_5_to_tile_21_5_1),
		.out_wire_3_2(vertical_tile_22_5_to_tile_21_5_2),
		.out_wire_3_3(vertical_tile_22_5_to_tile_21_5_3),
		.in_wire_3_0(vertical_tile_21_5_to_tile_22_5_0),
		.in_wire_3_1(vertical_tile_21_5_to_tile_22_5_1),
		.in_wire_3_2(vertical_tile_21_5_to_tile_22_5_2),
		.in_wire_3_3(vertical_tile_21_5_to_tile_22_5_3),
		.out_wire_1_0(vertical_tile_22_5_to_tile_23_5_0),
		.out_wire_1_1(vertical_tile_22_5_to_tile_23_5_1),
		.out_wire_1_2(vertical_tile_22_5_to_tile_23_5_2),
		.out_wire_1_3(vertical_tile_22_5_to_tile_23_5_3),
		.in_wire_1_0(vertical_tile_23_5_to_tile_22_5_0),
		.in_wire_1_1(vertical_tile_23_5_to_tile_22_5_1),
		.in_wire_1_2(vertical_tile_23_5_to_tile_22_5_2),
		.in_wire_1_3(vertical_tile_23_5_to_tile_22_5_3),
		.out_wire_2_0(horizontal_tile_22_5_to_tile_22_4_0),
		.out_wire_2_1(horizontal_tile_22_5_to_tile_22_4_1),
		.out_wire_2_2(horizontal_tile_22_5_to_tile_22_4_2),
		.out_wire_2_3(horizontal_tile_22_5_to_tile_22_4_3),
		.in_wire_2_0(horizontal_tile_22_4_to_tile_22_5_0),
		.in_wire_2_1(horizontal_tile_22_4_to_tile_22_5_1),
		.in_wire_2_2(horizontal_tile_22_4_to_tile_22_5_2),
		.in_wire_2_3(horizontal_tile_22_4_to_tile_22_5_3),
		.out_wire_0_0(horizontal_tile_22_5_to_tile_22_6_0),
		.out_wire_0_1(horizontal_tile_22_5_to_tile_22_6_1),
		.out_wire_0_2(horizontal_tile_22_5_to_tile_22_6_2),
		.out_wire_0_3(horizontal_tile_22_5_to_tile_22_6_3),
		.in_wire_0_0(horizontal_tile_22_6_to_tile_22_5_0),
		.in_wire_0_1(horizontal_tile_22_6_to_tile_22_5_1),
		.in_wire_0_2(horizontal_tile_22_6_to_tile_22_5_2),
		.in_wire_0_3(horizontal_tile_22_6_to_tile_22_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(710)
	);

	pe_tile pe_tile_22_6(
		.out_wire_3_0(vertical_tile_22_6_to_tile_21_6_0),
		.out_wire_3_1(vertical_tile_22_6_to_tile_21_6_1),
		.out_wire_3_2(vertical_tile_22_6_to_tile_21_6_2),
		.out_wire_3_3(vertical_tile_22_6_to_tile_21_6_3),
		.in_wire_3_0(vertical_tile_21_6_to_tile_22_6_0),
		.in_wire_3_1(vertical_tile_21_6_to_tile_22_6_1),
		.in_wire_3_2(vertical_tile_21_6_to_tile_22_6_2),
		.in_wire_3_3(vertical_tile_21_6_to_tile_22_6_3),
		.out_wire_1_0(vertical_tile_22_6_to_tile_23_6_0),
		.out_wire_1_1(vertical_tile_22_6_to_tile_23_6_1),
		.out_wire_1_2(vertical_tile_22_6_to_tile_23_6_2),
		.out_wire_1_3(vertical_tile_22_6_to_tile_23_6_3),
		.in_wire_1_0(vertical_tile_23_6_to_tile_22_6_0),
		.in_wire_1_1(vertical_tile_23_6_to_tile_22_6_1),
		.in_wire_1_2(vertical_tile_23_6_to_tile_22_6_2),
		.in_wire_1_3(vertical_tile_23_6_to_tile_22_6_3),
		.out_wire_2_0(horizontal_tile_22_6_to_tile_22_5_0),
		.out_wire_2_1(horizontal_tile_22_6_to_tile_22_5_1),
		.out_wire_2_2(horizontal_tile_22_6_to_tile_22_5_2),
		.out_wire_2_3(horizontal_tile_22_6_to_tile_22_5_3),
		.in_wire_2_0(horizontal_tile_22_5_to_tile_22_6_0),
		.in_wire_2_1(horizontal_tile_22_5_to_tile_22_6_1),
		.in_wire_2_2(horizontal_tile_22_5_to_tile_22_6_2),
		.in_wire_2_3(horizontal_tile_22_5_to_tile_22_6_3),
		.out_wire_0_0(horizontal_tile_22_6_to_tile_22_7_0),
		.out_wire_0_1(horizontal_tile_22_6_to_tile_22_7_1),
		.out_wire_0_2(horizontal_tile_22_6_to_tile_22_7_2),
		.out_wire_0_3(horizontal_tile_22_6_to_tile_22_7_3),
		.in_wire_0_0(horizontal_tile_22_7_to_tile_22_6_0),
		.in_wire_0_1(horizontal_tile_22_7_to_tile_22_6_1),
		.in_wire_0_2(horizontal_tile_22_7_to_tile_22_6_2),
		.in_wire_0_3(horizontal_tile_22_7_to_tile_22_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(711)
	);

	pe_tile pe_tile_22_7(
		.out_wire_3_0(vertical_tile_22_7_to_tile_21_7_0),
		.out_wire_3_1(vertical_tile_22_7_to_tile_21_7_1),
		.out_wire_3_2(vertical_tile_22_7_to_tile_21_7_2),
		.out_wire_3_3(vertical_tile_22_7_to_tile_21_7_3),
		.in_wire_3_0(vertical_tile_21_7_to_tile_22_7_0),
		.in_wire_3_1(vertical_tile_21_7_to_tile_22_7_1),
		.in_wire_3_2(vertical_tile_21_7_to_tile_22_7_2),
		.in_wire_3_3(vertical_tile_21_7_to_tile_22_7_3),
		.out_wire_1_0(vertical_tile_22_7_to_tile_23_7_0),
		.out_wire_1_1(vertical_tile_22_7_to_tile_23_7_1),
		.out_wire_1_2(vertical_tile_22_7_to_tile_23_7_2),
		.out_wire_1_3(vertical_tile_22_7_to_tile_23_7_3),
		.in_wire_1_0(vertical_tile_23_7_to_tile_22_7_0),
		.in_wire_1_1(vertical_tile_23_7_to_tile_22_7_1),
		.in_wire_1_2(vertical_tile_23_7_to_tile_22_7_2),
		.in_wire_1_3(vertical_tile_23_7_to_tile_22_7_3),
		.out_wire_2_0(horizontal_tile_22_7_to_tile_22_6_0),
		.out_wire_2_1(horizontal_tile_22_7_to_tile_22_6_1),
		.out_wire_2_2(horizontal_tile_22_7_to_tile_22_6_2),
		.out_wire_2_3(horizontal_tile_22_7_to_tile_22_6_3),
		.in_wire_2_0(horizontal_tile_22_6_to_tile_22_7_0),
		.in_wire_2_1(horizontal_tile_22_6_to_tile_22_7_1),
		.in_wire_2_2(horizontal_tile_22_6_to_tile_22_7_2),
		.in_wire_2_3(horizontal_tile_22_6_to_tile_22_7_3),
		.out_wire_0_0(horizontal_tile_22_7_to_tile_22_8_0),
		.out_wire_0_1(horizontal_tile_22_7_to_tile_22_8_1),
		.out_wire_0_2(horizontal_tile_22_7_to_tile_22_8_2),
		.out_wire_0_3(horizontal_tile_22_7_to_tile_22_8_3),
		.in_wire_0_0(horizontal_tile_22_8_to_tile_22_7_0),
		.in_wire_0_1(horizontal_tile_22_8_to_tile_22_7_1),
		.in_wire_0_2(horizontal_tile_22_8_to_tile_22_7_2),
		.in_wire_0_3(horizontal_tile_22_8_to_tile_22_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(712)
	);

	pe_tile pe_tile_22_8(
		.out_wire_3_0(vertical_tile_22_8_to_tile_21_8_0),
		.out_wire_3_1(vertical_tile_22_8_to_tile_21_8_1),
		.out_wire_3_2(vertical_tile_22_8_to_tile_21_8_2),
		.out_wire_3_3(vertical_tile_22_8_to_tile_21_8_3),
		.in_wire_3_0(vertical_tile_21_8_to_tile_22_8_0),
		.in_wire_3_1(vertical_tile_21_8_to_tile_22_8_1),
		.in_wire_3_2(vertical_tile_21_8_to_tile_22_8_2),
		.in_wire_3_3(vertical_tile_21_8_to_tile_22_8_3),
		.out_wire_1_0(vertical_tile_22_8_to_tile_23_8_0),
		.out_wire_1_1(vertical_tile_22_8_to_tile_23_8_1),
		.out_wire_1_2(vertical_tile_22_8_to_tile_23_8_2),
		.out_wire_1_3(vertical_tile_22_8_to_tile_23_8_3),
		.in_wire_1_0(vertical_tile_23_8_to_tile_22_8_0),
		.in_wire_1_1(vertical_tile_23_8_to_tile_22_8_1),
		.in_wire_1_2(vertical_tile_23_8_to_tile_22_8_2),
		.in_wire_1_3(vertical_tile_23_8_to_tile_22_8_3),
		.out_wire_2_0(horizontal_tile_22_8_to_tile_22_7_0),
		.out_wire_2_1(horizontal_tile_22_8_to_tile_22_7_1),
		.out_wire_2_2(horizontal_tile_22_8_to_tile_22_7_2),
		.out_wire_2_3(horizontal_tile_22_8_to_tile_22_7_3),
		.in_wire_2_0(horizontal_tile_22_7_to_tile_22_8_0),
		.in_wire_2_1(horizontal_tile_22_7_to_tile_22_8_1),
		.in_wire_2_2(horizontal_tile_22_7_to_tile_22_8_2),
		.in_wire_2_3(horizontal_tile_22_7_to_tile_22_8_3),
		.out_wire_0_0(horizontal_tile_22_8_to_tile_22_9_0),
		.out_wire_0_1(horizontal_tile_22_8_to_tile_22_9_1),
		.out_wire_0_2(horizontal_tile_22_8_to_tile_22_9_2),
		.out_wire_0_3(horizontal_tile_22_8_to_tile_22_9_3),
		.in_wire_0_0(horizontal_tile_22_9_to_tile_22_8_0),
		.in_wire_0_1(horizontal_tile_22_9_to_tile_22_8_1),
		.in_wire_0_2(horizontal_tile_22_9_to_tile_22_8_2),
		.in_wire_0_3(horizontal_tile_22_9_to_tile_22_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(713)
	);

	pe_tile pe_tile_22_9(
		.out_wire_3_0(vertical_tile_22_9_to_tile_21_9_0),
		.out_wire_3_1(vertical_tile_22_9_to_tile_21_9_1),
		.out_wire_3_2(vertical_tile_22_9_to_tile_21_9_2),
		.out_wire_3_3(vertical_tile_22_9_to_tile_21_9_3),
		.in_wire_3_0(vertical_tile_21_9_to_tile_22_9_0),
		.in_wire_3_1(vertical_tile_21_9_to_tile_22_9_1),
		.in_wire_3_2(vertical_tile_21_9_to_tile_22_9_2),
		.in_wire_3_3(vertical_tile_21_9_to_tile_22_9_3),
		.out_wire_1_0(vertical_tile_22_9_to_tile_23_9_0),
		.out_wire_1_1(vertical_tile_22_9_to_tile_23_9_1),
		.out_wire_1_2(vertical_tile_22_9_to_tile_23_9_2),
		.out_wire_1_3(vertical_tile_22_9_to_tile_23_9_3),
		.in_wire_1_0(vertical_tile_23_9_to_tile_22_9_0),
		.in_wire_1_1(vertical_tile_23_9_to_tile_22_9_1),
		.in_wire_1_2(vertical_tile_23_9_to_tile_22_9_2),
		.in_wire_1_3(vertical_tile_23_9_to_tile_22_9_3),
		.out_wire_2_0(horizontal_tile_22_9_to_tile_22_8_0),
		.out_wire_2_1(horizontal_tile_22_9_to_tile_22_8_1),
		.out_wire_2_2(horizontal_tile_22_9_to_tile_22_8_2),
		.out_wire_2_3(horizontal_tile_22_9_to_tile_22_8_3),
		.in_wire_2_0(horizontal_tile_22_8_to_tile_22_9_0),
		.in_wire_2_1(horizontal_tile_22_8_to_tile_22_9_1),
		.in_wire_2_2(horizontal_tile_22_8_to_tile_22_9_2),
		.in_wire_2_3(horizontal_tile_22_8_to_tile_22_9_3),
		.out_wire_0_0(horizontal_tile_22_9_to_tile_22_10_0),
		.out_wire_0_1(horizontal_tile_22_9_to_tile_22_10_1),
		.out_wire_0_2(horizontal_tile_22_9_to_tile_22_10_2),
		.out_wire_0_3(horizontal_tile_22_9_to_tile_22_10_3),
		.in_wire_0_0(horizontal_tile_22_10_to_tile_22_9_0),
		.in_wire_0_1(horizontal_tile_22_10_to_tile_22_9_1),
		.in_wire_0_2(horizontal_tile_22_10_to_tile_22_9_2),
		.in_wire_0_3(horizontal_tile_22_10_to_tile_22_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(714)
	);

	pe_tile pe_tile_22_10(
		.out_wire_3_0(vertical_tile_22_10_to_tile_21_10_0),
		.out_wire_3_1(vertical_tile_22_10_to_tile_21_10_1),
		.out_wire_3_2(vertical_tile_22_10_to_tile_21_10_2),
		.out_wire_3_3(vertical_tile_22_10_to_tile_21_10_3),
		.in_wire_3_0(vertical_tile_21_10_to_tile_22_10_0),
		.in_wire_3_1(vertical_tile_21_10_to_tile_22_10_1),
		.in_wire_3_2(vertical_tile_21_10_to_tile_22_10_2),
		.in_wire_3_3(vertical_tile_21_10_to_tile_22_10_3),
		.out_wire_1_0(vertical_tile_22_10_to_tile_23_10_0),
		.out_wire_1_1(vertical_tile_22_10_to_tile_23_10_1),
		.out_wire_1_2(vertical_tile_22_10_to_tile_23_10_2),
		.out_wire_1_3(vertical_tile_22_10_to_tile_23_10_3),
		.in_wire_1_0(vertical_tile_23_10_to_tile_22_10_0),
		.in_wire_1_1(vertical_tile_23_10_to_tile_22_10_1),
		.in_wire_1_2(vertical_tile_23_10_to_tile_22_10_2),
		.in_wire_1_3(vertical_tile_23_10_to_tile_22_10_3),
		.out_wire_2_0(horizontal_tile_22_10_to_tile_22_9_0),
		.out_wire_2_1(horizontal_tile_22_10_to_tile_22_9_1),
		.out_wire_2_2(horizontal_tile_22_10_to_tile_22_9_2),
		.out_wire_2_3(horizontal_tile_22_10_to_tile_22_9_3),
		.in_wire_2_0(horizontal_tile_22_9_to_tile_22_10_0),
		.in_wire_2_1(horizontal_tile_22_9_to_tile_22_10_1),
		.in_wire_2_2(horizontal_tile_22_9_to_tile_22_10_2),
		.in_wire_2_3(horizontal_tile_22_9_to_tile_22_10_3),
		.out_wire_0_0(horizontal_tile_22_10_to_tile_22_11_0),
		.out_wire_0_1(horizontal_tile_22_10_to_tile_22_11_1),
		.out_wire_0_2(horizontal_tile_22_10_to_tile_22_11_2),
		.out_wire_0_3(horizontal_tile_22_10_to_tile_22_11_3),
		.in_wire_0_0(horizontal_tile_22_11_to_tile_22_10_0),
		.in_wire_0_1(horizontal_tile_22_11_to_tile_22_10_1),
		.in_wire_0_2(horizontal_tile_22_11_to_tile_22_10_2),
		.in_wire_0_3(horizontal_tile_22_11_to_tile_22_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(715)
	);

	pe_tile pe_tile_22_11(
		.out_wire_3_0(vertical_tile_22_11_to_tile_21_11_0),
		.out_wire_3_1(vertical_tile_22_11_to_tile_21_11_1),
		.out_wire_3_2(vertical_tile_22_11_to_tile_21_11_2),
		.out_wire_3_3(vertical_tile_22_11_to_tile_21_11_3),
		.in_wire_3_0(vertical_tile_21_11_to_tile_22_11_0),
		.in_wire_3_1(vertical_tile_21_11_to_tile_22_11_1),
		.in_wire_3_2(vertical_tile_21_11_to_tile_22_11_2),
		.in_wire_3_3(vertical_tile_21_11_to_tile_22_11_3),
		.out_wire_1_0(vertical_tile_22_11_to_tile_23_11_0),
		.out_wire_1_1(vertical_tile_22_11_to_tile_23_11_1),
		.out_wire_1_2(vertical_tile_22_11_to_tile_23_11_2),
		.out_wire_1_3(vertical_tile_22_11_to_tile_23_11_3),
		.in_wire_1_0(vertical_tile_23_11_to_tile_22_11_0),
		.in_wire_1_1(vertical_tile_23_11_to_tile_22_11_1),
		.in_wire_1_2(vertical_tile_23_11_to_tile_22_11_2),
		.in_wire_1_3(vertical_tile_23_11_to_tile_22_11_3),
		.out_wire_2_0(horizontal_tile_22_11_to_tile_22_10_0),
		.out_wire_2_1(horizontal_tile_22_11_to_tile_22_10_1),
		.out_wire_2_2(horizontal_tile_22_11_to_tile_22_10_2),
		.out_wire_2_3(horizontal_tile_22_11_to_tile_22_10_3),
		.in_wire_2_0(horizontal_tile_22_10_to_tile_22_11_0),
		.in_wire_2_1(horizontal_tile_22_10_to_tile_22_11_1),
		.in_wire_2_2(horizontal_tile_22_10_to_tile_22_11_2),
		.in_wire_2_3(horizontal_tile_22_10_to_tile_22_11_3),
		.out_wire_0_0(horizontal_tile_22_11_to_tile_22_12_0),
		.out_wire_0_1(horizontal_tile_22_11_to_tile_22_12_1),
		.out_wire_0_2(horizontal_tile_22_11_to_tile_22_12_2),
		.out_wire_0_3(horizontal_tile_22_11_to_tile_22_12_3),
		.in_wire_0_0(horizontal_tile_22_12_to_tile_22_11_0),
		.in_wire_0_1(horizontal_tile_22_12_to_tile_22_11_1),
		.in_wire_0_2(horizontal_tile_22_12_to_tile_22_11_2),
		.in_wire_0_3(horizontal_tile_22_12_to_tile_22_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(716)
	);

	pe_tile pe_tile_22_12(
		.out_wire_3_0(vertical_tile_22_12_to_tile_21_12_0),
		.out_wire_3_1(vertical_tile_22_12_to_tile_21_12_1),
		.out_wire_3_2(vertical_tile_22_12_to_tile_21_12_2),
		.out_wire_3_3(vertical_tile_22_12_to_tile_21_12_3),
		.in_wire_3_0(vertical_tile_21_12_to_tile_22_12_0),
		.in_wire_3_1(vertical_tile_21_12_to_tile_22_12_1),
		.in_wire_3_2(vertical_tile_21_12_to_tile_22_12_2),
		.in_wire_3_3(vertical_tile_21_12_to_tile_22_12_3),
		.out_wire_1_0(vertical_tile_22_12_to_tile_23_12_0),
		.out_wire_1_1(vertical_tile_22_12_to_tile_23_12_1),
		.out_wire_1_2(vertical_tile_22_12_to_tile_23_12_2),
		.out_wire_1_3(vertical_tile_22_12_to_tile_23_12_3),
		.in_wire_1_0(vertical_tile_23_12_to_tile_22_12_0),
		.in_wire_1_1(vertical_tile_23_12_to_tile_22_12_1),
		.in_wire_1_2(vertical_tile_23_12_to_tile_22_12_2),
		.in_wire_1_3(vertical_tile_23_12_to_tile_22_12_3),
		.out_wire_2_0(horizontal_tile_22_12_to_tile_22_11_0),
		.out_wire_2_1(horizontal_tile_22_12_to_tile_22_11_1),
		.out_wire_2_2(horizontal_tile_22_12_to_tile_22_11_2),
		.out_wire_2_3(horizontal_tile_22_12_to_tile_22_11_3),
		.in_wire_2_0(horizontal_tile_22_11_to_tile_22_12_0),
		.in_wire_2_1(horizontal_tile_22_11_to_tile_22_12_1),
		.in_wire_2_2(horizontal_tile_22_11_to_tile_22_12_2),
		.in_wire_2_3(horizontal_tile_22_11_to_tile_22_12_3),
		.out_wire_0_0(horizontal_tile_22_12_to_tile_22_13_0),
		.out_wire_0_1(horizontal_tile_22_12_to_tile_22_13_1),
		.out_wire_0_2(horizontal_tile_22_12_to_tile_22_13_2),
		.out_wire_0_3(horizontal_tile_22_12_to_tile_22_13_3),
		.in_wire_0_0(horizontal_tile_22_13_to_tile_22_12_0),
		.in_wire_0_1(horizontal_tile_22_13_to_tile_22_12_1),
		.in_wire_0_2(horizontal_tile_22_13_to_tile_22_12_2),
		.in_wire_0_3(horizontal_tile_22_13_to_tile_22_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(717)
	);

	pe_tile pe_tile_22_13(
		.out_wire_3_0(vertical_tile_22_13_to_tile_21_13_0),
		.out_wire_3_1(vertical_tile_22_13_to_tile_21_13_1),
		.out_wire_3_2(vertical_tile_22_13_to_tile_21_13_2),
		.out_wire_3_3(vertical_tile_22_13_to_tile_21_13_3),
		.in_wire_3_0(vertical_tile_21_13_to_tile_22_13_0),
		.in_wire_3_1(vertical_tile_21_13_to_tile_22_13_1),
		.in_wire_3_2(vertical_tile_21_13_to_tile_22_13_2),
		.in_wire_3_3(vertical_tile_21_13_to_tile_22_13_3),
		.out_wire_1_0(vertical_tile_22_13_to_tile_23_13_0),
		.out_wire_1_1(vertical_tile_22_13_to_tile_23_13_1),
		.out_wire_1_2(vertical_tile_22_13_to_tile_23_13_2),
		.out_wire_1_3(vertical_tile_22_13_to_tile_23_13_3),
		.in_wire_1_0(vertical_tile_23_13_to_tile_22_13_0),
		.in_wire_1_1(vertical_tile_23_13_to_tile_22_13_1),
		.in_wire_1_2(vertical_tile_23_13_to_tile_22_13_2),
		.in_wire_1_3(vertical_tile_23_13_to_tile_22_13_3),
		.out_wire_2_0(horizontal_tile_22_13_to_tile_22_12_0),
		.out_wire_2_1(horizontal_tile_22_13_to_tile_22_12_1),
		.out_wire_2_2(horizontal_tile_22_13_to_tile_22_12_2),
		.out_wire_2_3(horizontal_tile_22_13_to_tile_22_12_3),
		.in_wire_2_0(horizontal_tile_22_12_to_tile_22_13_0),
		.in_wire_2_1(horizontal_tile_22_12_to_tile_22_13_1),
		.in_wire_2_2(horizontal_tile_22_12_to_tile_22_13_2),
		.in_wire_2_3(horizontal_tile_22_12_to_tile_22_13_3),
		.out_wire_0_0(horizontal_tile_22_13_to_tile_22_14_0),
		.out_wire_0_1(horizontal_tile_22_13_to_tile_22_14_1),
		.out_wire_0_2(horizontal_tile_22_13_to_tile_22_14_2),
		.out_wire_0_3(horizontal_tile_22_13_to_tile_22_14_3),
		.in_wire_0_0(horizontal_tile_22_14_to_tile_22_13_0),
		.in_wire_0_1(horizontal_tile_22_14_to_tile_22_13_1),
		.in_wire_0_2(horizontal_tile_22_14_to_tile_22_13_2),
		.in_wire_0_3(horizontal_tile_22_14_to_tile_22_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(718)
	);

	pe_tile pe_tile_22_14(
		.out_wire_3_0(vertical_tile_22_14_to_tile_21_14_0),
		.out_wire_3_1(vertical_tile_22_14_to_tile_21_14_1),
		.out_wire_3_2(vertical_tile_22_14_to_tile_21_14_2),
		.out_wire_3_3(vertical_tile_22_14_to_tile_21_14_3),
		.in_wire_3_0(vertical_tile_21_14_to_tile_22_14_0),
		.in_wire_3_1(vertical_tile_21_14_to_tile_22_14_1),
		.in_wire_3_2(vertical_tile_21_14_to_tile_22_14_2),
		.in_wire_3_3(vertical_tile_21_14_to_tile_22_14_3),
		.out_wire_1_0(vertical_tile_22_14_to_tile_23_14_0),
		.out_wire_1_1(vertical_tile_22_14_to_tile_23_14_1),
		.out_wire_1_2(vertical_tile_22_14_to_tile_23_14_2),
		.out_wire_1_3(vertical_tile_22_14_to_tile_23_14_3),
		.in_wire_1_0(vertical_tile_23_14_to_tile_22_14_0),
		.in_wire_1_1(vertical_tile_23_14_to_tile_22_14_1),
		.in_wire_1_2(vertical_tile_23_14_to_tile_22_14_2),
		.in_wire_1_3(vertical_tile_23_14_to_tile_22_14_3),
		.out_wire_2_0(horizontal_tile_22_14_to_tile_22_13_0),
		.out_wire_2_1(horizontal_tile_22_14_to_tile_22_13_1),
		.out_wire_2_2(horizontal_tile_22_14_to_tile_22_13_2),
		.out_wire_2_3(horizontal_tile_22_14_to_tile_22_13_3),
		.in_wire_2_0(horizontal_tile_22_13_to_tile_22_14_0),
		.in_wire_2_1(horizontal_tile_22_13_to_tile_22_14_1),
		.in_wire_2_2(horizontal_tile_22_13_to_tile_22_14_2),
		.in_wire_2_3(horizontal_tile_22_13_to_tile_22_14_3),
		.out_wire_0_0(horizontal_tile_22_14_to_tile_22_15_0),
		.out_wire_0_1(horizontal_tile_22_14_to_tile_22_15_1),
		.out_wire_0_2(horizontal_tile_22_14_to_tile_22_15_2),
		.out_wire_0_3(horizontal_tile_22_14_to_tile_22_15_3),
		.in_wire_0_0(horizontal_tile_22_15_to_tile_22_14_0),
		.in_wire_0_1(horizontal_tile_22_15_to_tile_22_14_1),
		.in_wire_0_2(horizontal_tile_22_15_to_tile_22_14_2),
		.in_wire_0_3(horizontal_tile_22_15_to_tile_22_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(719)
	);

	pe_tile pe_tile_22_15(
		.out_wire_3_0(vertical_tile_22_15_to_tile_21_15_0),
		.out_wire_3_1(vertical_tile_22_15_to_tile_21_15_1),
		.out_wire_3_2(vertical_tile_22_15_to_tile_21_15_2),
		.out_wire_3_3(vertical_tile_22_15_to_tile_21_15_3),
		.in_wire_3_0(vertical_tile_21_15_to_tile_22_15_0),
		.in_wire_3_1(vertical_tile_21_15_to_tile_22_15_1),
		.in_wire_3_2(vertical_tile_21_15_to_tile_22_15_2),
		.in_wire_3_3(vertical_tile_21_15_to_tile_22_15_3),
		.out_wire_1_0(vertical_tile_22_15_to_tile_23_15_0),
		.out_wire_1_1(vertical_tile_22_15_to_tile_23_15_1),
		.out_wire_1_2(vertical_tile_22_15_to_tile_23_15_2),
		.out_wire_1_3(vertical_tile_22_15_to_tile_23_15_3),
		.in_wire_1_0(vertical_tile_23_15_to_tile_22_15_0),
		.in_wire_1_1(vertical_tile_23_15_to_tile_22_15_1),
		.in_wire_1_2(vertical_tile_23_15_to_tile_22_15_2),
		.in_wire_1_3(vertical_tile_23_15_to_tile_22_15_3),
		.out_wire_2_0(horizontal_tile_22_15_to_tile_22_14_0),
		.out_wire_2_1(horizontal_tile_22_15_to_tile_22_14_1),
		.out_wire_2_2(horizontal_tile_22_15_to_tile_22_14_2),
		.out_wire_2_3(horizontal_tile_22_15_to_tile_22_14_3),
		.in_wire_2_0(horizontal_tile_22_14_to_tile_22_15_0),
		.in_wire_2_1(horizontal_tile_22_14_to_tile_22_15_1),
		.in_wire_2_2(horizontal_tile_22_14_to_tile_22_15_2),
		.in_wire_2_3(horizontal_tile_22_14_to_tile_22_15_3),
		.out_wire_0_0(horizontal_tile_22_15_to_tile_22_16_0),
		.out_wire_0_1(horizontal_tile_22_15_to_tile_22_16_1),
		.out_wire_0_2(horizontal_tile_22_15_to_tile_22_16_2),
		.out_wire_0_3(horizontal_tile_22_15_to_tile_22_16_3),
		.in_wire_0_0(horizontal_tile_22_16_to_tile_22_15_0),
		.in_wire_0_1(horizontal_tile_22_16_to_tile_22_15_1),
		.in_wire_0_2(horizontal_tile_22_16_to_tile_22_15_2),
		.in_wire_0_3(horizontal_tile_22_16_to_tile_22_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(720)
	);

	pe_tile pe_tile_22_16(
		.out_wire_3_0(vertical_tile_22_16_to_tile_21_16_0),
		.out_wire_3_1(vertical_tile_22_16_to_tile_21_16_1),
		.out_wire_3_2(vertical_tile_22_16_to_tile_21_16_2),
		.out_wire_3_3(vertical_tile_22_16_to_tile_21_16_3),
		.in_wire_3_0(vertical_tile_21_16_to_tile_22_16_0),
		.in_wire_3_1(vertical_tile_21_16_to_tile_22_16_1),
		.in_wire_3_2(vertical_tile_21_16_to_tile_22_16_2),
		.in_wire_3_3(vertical_tile_21_16_to_tile_22_16_3),
		.out_wire_1_0(vertical_tile_22_16_to_tile_23_16_0),
		.out_wire_1_1(vertical_tile_22_16_to_tile_23_16_1),
		.out_wire_1_2(vertical_tile_22_16_to_tile_23_16_2),
		.out_wire_1_3(vertical_tile_22_16_to_tile_23_16_3),
		.in_wire_1_0(vertical_tile_23_16_to_tile_22_16_0),
		.in_wire_1_1(vertical_tile_23_16_to_tile_22_16_1),
		.in_wire_1_2(vertical_tile_23_16_to_tile_22_16_2),
		.in_wire_1_3(vertical_tile_23_16_to_tile_22_16_3),
		.out_wire_2_0(horizontal_tile_22_16_to_tile_22_15_0),
		.out_wire_2_1(horizontal_tile_22_16_to_tile_22_15_1),
		.out_wire_2_2(horizontal_tile_22_16_to_tile_22_15_2),
		.out_wire_2_3(horizontal_tile_22_16_to_tile_22_15_3),
		.in_wire_2_0(horizontal_tile_22_15_to_tile_22_16_0),
		.in_wire_2_1(horizontal_tile_22_15_to_tile_22_16_1),
		.in_wire_2_2(horizontal_tile_22_15_to_tile_22_16_2),
		.in_wire_2_3(horizontal_tile_22_15_to_tile_22_16_3),
		.out_wire_0_0(horizontal_tile_22_16_to_tile_22_17_0),
		.out_wire_0_1(horizontal_tile_22_16_to_tile_22_17_1),
		.out_wire_0_2(horizontal_tile_22_16_to_tile_22_17_2),
		.out_wire_0_3(horizontal_tile_22_16_to_tile_22_17_3),
		.in_wire_0_0(horizontal_tile_22_17_to_tile_22_16_0),
		.in_wire_0_1(horizontal_tile_22_17_to_tile_22_16_1),
		.in_wire_0_2(horizontal_tile_22_17_to_tile_22_16_2),
		.in_wire_0_3(horizontal_tile_22_17_to_tile_22_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(721)
	);

	pe_tile pe_tile_22_17(
		.out_wire_3_0(vertical_tile_22_17_to_tile_21_17_0),
		.out_wire_3_1(vertical_tile_22_17_to_tile_21_17_1),
		.out_wire_3_2(vertical_tile_22_17_to_tile_21_17_2),
		.out_wire_3_3(vertical_tile_22_17_to_tile_21_17_3),
		.in_wire_3_0(vertical_tile_21_17_to_tile_22_17_0),
		.in_wire_3_1(vertical_tile_21_17_to_tile_22_17_1),
		.in_wire_3_2(vertical_tile_21_17_to_tile_22_17_2),
		.in_wire_3_3(vertical_tile_21_17_to_tile_22_17_3),
		.out_wire_1_0(vertical_tile_22_17_to_tile_23_17_0),
		.out_wire_1_1(vertical_tile_22_17_to_tile_23_17_1),
		.out_wire_1_2(vertical_tile_22_17_to_tile_23_17_2),
		.out_wire_1_3(vertical_tile_22_17_to_tile_23_17_3),
		.in_wire_1_0(vertical_tile_23_17_to_tile_22_17_0),
		.in_wire_1_1(vertical_tile_23_17_to_tile_22_17_1),
		.in_wire_1_2(vertical_tile_23_17_to_tile_22_17_2),
		.in_wire_1_3(vertical_tile_23_17_to_tile_22_17_3),
		.out_wire_2_0(horizontal_tile_22_17_to_tile_22_16_0),
		.out_wire_2_1(horizontal_tile_22_17_to_tile_22_16_1),
		.out_wire_2_2(horizontal_tile_22_17_to_tile_22_16_2),
		.out_wire_2_3(horizontal_tile_22_17_to_tile_22_16_3),
		.in_wire_2_0(horizontal_tile_22_16_to_tile_22_17_0),
		.in_wire_2_1(horizontal_tile_22_16_to_tile_22_17_1),
		.in_wire_2_2(horizontal_tile_22_16_to_tile_22_17_2),
		.in_wire_2_3(horizontal_tile_22_16_to_tile_22_17_3),
		.out_wire_0_0(horizontal_tile_22_17_to_tile_22_18_0),
		.out_wire_0_1(horizontal_tile_22_17_to_tile_22_18_1),
		.out_wire_0_2(horizontal_tile_22_17_to_tile_22_18_2),
		.out_wire_0_3(horizontal_tile_22_17_to_tile_22_18_3),
		.in_wire_0_0(horizontal_tile_22_18_to_tile_22_17_0),
		.in_wire_0_1(horizontal_tile_22_18_to_tile_22_17_1),
		.in_wire_0_2(horizontal_tile_22_18_to_tile_22_17_2),
		.in_wire_0_3(horizontal_tile_22_18_to_tile_22_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(722)
	);

	pe_tile pe_tile_22_18(
		.out_wire_3_0(vertical_tile_22_18_to_tile_21_18_0),
		.out_wire_3_1(vertical_tile_22_18_to_tile_21_18_1),
		.out_wire_3_2(vertical_tile_22_18_to_tile_21_18_2),
		.out_wire_3_3(vertical_tile_22_18_to_tile_21_18_3),
		.in_wire_3_0(vertical_tile_21_18_to_tile_22_18_0),
		.in_wire_3_1(vertical_tile_21_18_to_tile_22_18_1),
		.in_wire_3_2(vertical_tile_21_18_to_tile_22_18_2),
		.in_wire_3_3(vertical_tile_21_18_to_tile_22_18_3),
		.out_wire_1_0(vertical_tile_22_18_to_tile_23_18_0),
		.out_wire_1_1(vertical_tile_22_18_to_tile_23_18_1),
		.out_wire_1_2(vertical_tile_22_18_to_tile_23_18_2),
		.out_wire_1_3(vertical_tile_22_18_to_tile_23_18_3),
		.in_wire_1_0(vertical_tile_23_18_to_tile_22_18_0),
		.in_wire_1_1(vertical_tile_23_18_to_tile_22_18_1),
		.in_wire_1_2(vertical_tile_23_18_to_tile_22_18_2),
		.in_wire_1_3(vertical_tile_23_18_to_tile_22_18_3),
		.out_wire_2_0(horizontal_tile_22_18_to_tile_22_17_0),
		.out_wire_2_1(horizontal_tile_22_18_to_tile_22_17_1),
		.out_wire_2_2(horizontal_tile_22_18_to_tile_22_17_2),
		.out_wire_2_3(horizontal_tile_22_18_to_tile_22_17_3),
		.in_wire_2_0(horizontal_tile_22_17_to_tile_22_18_0),
		.in_wire_2_1(horizontal_tile_22_17_to_tile_22_18_1),
		.in_wire_2_2(horizontal_tile_22_17_to_tile_22_18_2),
		.in_wire_2_3(horizontal_tile_22_17_to_tile_22_18_3),
		.out_wire_0_0(horizontal_tile_22_18_to_tile_22_19_0),
		.out_wire_0_1(horizontal_tile_22_18_to_tile_22_19_1),
		.out_wire_0_2(horizontal_tile_22_18_to_tile_22_19_2),
		.out_wire_0_3(horizontal_tile_22_18_to_tile_22_19_3),
		.in_wire_0_0(horizontal_tile_22_19_to_tile_22_18_0),
		.in_wire_0_1(horizontal_tile_22_19_to_tile_22_18_1),
		.in_wire_0_2(horizontal_tile_22_19_to_tile_22_18_2),
		.in_wire_0_3(horizontal_tile_22_19_to_tile_22_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(723)
	);

	pe_tile pe_tile_22_19(
		.out_wire_3_0(vertical_tile_22_19_to_tile_21_19_0),
		.out_wire_3_1(vertical_tile_22_19_to_tile_21_19_1),
		.out_wire_3_2(vertical_tile_22_19_to_tile_21_19_2),
		.out_wire_3_3(vertical_tile_22_19_to_tile_21_19_3),
		.in_wire_3_0(vertical_tile_21_19_to_tile_22_19_0),
		.in_wire_3_1(vertical_tile_21_19_to_tile_22_19_1),
		.in_wire_3_2(vertical_tile_21_19_to_tile_22_19_2),
		.in_wire_3_3(vertical_tile_21_19_to_tile_22_19_3),
		.out_wire_1_0(vertical_tile_22_19_to_tile_23_19_0),
		.out_wire_1_1(vertical_tile_22_19_to_tile_23_19_1),
		.out_wire_1_2(vertical_tile_22_19_to_tile_23_19_2),
		.out_wire_1_3(vertical_tile_22_19_to_tile_23_19_3),
		.in_wire_1_0(vertical_tile_23_19_to_tile_22_19_0),
		.in_wire_1_1(vertical_tile_23_19_to_tile_22_19_1),
		.in_wire_1_2(vertical_tile_23_19_to_tile_22_19_2),
		.in_wire_1_3(vertical_tile_23_19_to_tile_22_19_3),
		.out_wire_2_0(horizontal_tile_22_19_to_tile_22_18_0),
		.out_wire_2_1(horizontal_tile_22_19_to_tile_22_18_1),
		.out_wire_2_2(horizontal_tile_22_19_to_tile_22_18_2),
		.out_wire_2_3(horizontal_tile_22_19_to_tile_22_18_3),
		.in_wire_2_0(horizontal_tile_22_18_to_tile_22_19_0),
		.in_wire_2_1(horizontal_tile_22_18_to_tile_22_19_1),
		.in_wire_2_2(horizontal_tile_22_18_to_tile_22_19_2),
		.in_wire_2_3(horizontal_tile_22_18_to_tile_22_19_3),
		.out_wire_0_0(horizontal_tile_22_19_to_tile_22_20_0),
		.out_wire_0_1(horizontal_tile_22_19_to_tile_22_20_1),
		.out_wire_0_2(horizontal_tile_22_19_to_tile_22_20_2),
		.out_wire_0_3(horizontal_tile_22_19_to_tile_22_20_3),
		.in_wire_0_0(horizontal_tile_22_20_to_tile_22_19_0),
		.in_wire_0_1(horizontal_tile_22_20_to_tile_22_19_1),
		.in_wire_0_2(horizontal_tile_22_20_to_tile_22_19_2),
		.in_wire_0_3(horizontal_tile_22_20_to_tile_22_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(724)
	);

	pe_tile pe_tile_22_20(
		.out_wire_3_0(vertical_tile_22_20_to_tile_21_20_0),
		.out_wire_3_1(vertical_tile_22_20_to_tile_21_20_1),
		.out_wire_3_2(vertical_tile_22_20_to_tile_21_20_2),
		.out_wire_3_3(vertical_tile_22_20_to_tile_21_20_3),
		.in_wire_3_0(vertical_tile_21_20_to_tile_22_20_0),
		.in_wire_3_1(vertical_tile_21_20_to_tile_22_20_1),
		.in_wire_3_2(vertical_tile_21_20_to_tile_22_20_2),
		.in_wire_3_3(vertical_tile_21_20_to_tile_22_20_3),
		.out_wire_1_0(vertical_tile_22_20_to_tile_23_20_0),
		.out_wire_1_1(vertical_tile_22_20_to_tile_23_20_1),
		.out_wire_1_2(vertical_tile_22_20_to_tile_23_20_2),
		.out_wire_1_3(vertical_tile_22_20_to_tile_23_20_3),
		.in_wire_1_0(vertical_tile_23_20_to_tile_22_20_0),
		.in_wire_1_1(vertical_tile_23_20_to_tile_22_20_1),
		.in_wire_1_2(vertical_tile_23_20_to_tile_22_20_2),
		.in_wire_1_3(vertical_tile_23_20_to_tile_22_20_3),
		.out_wire_2_0(horizontal_tile_22_20_to_tile_22_19_0),
		.out_wire_2_1(horizontal_tile_22_20_to_tile_22_19_1),
		.out_wire_2_2(horizontal_tile_22_20_to_tile_22_19_2),
		.out_wire_2_3(horizontal_tile_22_20_to_tile_22_19_3),
		.in_wire_2_0(horizontal_tile_22_19_to_tile_22_20_0),
		.in_wire_2_1(horizontal_tile_22_19_to_tile_22_20_1),
		.in_wire_2_2(horizontal_tile_22_19_to_tile_22_20_2),
		.in_wire_2_3(horizontal_tile_22_19_to_tile_22_20_3),
		.out_wire_0_0(horizontal_tile_22_20_to_tile_22_21_0),
		.out_wire_0_1(horizontal_tile_22_20_to_tile_22_21_1),
		.out_wire_0_2(horizontal_tile_22_20_to_tile_22_21_2),
		.out_wire_0_3(horizontal_tile_22_20_to_tile_22_21_3),
		.in_wire_0_0(horizontal_tile_22_21_to_tile_22_20_0),
		.in_wire_0_1(horizontal_tile_22_21_to_tile_22_20_1),
		.in_wire_0_2(horizontal_tile_22_21_to_tile_22_20_2),
		.in_wire_0_3(horizontal_tile_22_21_to_tile_22_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(725)
	);

	pe_tile pe_tile_22_21(
		.out_wire_3_0(vertical_tile_22_21_to_tile_21_21_0),
		.out_wire_3_1(vertical_tile_22_21_to_tile_21_21_1),
		.out_wire_3_2(vertical_tile_22_21_to_tile_21_21_2),
		.out_wire_3_3(vertical_tile_22_21_to_tile_21_21_3),
		.in_wire_3_0(vertical_tile_21_21_to_tile_22_21_0),
		.in_wire_3_1(vertical_tile_21_21_to_tile_22_21_1),
		.in_wire_3_2(vertical_tile_21_21_to_tile_22_21_2),
		.in_wire_3_3(vertical_tile_21_21_to_tile_22_21_3),
		.out_wire_1_0(vertical_tile_22_21_to_tile_23_21_0),
		.out_wire_1_1(vertical_tile_22_21_to_tile_23_21_1),
		.out_wire_1_2(vertical_tile_22_21_to_tile_23_21_2),
		.out_wire_1_3(vertical_tile_22_21_to_tile_23_21_3),
		.in_wire_1_0(vertical_tile_23_21_to_tile_22_21_0),
		.in_wire_1_1(vertical_tile_23_21_to_tile_22_21_1),
		.in_wire_1_2(vertical_tile_23_21_to_tile_22_21_2),
		.in_wire_1_3(vertical_tile_23_21_to_tile_22_21_3),
		.out_wire_2_0(horizontal_tile_22_21_to_tile_22_20_0),
		.out_wire_2_1(horizontal_tile_22_21_to_tile_22_20_1),
		.out_wire_2_2(horizontal_tile_22_21_to_tile_22_20_2),
		.out_wire_2_3(horizontal_tile_22_21_to_tile_22_20_3),
		.in_wire_2_0(horizontal_tile_22_20_to_tile_22_21_0),
		.in_wire_2_1(horizontal_tile_22_20_to_tile_22_21_1),
		.in_wire_2_2(horizontal_tile_22_20_to_tile_22_21_2),
		.in_wire_2_3(horizontal_tile_22_20_to_tile_22_21_3),
		.out_wire_0_0(horizontal_tile_22_21_to_tile_22_22_0),
		.out_wire_0_1(horizontal_tile_22_21_to_tile_22_22_1),
		.out_wire_0_2(horizontal_tile_22_21_to_tile_22_22_2),
		.out_wire_0_3(horizontal_tile_22_21_to_tile_22_22_3),
		.in_wire_0_0(horizontal_tile_22_22_to_tile_22_21_0),
		.in_wire_0_1(horizontal_tile_22_22_to_tile_22_21_1),
		.in_wire_0_2(horizontal_tile_22_22_to_tile_22_21_2),
		.in_wire_0_3(horizontal_tile_22_22_to_tile_22_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(726)
	);

	pe_tile pe_tile_22_22(
		.out_wire_3_0(vertical_tile_22_22_to_tile_21_22_0),
		.out_wire_3_1(vertical_tile_22_22_to_tile_21_22_1),
		.out_wire_3_2(vertical_tile_22_22_to_tile_21_22_2),
		.out_wire_3_3(vertical_tile_22_22_to_tile_21_22_3),
		.in_wire_3_0(vertical_tile_21_22_to_tile_22_22_0),
		.in_wire_3_1(vertical_tile_21_22_to_tile_22_22_1),
		.in_wire_3_2(vertical_tile_21_22_to_tile_22_22_2),
		.in_wire_3_3(vertical_tile_21_22_to_tile_22_22_3),
		.out_wire_1_0(vertical_tile_22_22_to_tile_23_22_0),
		.out_wire_1_1(vertical_tile_22_22_to_tile_23_22_1),
		.out_wire_1_2(vertical_tile_22_22_to_tile_23_22_2),
		.out_wire_1_3(vertical_tile_22_22_to_tile_23_22_3),
		.in_wire_1_0(vertical_tile_23_22_to_tile_22_22_0),
		.in_wire_1_1(vertical_tile_23_22_to_tile_22_22_1),
		.in_wire_1_2(vertical_tile_23_22_to_tile_22_22_2),
		.in_wire_1_3(vertical_tile_23_22_to_tile_22_22_3),
		.out_wire_2_0(horizontal_tile_22_22_to_tile_22_21_0),
		.out_wire_2_1(horizontal_tile_22_22_to_tile_22_21_1),
		.out_wire_2_2(horizontal_tile_22_22_to_tile_22_21_2),
		.out_wire_2_3(horizontal_tile_22_22_to_tile_22_21_3),
		.in_wire_2_0(horizontal_tile_22_21_to_tile_22_22_0),
		.in_wire_2_1(horizontal_tile_22_21_to_tile_22_22_1),
		.in_wire_2_2(horizontal_tile_22_21_to_tile_22_22_2),
		.in_wire_2_3(horizontal_tile_22_21_to_tile_22_22_3),
		.out_wire_0_0(horizontal_tile_22_22_to_tile_22_23_0),
		.out_wire_0_1(horizontal_tile_22_22_to_tile_22_23_1),
		.out_wire_0_2(horizontal_tile_22_22_to_tile_22_23_2),
		.out_wire_0_3(horizontal_tile_22_22_to_tile_22_23_3),
		.in_wire_0_0(horizontal_tile_22_23_to_tile_22_22_0),
		.in_wire_0_1(horizontal_tile_22_23_to_tile_22_22_1),
		.in_wire_0_2(horizontal_tile_22_23_to_tile_22_22_2),
		.in_wire_0_3(horizontal_tile_22_23_to_tile_22_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(727)
	);

	pe_tile pe_tile_22_23(
		.out_wire_3_0(vertical_tile_22_23_to_tile_21_23_0),
		.out_wire_3_1(vertical_tile_22_23_to_tile_21_23_1),
		.out_wire_3_2(vertical_tile_22_23_to_tile_21_23_2),
		.out_wire_3_3(vertical_tile_22_23_to_tile_21_23_3),
		.in_wire_3_0(vertical_tile_21_23_to_tile_22_23_0),
		.in_wire_3_1(vertical_tile_21_23_to_tile_22_23_1),
		.in_wire_3_2(vertical_tile_21_23_to_tile_22_23_2),
		.in_wire_3_3(vertical_tile_21_23_to_tile_22_23_3),
		.out_wire_1_0(vertical_tile_22_23_to_tile_23_23_0),
		.out_wire_1_1(vertical_tile_22_23_to_tile_23_23_1),
		.out_wire_1_2(vertical_tile_22_23_to_tile_23_23_2),
		.out_wire_1_3(vertical_tile_22_23_to_tile_23_23_3),
		.in_wire_1_0(vertical_tile_23_23_to_tile_22_23_0),
		.in_wire_1_1(vertical_tile_23_23_to_tile_22_23_1),
		.in_wire_1_2(vertical_tile_23_23_to_tile_22_23_2),
		.in_wire_1_3(vertical_tile_23_23_to_tile_22_23_3),
		.out_wire_2_0(horizontal_tile_22_23_to_tile_22_22_0),
		.out_wire_2_1(horizontal_tile_22_23_to_tile_22_22_1),
		.out_wire_2_2(horizontal_tile_22_23_to_tile_22_22_2),
		.out_wire_2_3(horizontal_tile_22_23_to_tile_22_22_3),
		.in_wire_2_0(horizontal_tile_22_22_to_tile_22_23_0),
		.in_wire_2_1(horizontal_tile_22_22_to_tile_22_23_1),
		.in_wire_2_2(horizontal_tile_22_22_to_tile_22_23_2),
		.in_wire_2_3(horizontal_tile_22_22_to_tile_22_23_3),
		.out_wire_0_0(horizontal_tile_22_23_to_tile_22_24_0),
		.out_wire_0_1(horizontal_tile_22_23_to_tile_22_24_1),
		.out_wire_0_2(horizontal_tile_22_23_to_tile_22_24_2),
		.out_wire_0_3(horizontal_tile_22_23_to_tile_22_24_3),
		.in_wire_0_0(horizontal_tile_22_24_to_tile_22_23_0),
		.in_wire_0_1(horizontal_tile_22_24_to_tile_22_23_1),
		.in_wire_0_2(horizontal_tile_22_24_to_tile_22_23_2),
		.in_wire_0_3(horizontal_tile_22_24_to_tile_22_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(728)
	);

	pe_tile pe_tile_22_24(
		.out_wire_3_0(vertical_tile_22_24_to_tile_21_24_0),
		.out_wire_3_1(vertical_tile_22_24_to_tile_21_24_1),
		.out_wire_3_2(vertical_tile_22_24_to_tile_21_24_2),
		.out_wire_3_3(vertical_tile_22_24_to_tile_21_24_3),
		.in_wire_3_0(vertical_tile_21_24_to_tile_22_24_0),
		.in_wire_3_1(vertical_tile_21_24_to_tile_22_24_1),
		.in_wire_3_2(vertical_tile_21_24_to_tile_22_24_2),
		.in_wire_3_3(vertical_tile_21_24_to_tile_22_24_3),
		.out_wire_1_0(vertical_tile_22_24_to_tile_23_24_0),
		.out_wire_1_1(vertical_tile_22_24_to_tile_23_24_1),
		.out_wire_1_2(vertical_tile_22_24_to_tile_23_24_2),
		.out_wire_1_3(vertical_tile_22_24_to_tile_23_24_3),
		.in_wire_1_0(vertical_tile_23_24_to_tile_22_24_0),
		.in_wire_1_1(vertical_tile_23_24_to_tile_22_24_1),
		.in_wire_1_2(vertical_tile_23_24_to_tile_22_24_2),
		.in_wire_1_3(vertical_tile_23_24_to_tile_22_24_3),
		.out_wire_2_0(horizontal_tile_22_24_to_tile_22_23_0),
		.out_wire_2_1(horizontal_tile_22_24_to_tile_22_23_1),
		.out_wire_2_2(horizontal_tile_22_24_to_tile_22_23_2),
		.out_wire_2_3(horizontal_tile_22_24_to_tile_22_23_3),
		.in_wire_2_0(horizontal_tile_22_23_to_tile_22_24_0),
		.in_wire_2_1(horizontal_tile_22_23_to_tile_22_24_1),
		.in_wire_2_2(horizontal_tile_22_23_to_tile_22_24_2),
		.in_wire_2_3(horizontal_tile_22_23_to_tile_22_24_3),
		.out_wire_0_0(horizontal_tile_22_24_to_tile_22_25_0),
		.out_wire_0_1(horizontal_tile_22_24_to_tile_22_25_1),
		.out_wire_0_2(horizontal_tile_22_24_to_tile_22_25_2),
		.out_wire_0_3(horizontal_tile_22_24_to_tile_22_25_3),
		.in_wire_0_0(horizontal_tile_22_25_to_tile_22_24_0),
		.in_wire_0_1(horizontal_tile_22_25_to_tile_22_24_1),
		.in_wire_0_2(horizontal_tile_22_25_to_tile_22_24_2),
		.in_wire_0_3(horizontal_tile_22_25_to_tile_22_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(729)
	);

	pe_tile pe_tile_22_25(
		.out_wire_3_0(vertical_tile_22_25_to_tile_21_25_0),
		.out_wire_3_1(vertical_tile_22_25_to_tile_21_25_1),
		.out_wire_3_2(vertical_tile_22_25_to_tile_21_25_2),
		.out_wire_3_3(vertical_tile_22_25_to_tile_21_25_3),
		.in_wire_3_0(vertical_tile_21_25_to_tile_22_25_0),
		.in_wire_3_1(vertical_tile_21_25_to_tile_22_25_1),
		.in_wire_3_2(vertical_tile_21_25_to_tile_22_25_2),
		.in_wire_3_3(vertical_tile_21_25_to_tile_22_25_3),
		.out_wire_1_0(vertical_tile_22_25_to_tile_23_25_0),
		.out_wire_1_1(vertical_tile_22_25_to_tile_23_25_1),
		.out_wire_1_2(vertical_tile_22_25_to_tile_23_25_2),
		.out_wire_1_3(vertical_tile_22_25_to_tile_23_25_3),
		.in_wire_1_0(vertical_tile_23_25_to_tile_22_25_0),
		.in_wire_1_1(vertical_tile_23_25_to_tile_22_25_1),
		.in_wire_1_2(vertical_tile_23_25_to_tile_22_25_2),
		.in_wire_1_3(vertical_tile_23_25_to_tile_22_25_3),
		.out_wire_2_0(horizontal_tile_22_25_to_tile_22_24_0),
		.out_wire_2_1(horizontal_tile_22_25_to_tile_22_24_1),
		.out_wire_2_2(horizontal_tile_22_25_to_tile_22_24_2),
		.out_wire_2_3(horizontal_tile_22_25_to_tile_22_24_3),
		.in_wire_2_0(horizontal_tile_22_24_to_tile_22_25_0),
		.in_wire_2_1(horizontal_tile_22_24_to_tile_22_25_1),
		.in_wire_2_2(horizontal_tile_22_24_to_tile_22_25_2),
		.in_wire_2_3(horizontal_tile_22_24_to_tile_22_25_3),
		.out_wire_0_0(horizontal_tile_22_25_to_tile_22_26_0),
		.out_wire_0_1(horizontal_tile_22_25_to_tile_22_26_1),
		.out_wire_0_2(horizontal_tile_22_25_to_tile_22_26_2),
		.out_wire_0_3(horizontal_tile_22_25_to_tile_22_26_3),
		.in_wire_0_0(horizontal_tile_22_26_to_tile_22_25_0),
		.in_wire_0_1(horizontal_tile_22_26_to_tile_22_25_1),
		.in_wire_0_2(horizontal_tile_22_26_to_tile_22_25_2),
		.in_wire_0_3(horizontal_tile_22_26_to_tile_22_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(730)
	);

	pe_tile pe_tile_22_26(
		.out_wire_3_0(vertical_tile_22_26_to_tile_21_26_0),
		.out_wire_3_1(vertical_tile_22_26_to_tile_21_26_1),
		.out_wire_3_2(vertical_tile_22_26_to_tile_21_26_2),
		.out_wire_3_3(vertical_tile_22_26_to_tile_21_26_3),
		.in_wire_3_0(vertical_tile_21_26_to_tile_22_26_0),
		.in_wire_3_1(vertical_tile_21_26_to_tile_22_26_1),
		.in_wire_3_2(vertical_tile_21_26_to_tile_22_26_2),
		.in_wire_3_3(vertical_tile_21_26_to_tile_22_26_3),
		.out_wire_1_0(vertical_tile_22_26_to_tile_23_26_0),
		.out_wire_1_1(vertical_tile_22_26_to_tile_23_26_1),
		.out_wire_1_2(vertical_tile_22_26_to_tile_23_26_2),
		.out_wire_1_3(vertical_tile_22_26_to_tile_23_26_3),
		.in_wire_1_0(vertical_tile_23_26_to_tile_22_26_0),
		.in_wire_1_1(vertical_tile_23_26_to_tile_22_26_1),
		.in_wire_1_2(vertical_tile_23_26_to_tile_22_26_2),
		.in_wire_1_3(vertical_tile_23_26_to_tile_22_26_3),
		.out_wire_2_0(horizontal_tile_22_26_to_tile_22_25_0),
		.out_wire_2_1(horizontal_tile_22_26_to_tile_22_25_1),
		.out_wire_2_2(horizontal_tile_22_26_to_tile_22_25_2),
		.out_wire_2_3(horizontal_tile_22_26_to_tile_22_25_3),
		.in_wire_2_0(horizontal_tile_22_25_to_tile_22_26_0),
		.in_wire_2_1(horizontal_tile_22_25_to_tile_22_26_1),
		.in_wire_2_2(horizontal_tile_22_25_to_tile_22_26_2),
		.in_wire_2_3(horizontal_tile_22_25_to_tile_22_26_3),
		.out_wire_0_0(horizontal_tile_22_26_to_tile_22_27_0),
		.out_wire_0_1(horizontal_tile_22_26_to_tile_22_27_1),
		.out_wire_0_2(horizontal_tile_22_26_to_tile_22_27_2),
		.out_wire_0_3(horizontal_tile_22_26_to_tile_22_27_3),
		.in_wire_0_0(horizontal_tile_22_27_to_tile_22_26_0),
		.in_wire_0_1(horizontal_tile_22_27_to_tile_22_26_1),
		.in_wire_0_2(horizontal_tile_22_27_to_tile_22_26_2),
		.in_wire_0_3(horizontal_tile_22_27_to_tile_22_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(731)
	);

	pe_tile pe_tile_22_27(
		.out_wire_3_0(vertical_tile_22_27_to_tile_21_27_0),
		.out_wire_3_1(vertical_tile_22_27_to_tile_21_27_1),
		.out_wire_3_2(vertical_tile_22_27_to_tile_21_27_2),
		.out_wire_3_3(vertical_tile_22_27_to_tile_21_27_3),
		.in_wire_3_0(vertical_tile_21_27_to_tile_22_27_0),
		.in_wire_3_1(vertical_tile_21_27_to_tile_22_27_1),
		.in_wire_3_2(vertical_tile_21_27_to_tile_22_27_2),
		.in_wire_3_3(vertical_tile_21_27_to_tile_22_27_3),
		.out_wire_1_0(vertical_tile_22_27_to_tile_23_27_0),
		.out_wire_1_1(vertical_tile_22_27_to_tile_23_27_1),
		.out_wire_1_2(vertical_tile_22_27_to_tile_23_27_2),
		.out_wire_1_3(vertical_tile_22_27_to_tile_23_27_3),
		.in_wire_1_0(vertical_tile_23_27_to_tile_22_27_0),
		.in_wire_1_1(vertical_tile_23_27_to_tile_22_27_1),
		.in_wire_1_2(vertical_tile_23_27_to_tile_22_27_2),
		.in_wire_1_3(vertical_tile_23_27_to_tile_22_27_3),
		.out_wire_2_0(horizontal_tile_22_27_to_tile_22_26_0),
		.out_wire_2_1(horizontal_tile_22_27_to_tile_22_26_1),
		.out_wire_2_2(horizontal_tile_22_27_to_tile_22_26_2),
		.out_wire_2_3(horizontal_tile_22_27_to_tile_22_26_3),
		.in_wire_2_0(horizontal_tile_22_26_to_tile_22_27_0),
		.in_wire_2_1(horizontal_tile_22_26_to_tile_22_27_1),
		.in_wire_2_2(horizontal_tile_22_26_to_tile_22_27_2),
		.in_wire_2_3(horizontal_tile_22_26_to_tile_22_27_3),
		.out_wire_0_0(horizontal_tile_22_27_to_tile_22_28_0),
		.out_wire_0_1(horizontal_tile_22_27_to_tile_22_28_1),
		.out_wire_0_2(horizontal_tile_22_27_to_tile_22_28_2),
		.out_wire_0_3(horizontal_tile_22_27_to_tile_22_28_3),
		.in_wire_0_0(horizontal_tile_22_28_to_tile_22_27_0),
		.in_wire_0_1(horizontal_tile_22_28_to_tile_22_27_1),
		.in_wire_0_2(horizontal_tile_22_28_to_tile_22_27_2),
		.in_wire_0_3(horizontal_tile_22_28_to_tile_22_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(732)
	);

	pe_tile pe_tile_22_28(
		.out_wire_3_0(vertical_tile_22_28_to_tile_21_28_0),
		.out_wire_3_1(vertical_tile_22_28_to_tile_21_28_1),
		.out_wire_3_2(vertical_tile_22_28_to_tile_21_28_2),
		.out_wire_3_3(vertical_tile_22_28_to_tile_21_28_3),
		.in_wire_3_0(vertical_tile_21_28_to_tile_22_28_0),
		.in_wire_3_1(vertical_tile_21_28_to_tile_22_28_1),
		.in_wire_3_2(vertical_tile_21_28_to_tile_22_28_2),
		.in_wire_3_3(vertical_tile_21_28_to_tile_22_28_3),
		.out_wire_1_0(vertical_tile_22_28_to_tile_23_28_0),
		.out_wire_1_1(vertical_tile_22_28_to_tile_23_28_1),
		.out_wire_1_2(vertical_tile_22_28_to_tile_23_28_2),
		.out_wire_1_3(vertical_tile_22_28_to_tile_23_28_3),
		.in_wire_1_0(vertical_tile_23_28_to_tile_22_28_0),
		.in_wire_1_1(vertical_tile_23_28_to_tile_22_28_1),
		.in_wire_1_2(vertical_tile_23_28_to_tile_22_28_2),
		.in_wire_1_3(vertical_tile_23_28_to_tile_22_28_3),
		.out_wire_2_0(horizontal_tile_22_28_to_tile_22_27_0),
		.out_wire_2_1(horizontal_tile_22_28_to_tile_22_27_1),
		.out_wire_2_2(horizontal_tile_22_28_to_tile_22_27_2),
		.out_wire_2_3(horizontal_tile_22_28_to_tile_22_27_3),
		.in_wire_2_0(horizontal_tile_22_27_to_tile_22_28_0),
		.in_wire_2_1(horizontal_tile_22_27_to_tile_22_28_1),
		.in_wire_2_2(horizontal_tile_22_27_to_tile_22_28_2),
		.in_wire_2_3(horizontal_tile_22_27_to_tile_22_28_3),
		.out_wire_0_0(horizontal_tile_22_28_to_tile_22_29_0),
		.out_wire_0_1(horizontal_tile_22_28_to_tile_22_29_1),
		.out_wire_0_2(horizontal_tile_22_28_to_tile_22_29_2),
		.out_wire_0_3(horizontal_tile_22_28_to_tile_22_29_3),
		.in_wire_0_0(horizontal_tile_22_29_to_tile_22_28_0),
		.in_wire_0_1(horizontal_tile_22_29_to_tile_22_28_1),
		.in_wire_0_2(horizontal_tile_22_29_to_tile_22_28_2),
		.in_wire_0_3(horizontal_tile_22_29_to_tile_22_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(733)
	);

	pe_tile pe_tile_22_29(
		.out_wire_3_0(vertical_tile_22_29_to_tile_21_29_0),
		.out_wire_3_1(vertical_tile_22_29_to_tile_21_29_1),
		.out_wire_3_2(vertical_tile_22_29_to_tile_21_29_2),
		.out_wire_3_3(vertical_tile_22_29_to_tile_21_29_3),
		.in_wire_3_0(vertical_tile_21_29_to_tile_22_29_0),
		.in_wire_3_1(vertical_tile_21_29_to_tile_22_29_1),
		.in_wire_3_2(vertical_tile_21_29_to_tile_22_29_2),
		.in_wire_3_3(vertical_tile_21_29_to_tile_22_29_3),
		.out_wire_1_0(vertical_tile_22_29_to_tile_23_29_0),
		.out_wire_1_1(vertical_tile_22_29_to_tile_23_29_1),
		.out_wire_1_2(vertical_tile_22_29_to_tile_23_29_2),
		.out_wire_1_3(vertical_tile_22_29_to_tile_23_29_3),
		.in_wire_1_0(vertical_tile_23_29_to_tile_22_29_0),
		.in_wire_1_1(vertical_tile_23_29_to_tile_22_29_1),
		.in_wire_1_2(vertical_tile_23_29_to_tile_22_29_2),
		.in_wire_1_3(vertical_tile_23_29_to_tile_22_29_3),
		.out_wire_2_0(horizontal_tile_22_29_to_tile_22_28_0),
		.out_wire_2_1(horizontal_tile_22_29_to_tile_22_28_1),
		.out_wire_2_2(horizontal_tile_22_29_to_tile_22_28_2),
		.out_wire_2_3(horizontal_tile_22_29_to_tile_22_28_3),
		.in_wire_2_0(horizontal_tile_22_28_to_tile_22_29_0),
		.in_wire_2_1(horizontal_tile_22_28_to_tile_22_29_1),
		.in_wire_2_2(horizontal_tile_22_28_to_tile_22_29_2),
		.in_wire_2_3(horizontal_tile_22_28_to_tile_22_29_3),
		.out_wire_0_0(horizontal_tile_22_29_to_tile_22_30_0),
		.out_wire_0_1(horizontal_tile_22_29_to_tile_22_30_1),
		.out_wire_0_2(horizontal_tile_22_29_to_tile_22_30_2),
		.out_wire_0_3(horizontal_tile_22_29_to_tile_22_30_3),
		.in_wire_0_0(horizontal_tile_22_30_to_tile_22_29_0),
		.in_wire_0_1(horizontal_tile_22_30_to_tile_22_29_1),
		.in_wire_0_2(horizontal_tile_22_30_to_tile_22_29_2),
		.in_wire_0_3(horizontal_tile_22_30_to_tile_22_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(734)
	);

	pe_tile pe_tile_22_30(
		.out_wire_3_0(vertical_tile_22_30_to_tile_21_30_0),
		.out_wire_3_1(vertical_tile_22_30_to_tile_21_30_1),
		.out_wire_3_2(vertical_tile_22_30_to_tile_21_30_2),
		.out_wire_3_3(vertical_tile_22_30_to_tile_21_30_3),
		.in_wire_3_0(vertical_tile_21_30_to_tile_22_30_0),
		.in_wire_3_1(vertical_tile_21_30_to_tile_22_30_1),
		.in_wire_3_2(vertical_tile_21_30_to_tile_22_30_2),
		.in_wire_3_3(vertical_tile_21_30_to_tile_22_30_3),
		.out_wire_1_0(vertical_tile_22_30_to_tile_23_30_0),
		.out_wire_1_1(vertical_tile_22_30_to_tile_23_30_1),
		.out_wire_1_2(vertical_tile_22_30_to_tile_23_30_2),
		.out_wire_1_3(vertical_tile_22_30_to_tile_23_30_3),
		.in_wire_1_0(vertical_tile_23_30_to_tile_22_30_0),
		.in_wire_1_1(vertical_tile_23_30_to_tile_22_30_1),
		.in_wire_1_2(vertical_tile_23_30_to_tile_22_30_2),
		.in_wire_1_3(vertical_tile_23_30_to_tile_22_30_3),
		.out_wire_2_0(horizontal_tile_22_30_to_tile_22_29_0),
		.out_wire_2_1(horizontal_tile_22_30_to_tile_22_29_1),
		.out_wire_2_2(horizontal_tile_22_30_to_tile_22_29_2),
		.out_wire_2_3(horizontal_tile_22_30_to_tile_22_29_3),
		.in_wire_2_0(horizontal_tile_22_29_to_tile_22_30_0),
		.in_wire_2_1(horizontal_tile_22_29_to_tile_22_30_1),
		.in_wire_2_2(horizontal_tile_22_29_to_tile_22_30_2),
		.in_wire_2_3(horizontal_tile_22_29_to_tile_22_30_3),
		.out_wire_0_0(horizontal_tile_22_30_to_tile_22_31_0),
		.out_wire_0_1(horizontal_tile_22_30_to_tile_22_31_1),
		.out_wire_0_2(horizontal_tile_22_30_to_tile_22_31_2),
		.out_wire_0_3(horizontal_tile_22_30_to_tile_22_31_3),
		.in_wire_0_0(horizontal_tile_22_31_to_tile_22_30_0),
		.in_wire_0_1(horizontal_tile_22_31_to_tile_22_30_1),
		.in_wire_0_2(horizontal_tile_22_31_to_tile_22_30_2),
		.in_wire_0_3(horizontal_tile_22_31_to_tile_22_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(735)
	);

	pe_tile_right pe_tile_22_31(
		.out_wire_3_0(vertical_tile_22_31_to_tile_21_31_0),
		.out_wire_3_1(vertical_tile_22_31_to_tile_21_31_1),
		.out_wire_3_2(vertical_tile_22_31_to_tile_21_31_2),
		.out_wire_3_3(vertical_tile_22_31_to_tile_21_31_3),
		.in_wire_3_0(vertical_tile_21_31_to_tile_22_31_0),
		.in_wire_3_1(vertical_tile_21_31_to_tile_22_31_1),
		.in_wire_3_2(vertical_tile_21_31_to_tile_22_31_2),
		.in_wire_3_3(vertical_tile_21_31_to_tile_22_31_3),
		.out_wire_1_0(vertical_tile_22_31_to_tile_23_31_0),
		.out_wire_1_1(vertical_tile_22_31_to_tile_23_31_1),
		.out_wire_1_2(vertical_tile_22_31_to_tile_23_31_2),
		.out_wire_1_3(vertical_tile_22_31_to_tile_23_31_3),
		.in_wire_1_0(vertical_tile_23_31_to_tile_22_31_0),
		.in_wire_1_1(vertical_tile_23_31_to_tile_22_31_1),
		.in_wire_1_2(vertical_tile_23_31_to_tile_22_31_2),
		.in_wire_1_3(vertical_tile_23_31_to_tile_22_31_3),
		.out_wire_2_0(horizontal_tile_22_31_to_tile_22_30_0),
		.out_wire_2_1(horizontal_tile_22_31_to_tile_22_30_1),
		.out_wire_2_2(horizontal_tile_22_31_to_tile_22_30_2),
		.out_wire_2_3(horizontal_tile_22_31_to_tile_22_30_3),
		.in_wire_2_0(horizontal_tile_22_30_to_tile_22_31_0),
		.in_wire_2_1(horizontal_tile_22_30_to_tile_22_31_1),
		.in_wire_2_2(horizontal_tile_22_30_to_tile_22_31_2),
		.in_wire_2_3(horizontal_tile_22_30_to_tile_22_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(736)
	);

	pe_tile_left pe_tile_23_0(
		.out_wire_3_0(vertical_tile_23_0_to_tile_22_0_0),
		.out_wire_3_1(vertical_tile_23_0_to_tile_22_0_1),
		.out_wire_3_2(vertical_tile_23_0_to_tile_22_0_2),
		.out_wire_3_3(vertical_tile_23_0_to_tile_22_0_3),
		.in_wire_3_0(vertical_tile_22_0_to_tile_23_0_0),
		.in_wire_3_1(vertical_tile_22_0_to_tile_23_0_1),
		.in_wire_3_2(vertical_tile_22_0_to_tile_23_0_2),
		.in_wire_3_3(vertical_tile_22_0_to_tile_23_0_3),
		.out_wire_1_0(vertical_tile_23_0_to_tile_24_0_0),
		.out_wire_1_1(vertical_tile_23_0_to_tile_24_0_1),
		.out_wire_1_2(vertical_tile_23_0_to_tile_24_0_2),
		.out_wire_1_3(vertical_tile_23_0_to_tile_24_0_3),
		.in_wire_1_0(vertical_tile_24_0_to_tile_23_0_0),
		.in_wire_1_1(vertical_tile_24_0_to_tile_23_0_1),
		.in_wire_1_2(vertical_tile_24_0_to_tile_23_0_2),
		.in_wire_1_3(vertical_tile_24_0_to_tile_23_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_23_0_to_tile_23_1_0),
		.out_wire_0_1(horizontal_tile_23_0_to_tile_23_1_1),
		.out_wire_0_2(horizontal_tile_23_0_to_tile_23_1_2),
		.out_wire_0_3(horizontal_tile_23_0_to_tile_23_1_3),
		.in_wire_0_0(horizontal_tile_23_1_to_tile_23_0_0),
		.in_wire_0_1(horizontal_tile_23_1_to_tile_23_0_1),
		.in_wire_0_2(horizontal_tile_23_1_to_tile_23_0_2),
		.in_wire_0_3(horizontal_tile_23_1_to_tile_23_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(737)
	);

	pe_tile pe_tile_23_1(
		.out_wire_3_0(vertical_tile_23_1_to_tile_22_1_0),
		.out_wire_3_1(vertical_tile_23_1_to_tile_22_1_1),
		.out_wire_3_2(vertical_tile_23_1_to_tile_22_1_2),
		.out_wire_3_3(vertical_tile_23_1_to_tile_22_1_3),
		.in_wire_3_0(vertical_tile_22_1_to_tile_23_1_0),
		.in_wire_3_1(vertical_tile_22_1_to_tile_23_1_1),
		.in_wire_3_2(vertical_tile_22_1_to_tile_23_1_2),
		.in_wire_3_3(vertical_tile_22_1_to_tile_23_1_3),
		.out_wire_1_0(vertical_tile_23_1_to_tile_24_1_0),
		.out_wire_1_1(vertical_tile_23_1_to_tile_24_1_1),
		.out_wire_1_2(vertical_tile_23_1_to_tile_24_1_2),
		.out_wire_1_3(vertical_tile_23_1_to_tile_24_1_3),
		.in_wire_1_0(vertical_tile_24_1_to_tile_23_1_0),
		.in_wire_1_1(vertical_tile_24_1_to_tile_23_1_1),
		.in_wire_1_2(vertical_tile_24_1_to_tile_23_1_2),
		.in_wire_1_3(vertical_tile_24_1_to_tile_23_1_3),
		.out_wire_2_0(horizontal_tile_23_1_to_tile_23_0_0),
		.out_wire_2_1(horizontal_tile_23_1_to_tile_23_0_1),
		.out_wire_2_2(horizontal_tile_23_1_to_tile_23_0_2),
		.out_wire_2_3(horizontal_tile_23_1_to_tile_23_0_3),
		.in_wire_2_0(horizontal_tile_23_0_to_tile_23_1_0),
		.in_wire_2_1(horizontal_tile_23_0_to_tile_23_1_1),
		.in_wire_2_2(horizontal_tile_23_0_to_tile_23_1_2),
		.in_wire_2_3(horizontal_tile_23_0_to_tile_23_1_3),
		.out_wire_0_0(horizontal_tile_23_1_to_tile_23_2_0),
		.out_wire_0_1(horizontal_tile_23_1_to_tile_23_2_1),
		.out_wire_0_2(horizontal_tile_23_1_to_tile_23_2_2),
		.out_wire_0_3(horizontal_tile_23_1_to_tile_23_2_3),
		.in_wire_0_0(horizontal_tile_23_2_to_tile_23_1_0),
		.in_wire_0_1(horizontal_tile_23_2_to_tile_23_1_1),
		.in_wire_0_2(horizontal_tile_23_2_to_tile_23_1_2),
		.in_wire_0_3(horizontal_tile_23_2_to_tile_23_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(738)
	);

	pe_tile pe_tile_23_2(
		.out_wire_3_0(vertical_tile_23_2_to_tile_22_2_0),
		.out_wire_3_1(vertical_tile_23_2_to_tile_22_2_1),
		.out_wire_3_2(vertical_tile_23_2_to_tile_22_2_2),
		.out_wire_3_3(vertical_tile_23_2_to_tile_22_2_3),
		.in_wire_3_0(vertical_tile_22_2_to_tile_23_2_0),
		.in_wire_3_1(vertical_tile_22_2_to_tile_23_2_1),
		.in_wire_3_2(vertical_tile_22_2_to_tile_23_2_2),
		.in_wire_3_3(vertical_tile_22_2_to_tile_23_2_3),
		.out_wire_1_0(vertical_tile_23_2_to_tile_24_2_0),
		.out_wire_1_1(vertical_tile_23_2_to_tile_24_2_1),
		.out_wire_1_2(vertical_tile_23_2_to_tile_24_2_2),
		.out_wire_1_3(vertical_tile_23_2_to_tile_24_2_3),
		.in_wire_1_0(vertical_tile_24_2_to_tile_23_2_0),
		.in_wire_1_1(vertical_tile_24_2_to_tile_23_2_1),
		.in_wire_1_2(vertical_tile_24_2_to_tile_23_2_2),
		.in_wire_1_3(vertical_tile_24_2_to_tile_23_2_3),
		.out_wire_2_0(horizontal_tile_23_2_to_tile_23_1_0),
		.out_wire_2_1(horizontal_tile_23_2_to_tile_23_1_1),
		.out_wire_2_2(horizontal_tile_23_2_to_tile_23_1_2),
		.out_wire_2_3(horizontal_tile_23_2_to_tile_23_1_3),
		.in_wire_2_0(horizontal_tile_23_1_to_tile_23_2_0),
		.in_wire_2_1(horizontal_tile_23_1_to_tile_23_2_1),
		.in_wire_2_2(horizontal_tile_23_1_to_tile_23_2_2),
		.in_wire_2_3(horizontal_tile_23_1_to_tile_23_2_3),
		.out_wire_0_0(horizontal_tile_23_2_to_tile_23_3_0),
		.out_wire_0_1(horizontal_tile_23_2_to_tile_23_3_1),
		.out_wire_0_2(horizontal_tile_23_2_to_tile_23_3_2),
		.out_wire_0_3(horizontal_tile_23_2_to_tile_23_3_3),
		.in_wire_0_0(horizontal_tile_23_3_to_tile_23_2_0),
		.in_wire_0_1(horizontal_tile_23_3_to_tile_23_2_1),
		.in_wire_0_2(horizontal_tile_23_3_to_tile_23_2_2),
		.in_wire_0_3(horizontal_tile_23_3_to_tile_23_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(739)
	);

	pe_tile pe_tile_23_3(
		.out_wire_3_0(vertical_tile_23_3_to_tile_22_3_0),
		.out_wire_3_1(vertical_tile_23_3_to_tile_22_3_1),
		.out_wire_3_2(vertical_tile_23_3_to_tile_22_3_2),
		.out_wire_3_3(vertical_tile_23_3_to_tile_22_3_3),
		.in_wire_3_0(vertical_tile_22_3_to_tile_23_3_0),
		.in_wire_3_1(vertical_tile_22_3_to_tile_23_3_1),
		.in_wire_3_2(vertical_tile_22_3_to_tile_23_3_2),
		.in_wire_3_3(vertical_tile_22_3_to_tile_23_3_3),
		.out_wire_1_0(vertical_tile_23_3_to_tile_24_3_0),
		.out_wire_1_1(vertical_tile_23_3_to_tile_24_3_1),
		.out_wire_1_2(vertical_tile_23_3_to_tile_24_3_2),
		.out_wire_1_3(vertical_tile_23_3_to_tile_24_3_3),
		.in_wire_1_0(vertical_tile_24_3_to_tile_23_3_0),
		.in_wire_1_1(vertical_tile_24_3_to_tile_23_3_1),
		.in_wire_1_2(vertical_tile_24_3_to_tile_23_3_2),
		.in_wire_1_3(vertical_tile_24_3_to_tile_23_3_3),
		.out_wire_2_0(horizontal_tile_23_3_to_tile_23_2_0),
		.out_wire_2_1(horizontal_tile_23_3_to_tile_23_2_1),
		.out_wire_2_2(horizontal_tile_23_3_to_tile_23_2_2),
		.out_wire_2_3(horizontal_tile_23_3_to_tile_23_2_3),
		.in_wire_2_0(horizontal_tile_23_2_to_tile_23_3_0),
		.in_wire_2_1(horizontal_tile_23_2_to_tile_23_3_1),
		.in_wire_2_2(horizontal_tile_23_2_to_tile_23_3_2),
		.in_wire_2_3(horizontal_tile_23_2_to_tile_23_3_3),
		.out_wire_0_0(horizontal_tile_23_3_to_tile_23_4_0),
		.out_wire_0_1(horizontal_tile_23_3_to_tile_23_4_1),
		.out_wire_0_2(horizontal_tile_23_3_to_tile_23_4_2),
		.out_wire_0_3(horizontal_tile_23_3_to_tile_23_4_3),
		.in_wire_0_0(horizontal_tile_23_4_to_tile_23_3_0),
		.in_wire_0_1(horizontal_tile_23_4_to_tile_23_3_1),
		.in_wire_0_2(horizontal_tile_23_4_to_tile_23_3_2),
		.in_wire_0_3(horizontal_tile_23_4_to_tile_23_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(740)
	);

	pe_tile pe_tile_23_4(
		.out_wire_3_0(vertical_tile_23_4_to_tile_22_4_0),
		.out_wire_3_1(vertical_tile_23_4_to_tile_22_4_1),
		.out_wire_3_2(vertical_tile_23_4_to_tile_22_4_2),
		.out_wire_3_3(vertical_tile_23_4_to_tile_22_4_3),
		.in_wire_3_0(vertical_tile_22_4_to_tile_23_4_0),
		.in_wire_3_1(vertical_tile_22_4_to_tile_23_4_1),
		.in_wire_3_2(vertical_tile_22_4_to_tile_23_4_2),
		.in_wire_3_3(vertical_tile_22_4_to_tile_23_4_3),
		.out_wire_1_0(vertical_tile_23_4_to_tile_24_4_0),
		.out_wire_1_1(vertical_tile_23_4_to_tile_24_4_1),
		.out_wire_1_2(vertical_tile_23_4_to_tile_24_4_2),
		.out_wire_1_3(vertical_tile_23_4_to_tile_24_4_3),
		.in_wire_1_0(vertical_tile_24_4_to_tile_23_4_0),
		.in_wire_1_1(vertical_tile_24_4_to_tile_23_4_1),
		.in_wire_1_2(vertical_tile_24_4_to_tile_23_4_2),
		.in_wire_1_3(vertical_tile_24_4_to_tile_23_4_3),
		.out_wire_2_0(horizontal_tile_23_4_to_tile_23_3_0),
		.out_wire_2_1(horizontal_tile_23_4_to_tile_23_3_1),
		.out_wire_2_2(horizontal_tile_23_4_to_tile_23_3_2),
		.out_wire_2_3(horizontal_tile_23_4_to_tile_23_3_3),
		.in_wire_2_0(horizontal_tile_23_3_to_tile_23_4_0),
		.in_wire_2_1(horizontal_tile_23_3_to_tile_23_4_1),
		.in_wire_2_2(horizontal_tile_23_3_to_tile_23_4_2),
		.in_wire_2_3(horizontal_tile_23_3_to_tile_23_4_3),
		.out_wire_0_0(horizontal_tile_23_4_to_tile_23_5_0),
		.out_wire_0_1(horizontal_tile_23_4_to_tile_23_5_1),
		.out_wire_0_2(horizontal_tile_23_4_to_tile_23_5_2),
		.out_wire_0_3(horizontal_tile_23_4_to_tile_23_5_3),
		.in_wire_0_0(horizontal_tile_23_5_to_tile_23_4_0),
		.in_wire_0_1(horizontal_tile_23_5_to_tile_23_4_1),
		.in_wire_0_2(horizontal_tile_23_5_to_tile_23_4_2),
		.in_wire_0_3(horizontal_tile_23_5_to_tile_23_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(741)
	);

	pe_tile pe_tile_23_5(
		.out_wire_3_0(vertical_tile_23_5_to_tile_22_5_0),
		.out_wire_3_1(vertical_tile_23_5_to_tile_22_5_1),
		.out_wire_3_2(vertical_tile_23_5_to_tile_22_5_2),
		.out_wire_3_3(vertical_tile_23_5_to_tile_22_5_3),
		.in_wire_3_0(vertical_tile_22_5_to_tile_23_5_0),
		.in_wire_3_1(vertical_tile_22_5_to_tile_23_5_1),
		.in_wire_3_2(vertical_tile_22_5_to_tile_23_5_2),
		.in_wire_3_3(vertical_tile_22_5_to_tile_23_5_3),
		.out_wire_1_0(vertical_tile_23_5_to_tile_24_5_0),
		.out_wire_1_1(vertical_tile_23_5_to_tile_24_5_1),
		.out_wire_1_2(vertical_tile_23_5_to_tile_24_5_2),
		.out_wire_1_3(vertical_tile_23_5_to_tile_24_5_3),
		.in_wire_1_0(vertical_tile_24_5_to_tile_23_5_0),
		.in_wire_1_1(vertical_tile_24_5_to_tile_23_5_1),
		.in_wire_1_2(vertical_tile_24_5_to_tile_23_5_2),
		.in_wire_1_3(vertical_tile_24_5_to_tile_23_5_3),
		.out_wire_2_0(horizontal_tile_23_5_to_tile_23_4_0),
		.out_wire_2_1(horizontal_tile_23_5_to_tile_23_4_1),
		.out_wire_2_2(horizontal_tile_23_5_to_tile_23_4_2),
		.out_wire_2_3(horizontal_tile_23_5_to_tile_23_4_3),
		.in_wire_2_0(horizontal_tile_23_4_to_tile_23_5_0),
		.in_wire_2_1(horizontal_tile_23_4_to_tile_23_5_1),
		.in_wire_2_2(horizontal_tile_23_4_to_tile_23_5_2),
		.in_wire_2_3(horizontal_tile_23_4_to_tile_23_5_3),
		.out_wire_0_0(horizontal_tile_23_5_to_tile_23_6_0),
		.out_wire_0_1(horizontal_tile_23_5_to_tile_23_6_1),
		.out_wire_0_2(horizontal_tile_23_5_to_tile_23_6_2),
		.out_wire_0_3(horizontal_tile_23_5_to_tile_23_6_3),
		.in_wire_0_0(horizontal_tile_23_6_to_tile_23_5_0),
		.in_wire_0_1(horizontal_tile_23_6_to_tile_23_5_1),
		.in_wire_0_2(horizontal_tile_23_6_to_tile_23_5_2),
		.in_wire_0_3(horizontal_tile_23_6_to_tile_23_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(742)
	);

	pe_tile pe_tile_23_6(
		.out_wire_3_0(vertical_tile_23_6_to_tile_22_6_0),
		.out_wire_3_1(vertical_tile_23_6_to_tile_22_6_1),
		.out_wire_3_2(vertical_tile_23_6_to_tile_22_6_2),
		.out_wire_3_3(vertical_tile_23_6_to_tile_22_6_3),
		.in_wire_3_0(vertical_tile_22_6_to_tile_23_6_0),
		.in_wire_3_1(vertical_tile_22_6_to_tile_23_6_1),
		.in_wire_3_2(vertical_tile_22_6_to_tile_23_6_2),
		.in_wire_3_3(vertical_tile_22_6_to_tile_23_6_3),
		.out_wire_1_0(vertical_tile_23_6_to_tile_24_6_0),
		.out_wire_1_1(vertical_tile_23_6_to_tile_24_6_1),
		.out_wire_1_2(vertical_tile_23_6_to_tile_24_6_2),
		.out_wire_1_3(vertical_tile_23_6_to_tile_24_6_3),
		.in_wire_1_0(vertical_tile_24_6_to_tile_23_6_0),
		.in_wire_1_1(vertical_tile_24_6_to_tile_23_6_1),
		.in_wire_1_2(vertical_tile_24_6_to_tile_23_6_2),
		.in_wire_1_3(vertical_tile_24_6_to_tile_23_6_3),
		.out_wire_2_0(horizontal_tile_23_6_to_tile_23_5_0),
		.out_wire_2_1(horizontal_tile_23_6_to_tile_23_5_1),
		.out_wire_2_2(horizontal_tile_23_6_to_tile_23_5_2),
		.out_wire_2_3(horizontal_tile_23_6_to_tile_23_5_3),
		.in_wire_2_0(horizontal_tile_23_5_to_tile_23_6_0),
		.in_wire_2_1(horizontal_tile_23_5_to_tile_23_6_1),
		.in_wire_2_2(horizontal_tile_23_5_to_tile_23_6_2),
		.in_wire_2_3(horizontal_tile_23_5_to_tile_23_6_3),
		.out_wire_0_0(horizontal_tile_23_6_to_tile_23_7_0),
		.out_wire_0_1(horizontal_tile_23_6_to_tile_23_7_1),
		.out_wire_0_2(horizontal_tile_23_6_to_tile_23_7_2),
		.out_wire_0_3(horizontal_tile_23_6_to_tile_23_7_3),
		.in_wire_0_0(horizontal_tile_23_7_to_tile_23_6_0),
		.in_wire_0_1(horizontal_tile_23_7_to_tile_23_6_1),
		.in_wire_0_2(horizontal_tile_23_7_to_tile_23_6_2),
		.in_wire_0_3(horizontal_tile_23_7_to_tile_23_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(743)
	);

	pe_tile pe_tile_23_7(
		.out_wire_3_0(vertical_tile_23_7_to_tile_22_7_0),
		.out_wire_3_1(vertical_tile_23_7_to_tile_22_7_1),
		.out_wire_3_2(vertical_tile_23_7_to_tile_22_7_2),
		.out_wire_3_3(vertical_tile_23_7_to_tile_22_7_3),
		.in_wire_3_0(vertical_tile_22_7_to_tile_23_7_0),
		.in_wire_3_1(vertical_tile_22_7_to_tile_23_7_1),
		.in_wire_3_2(vertical_tile_22_7_to_tile_23_7_2),
		.in_wire_3_3(vertical_tile_22_7_to_tile_23_7_3),
		.out_wire_1_0(vertical_tile_23_7_to_tile_24_7_0),
		.out_wire_1_1(vertical_tile_23_7_to_tile_24_7_1),
		.out_wire_1_2(vertical_tile_23_7_to_tile_24_7_2),
		.out_wire_1_3(vertical_tile_23_7_to_tile_24_7_3),
		.in_wire_1_0(vertical_tile_24_7_to_tile_23_7_0),
		.in_wire_1_1(vertical_tile_24_7_to_tile_23_7_1),
		.in_wire_1_2(vertical_tile_24_7_to_tile_23_7_2),
		.in_wire_1_3(vertical_tile_24_7_to_tile_23_7_3),
		.out_wire_2_0(horizontal_tile_23_7_to_tile_23_6_0),
		.out_wire_2_1(horizontal_tile_23_7_to_tile_23_6_1),
		.out_wire_2_2(horizontal_tile_23_7_to_tile_23_6_2),
		.out_wire_2_3(horizontal_tile_23_7_to_tile_23_6_3),
		.in_wire_2_0(horizontal_tile_23_6_to_tile_23_7_0),
		.in_wire_2_1(horizontal_tile_23_6_to_tile_23_7_1),
		.in_wire_2_2(horizontal_tile_23_6_to_tile_23_7_2),
		.in_wire_2_3(horizontal_tile_23_6_to_tile_23_7_3),
		.out_wire_0_0(horizontal_tile_23_7_to_tile_23_8_0),
		.out_wire_0_1(horizontal_tile_23_7_to_tile_23_8_1),
		.out_wire_0_2(horizontal_tile_23_7_to_tile_23_8_2),
		.out_wire_0_3(horizontal_tile_23_7_to_tile_23_8_3),
		.in_wire_0_0(horizontal_tile_23_8_to_tile_23_7_0),
		.in_wire_0_1(horizontal_tile_23_8_to_tile_23_7_1),
		.in_wire_0_2(horizontal_tile_23_8_to_tile_23_7_2),
		.in_wire_0_3(horizontal_tile_23_8_to_tile_23_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(744)
	);

	pe_tile pe_tile_23_8(
		.out_wire_3_0(vertical_tile_23_8_to_tile_22_8_0),
		.out_wire_3_1(vertical_tile_23_8_to_tile_22_8_1),
		.out_wire_3_2(vertical_tile_23_8_to_tile_22_8_2),
		.out_wire_3_3(vertical_tile_23_8_to_tile_22_8_3),
		.in_wire_3_0(vertical_tile_22_8_to_tile_23_8_0),
		.in_wire_3_1(vertical_tile_22_8_to_tile_23_8_1),
		.in_wire_3_2(vertical_tile_22_8_to_tile_23_8_2),
		.in_wire_3_3(vertical_tile_22_8_to_tile_23_8_3),
		.out_wire_1_0(vertical_tile_23_8_to_tile_24_8_0),
		.out_wire_1_1(vertical_tile_23_8_to_tile_24_8_1),
		.out_wire_1_2(vertical_tile_23_8_to_tile_24_8_2),
		.out_wire_1_3(vertical_tile_23_8_to_tile_24_8_3),
		.in_wire_1_0(vertical_tile_24_8_to_tile_23_8_0),
		.in_wire_1_1(vertical_tile_24_8_to_tile_23_8_1),
		.in_wire_1_2(vertical_tile_24_8_to_tile_23_8_2),
		.in_wire_1_3(vertical_tile_24_8_to_tile_23_8_3),
		.out_wire_2_0(horizontal_tile_23_8_to_tile_23_7_0),
		.out_wire_2_1(horizontal_tile_23_8_to_tile_23_7_1),
		.out_wire_2_2(horizontal_tile_23_8_to_tile_23_7_2),
		.out_wire_2_3(horizontal_tile_23_8_to_tile_23_7_3),
		.in_wire_2_0(horizontal_tile_23_7_to_tile_23_8_0),
		.in_wire_2_1(horizontal_tile_23_7_to_tile_23_8_1),
		.in_wire_2_2(horizontal_tile_23_7_to_tile_23_8_2),
		.in_wire_2_3(horizontal_tile_23_7_to_tile_23_8_3),
		.out_wire_0_0(horizontal_tile_23_8_to_tile_23_9_0),
		.out_wire_0_1(horizontal_tile_23_8_to_tile_23_9_1),
		.out_wire_0_2(horizontal_tile_23_8_to_tile_23_9_2),
		.out_wire_0_3(horizontal_tile_23_8_to_tile_23_9_3),
		.in_wire_0_0(horizontal_tile_23_9_to_tile_23_8_0),
		.in_wire_0_1(horizontal_tile_23_9_to_tile_23_8_1),
		.in_wire_0_2(horizontal_tile_23_9_to_tile_23_8_2),
		.in_wire_0_3(horizontal_tile_23_9_to_tile_23_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(745)
	);

	pe_tile pe_tile_23_9(
		.out_wire_3_0(vertical_tile_23_9_to_tile_22_9_0),
		.out_wire_3_1(vertical_tile_23_9_to_tile_22_9_1),
		.out_wire_3_2(vertical_tile_23_9_to_tile_22_9_2),
		.out_wire_3_3(vertical_tile_23_9_to_tile_22_9_3),
		.in_wire_3_0(vertical_tile_22_9_to_tile_23_9_0),
		.in_wire_3_1(vertical_tile_22_9_to_tile_23_9_1),
		.in_wire_3_2(vertical_tile_22_9_to_tile_23_9_2),
		.in_wire_3_3(vertical_tile_22_9_to_tile_23_9_3),
		.out_wire_1_0(vertical_tile_23_9_to_tile_24_9_0),
		.out_wire_1_1(vertical_tile_23_9_to_tile_24_9_1),
		.out_wire_1_2(vertical_tile_23_9_to_tile_24_9_2),
		.out_wire_1_3(vertical_tile_23_9_to_tile_24_9_3),
		.in_wire_1_0(vertical_tile_24_9_to_tile_23_9_0),
		.in_wire_1_1(vertical_tile_24_9_to_tile_23_9_1),
		.in_wire_1_2(vertical_tile_24_9_to_tile_23_9_2),
		.in_wire_1_3(vertical_tile_24_9_to_tile_23_9_3),
		.out_wire_2_0(horizontal_tile_23_9_to_tile_23_8_0),
		.out_wire_2_1(horizontal_tile_23_9_to_tile_23_8_1),
		.out_wire_2_2(horizontal_tile_23_9_to_tile_23_8_2),
		.out_wire_2_3(horizontal_tile_23_9_to_tile_23_8_3),
		.in_wire_2_0(horizontal_tile_23_8_to_tile_23_9_0),
		.in_wire_2_1(horizontal_tile_23_8_to_tile_23_9_1),
		.in_wire_2_2(horizontal_tile_23_8_to_tile_23_9_2),
		.in_wire_2_3(horizontal_tile_23_8_to_tile_23_9_3),
		.out_wire_0_0(horizontal_tile_23_9_to_tile_23_10_0),
		.out_wire_0_1(horizontal_tile_23_9_to_tile_23_10_1),
		.out_wire_0_2(horizontal_tile_23_9_to_tile_23_10_2),
		.out_wire_0_3(horizontal_tile_23_9_to_tile_23_10_3),
		.in_wire_0_0(horizontal_tile_23_10_to_tile_23_9_0),
		.in_wire_0_1(horizontal_tile_23_10_to_tile_23_9_1),
		.in_wire_0_2(horizontal_tile_23_10_to_tile_23_9_2),
		.in_wire_0_3(horizontal_tile_23_10_to_tile_23_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(746)
	);

	pe_tile pe_tile_23_10(
		.out_wire_3_0(vertical_tile_23_10_to_tile_22_10_0),
		.out_wire_3_1(vertical_tile_23_10_to_tile_22_10_1),
		.out_wire_3_2(vertical_tile_23_10_to_tile_22_10_2),
		.out_wire_3_3(vertical_tile_23_10_to_tile_22_10_3),
		.in_wire_3_0(vertical_tile_22_10_to_tile_23_10_0),
		.in_wire_3_1(vertical_tile_22_10_to_tile_23_10_1),
		.in_wire_3_2(vertical_tile_22_10_to_tile_23_10_2),
		.in_wire_3_3(vertical_tile_22_10_to_tile_23_10_3),
		.out_wire_1_0(vertical_tile_23_10_to_tile_24_10_0),
		.out_wire_1_1(vertical_tile_23_10_to_tile_24_10_1),
		.out_wire_1_2(vertical_tile_23_10_to_tile_24_10_2),
		.out_wire_1_3(vertical_tile_23_10_to_tile_24_10_3),
		.in_wire_1_0(vertical_tile_24_10_to_tile_23_10_0),
		.in_wire_1_1(vertical_tile_24_10_to_tile_23_10_1),
		.in_wire_1_2(vertical_tile_24_10_to_tile_23_10_2),
		.in_wire_1_3(vertical_tile_24_10_to_tile_23_10_3),
		.out_wire_2_0(horizontal_tile_23_10_to_tile_23_9_0),
		.out_wire_2_1(horizontal_tile_23_10_to_tile_23_9_1),
		.out_wire_2_2(horizontal_tile_23_10_to_tile_23_9_2),
		.out_wire_2_3(horizontal_tile_23_10_to_tile_23_9_3),
		.in_wire_2_0(horizontal_tile_23_9_to_tile_23_10_0),
		.in_wire_2_1(horizontal_tile_23_9_to_tile_23_10_1),
		.in_wire_2_2(horizontal_tile_23_9_to_tile_23_10_2),
		.in_wire_2_3(horizontal_tile_23_9_to_tile_23_10_3),
		.out_wire_0_0(horizontal_tile_23_10_to_tile_23_11_0),
		.out_wire_0_1(horizontal_tile_23_10_to_tile_23_11_1),
		.out_wire_0_2(horizontal_tile_23_10_to_tile_23_11_2),
		.out_wire_0_3(horizontal_tile_23_10_to_tile_23_11_3),
		.in_wire_0_0(horizontal_tile_23_11_to_tile_23_10_0),
		.in_wire_0_1(horizontal_tile_23_11_to_tile_23_10_1),
		.in_wire_0_2(horizontal_tile_23_11_to_tile_23_10_2),
		.in_wire_0_3(horizontal_tile_23_11_to_tile_23_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(747)
	);

	pe_tile pe_tile_23_11(
		.out_wire_3_0(vertical_tile_23_11_to_tile_22_11_0),
		.out_wire_3_1(vertical_tile_23_11_to_tile_22_11_1),
		.out_wire_3_2(vertical_tile_23_11_to_tile_22_11_2),
		.out_wire_3_3(vertical_tile_23_11_to_tile_22_11_3),
		.in_wire_3_0(vertical_tile_22_11_to_tile_23_11_0),
		.in_wire_3_1(vertical_tile_22_11_to_tile_23_11_1),
		.in_wire_3_2(vertical_tile_22_11_to_tile_23_11_2),
		.in_wire_3_3(vertical_tile_22_11_to_tile_23_11_3),
		.out_wire_1_0(vertical_tile_23_11_to_tile_24_11_0),
		.out_wire_1_1(vertical_tile_23_11_to_tile_24_11_1),
		.out_wire_1_2(vertical_tile_23_11_to_tile_24_11_2),
		.out_wire_1_3(vertical_tile_23_11_to_tile_24_11_3),
		.in_wire_1_0(vertical_tile_24_11_to_tile_23_11_0),
		.in_wire_1_1(vertical_tile_24_11_to_tile_23_11_1),
		.in_wire_1_2(vertical_tile_24_11_to_tile_23_11_2),
		.in_wire_1_3(vertical_tile_24_11_to_tile_23_11_3),
		.out_wire_2_0(horizontal_tile_23_11_to_tile_23_10_0),
		.out_wire_2_1(horizontal_tile_23_11_to_tile_23_10_1),
		.out_wire_2_2(horizontal_tile_23_11_to_tile_23_10_2),
		.out_wire_2_3(horizontal_tile_23_11_to_tile_23_10_3),
		.in_wire_2_0(horizontal_tile_23_10_to_tile_23_11_0),
		.in_wire_2_1(horizontal_tile_23_10_to_tile_23_11_1),
		.in_wire_2_2(horizontal_tile_23_10_to_tile_23_11_2),
		.in_wire_2_3(horizontal_tile_23_10_to_tile_23_11_3),
		.out_wire_0_0(horizontal_tile_23_11_to_tile_23_12_0),
		.out_wire_0_1(horizontal_tile_23_11_to_tile_23_12_1),
		.out_wire_0_2(horizontal_tile_23_11_to_tile_23_12_2),
		.out_wire_0_3(horizontal_tile_23_11_to_tile_23_12_3),
		.in_wire_0_0(horizontal_tile_23_12_to_tile_23_11_0),
		.in_wire_0_1(horizontal_tile_23_12_to_tile_23_11_1),
		.in_wire_0_2(horizontal_tile_23_12_to_tile_23_11_2),
		.in_wire_0_3(horizontal_tile_23_12_to_tile_23_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(748)
	);

	pe_tile pe_tile_23_12(
		.out_wire_3_0(vertical_tile_23_12_to_tile_22_12_0),
		.out_wire_3_1(vertical_tile_23_12_to_tile_22_12_1),
		.out_wire_3_2(vertical_tile_23_12_to_tile_22_12_2),
		.out_wire_3_3(vertical_tile_23_12_to_tile_22_12_3),
		.in_wire_3_0(vertical_tile_22_12_to_tile_23_12_0),
		.in_wire_3_1(vertical_tile_22_12_to_tile_23_12_1),
		.in_wire_3_2(vertical_tile_22_12_to_tile_23_12_2),
		.in_wire_3_3(vertical_tile_22_12_to_tile_23_12_3),
		.out_wire_1_0(vertical_tile_23_12_to_tile_24_12_0),
		.out_wire_1_1(vertical_tile_23_12_to_tile_24_12_1),
		.out_wire_1_2(vertical_tile_23_12_to_tile_24_12_2),
		.out_wire_1_3(vertical_tile_23_12_to_tile_24_12_3),
		.in_wire_1_0(vertical_tile_24_12_to_tile_23_12_0),
		.in_wire_1_1(vertical_tile_24_12_to_tile_23_12_1),
		.in_wire_1_2(vertical_tile_24_12_to_tile_23_12_2),
		.in_wire_1_3(vertical_tile_24_12_to_tile_23_12_3),
		.out_wire_2_0(horizontal_tile_23_12_to_tile_23_11_0),
		.out_wire_2_1(horizontal_tile_23_12_to_tile_23_11_1),
		.out_wire_2_2(horizontal_tile_23_12_to_tile_23_11_2),
		.out_wire_2_3(horizontal_tile_23_12_to_tile_23_11_3),
		.in_wire_2_0(horizontal_tile_23_11_to_tile_23_12_0),
		.in_wire_2_1(horizontal_tile_23_11_to_tile_23_12_1),
		.in_wire_2_2(horizontal_tile_23_11_to_tile_23_12_2),
		.in_wire_2_3(horizontal_tile_23_11_to_tile_23_12_3),
		.out_wire_0_0(horizontal_tile_23_12_to_tile_23_13_0),
		.out_wire_0_1(horizontal_tile_23_12_to_tile_23_13_1),
		.out_wire_0_2(horizontal_tile_23_12_to_tile_23_13_2),
		.out_wire_0_3(horizontal_tile_23_12_to_tile_23_13_3),
		.in_wire_0_0(horizontal_tile_23_13_to_tile_23_12_0),
		.in_wire_0_1(horizontal_tile_23_13_to_tile_23_12_1),
		.in_wire_0_2(horizontal_tile_23_13_to_tile_23_12_2),
		.in_wire_0_3(horizontal_tile_23_13_to_tile_23_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(749)
	);

	pe_tile pe_tile_23_13(
		.out_wire_3_0(vertical_tile_23_13_to_tile_22_13_0),
		.out_wire_3_1(vertical_tile_23_13_to_tile_22_13_1),
		.out_wire_3_2(vertical_tile_23_13_to_tile_22_13_2),
		.out_wire_3_3(vertical_tile_23_13_to_tile_22_13_3),
		.in_wire_3_0(vertical_tile_22_13_to_tile_23_13_0),
		.in_wire_3_1(vertical_tile_22_13_to_tile_23_13_1),
		.in_wire_3_2(vertical_tile_22_13_to_tile_23_13_2),
		.in_wire_3_3(vertical_tile_22_13_to_tile_23_13_3),
		.out_wire_1_0(vertical_tile_23_13_to_tile_24_13_0),
		.out_wire_1_1(vertical_tile_23_13_to_tile_24_13_1),
		.out_wire_1_2(vertical_tile_23_13_to_tile_24_13_2),
		.out_wire_1_3(vertical_tile_23_13_to_tile_24_13_3),
		.in_wire_1_0(vertical_tile_24_13_to_tile_23_13_0),
		.in_wire_1_1(vertical_tile_24_13_to_tile_23_13_1),
		.in_wire_1_2(vertical_tile_24_13_to_tile_23_13_2),
		.in_wire_1_3(vertical_tile_24_13_to_tile_23_13_3),
		.out_wire_2_0(horizontal_tile_23_13_to_tile_23_12_0),
		.out_wire_2_1(horizontal_tile_23_13_to_tile_23_12_1),
		.out_wire_2_2(horizontal_tile_23_13_to_tile_23_12_2),
		.out_wire_2_3(horizontal_tile_23_13_to_tile_23_12_3),
		.in_wire_2_0(horizontal_tile_23_12_to_tile_23_13_0),
		.in_wire_2_1(horizontal_tile_23_12_to_tile_23_13_1),
		.in_wire_2_2(horizontal_tile_23_12_to_tile_23_13_2),
		.in_wire_2_3(horizontal_tile_23_12_to_tile_23_13_3),
		.out_wire_0_0(horizontal_tile_23_13_to_tile_23_14_0),
		.out_wire_0_1(horizontal_tile_23_13_to_tile_23_14_1),
		.out_wire_0_2(horizontal_tile_23_13_to_tile_23_14_2),
		.out_wire_0_3(horizontal_tile_23_13_to_tile_23_14_3),
		.in_wire_0_0(horizontal_tile_23_14_to_tile_23_13_0),
		.in_wire_0_1(horizontal_tile_23_14_to_tile_23_13_1),
		.in_wire_0_2(horizontal_tile_23_14_to_tile_23_13_2),
		.in_wire_0_3(horizontal_tile_23_14_to_tile_23_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(750)
	);

	pe_tile pe_tile_23_14(
		.out_wire_3_0(vertical_tile_23_14_to_tile_22_14_0),
		.out_wire_3_1(vertical_tile_23_14_to_tile_22_14_1),
		.out_wire_3_2(vertical_tile_23_14_to_tile_22_14_2),
		.out_wire_3_3(vertical_tile_23_14_to_tile_22_14_3),
		.in_wire_3_0(vertical_tile_22_14_to_tile_23_14_0),
		.in_wire_3_1(vertical_tile_22_14_to_tile_23_14_1),
		.in_wire_3_2(vertical_tile_22_14_to_tile_23_14_2),
		.in_wire_3_3(vertical_tile_22_14_to_tile_23_14_3),
		.out_wire_1_0(vertical_tile_23_14_to_tile_24_14_0),
		.out_wire_1_1(vertical_tile_23_14_to_tile_24_14_1),
		.out_wire_1_2(vertical_tile_23_14_to_tile_24_14_2),
		.out_wire_1_3(vertical_tile_23_14_to_tile_24_14_3),
		.in_wire_1_0(vertical_tile_24_14_to_tile_23_14_0),
		.in_wire_1_1(vertical_tile_24_14_to_tile_23_14_1),
		.in_wire_1_2(vertical_tile_24_14_to_tile_23_14_2),
		.in_wire_1_3(vertical_tile_24_14_to_tile_23_14_3),
		.out_wire_2_0(horizontal_tile_23_14_to_tile_23_13_0),
		.out_wire_2_1(horizontal_tile_23_14_to_tile_23_13_1),
		.out_wire_2_2(horizontal_tile_23_14_to_tile_23_13_2),
		.out_wire_2_3(horizontal_tile_23_14_to_tile_23_13_3),
		.in_wire_2_0(horizontal_tile_23_13_to_tile_23_14_0),
		.in_wire_2_1(horizontal_tile_23_13_to_tile_23_14_1),
		.in_wire_2_2(horizontal_tile_23_13_to_tile_23_14_2),
		.in_wire_2_3(horizontal_tile_23_13_to_tile_23_14_3),
		.out_wire_0_0(horizontal_tile_23_14_to_tile_23_15_0),
		.out_wire_0_1(horizontal_tile_23_14_to_tile_23_15_1),
		.out_wire_0_2(horizontal_tile_23_14_to_tile_23_15_2),
		.out_wire_0_3(horizontal_tile_23_14_to_tile_23_15_3),
		.in_wire_0_0(horizontal_tile_23_15_to_tile_23_14_0),
		.in_wire_0_1(horizontal_tile_23_15_to_tile_23_14_1),
		.in_wire_0_2(horizontal_tile_23_15_to_tile_23_14_2),
		.in_wire_0_3(horizontal_tile_23_15_to_tile_23_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(751)
	);

	pe_tile pe_tile_23_15(
		.out_wire_3_0(vertical_tile_23_15_to_tile_22_15_0),
		.out_wire_3_1(vertical_tile_23_15_to_tile_22_15_1),
		.out_wire_3_2(vertical_tile_23_15_to_tile_22_15_2),
		.out_wire_3_3(vertical_tile_23_15_to_tile_22_15_3),
		.in_wire_3_0(vertical_tile_22_15_to_tile_23_15_0),
		.in_wire_3_1(vertical_tile_22_15_to_tile_23_15_1),
		.in_wire_3_2(vertical_tile_22_15_to_tile_23_15_2),
		.in_wire_3_3(vertical_tile_22_15_to_tile_23_15_3),
		.out_wire_1_0(vertical_tile_23_15_to_tile_24_15_0),
		.out_wire_1_1(vertical_tile_23_15_to_tile_24_15_1),
		.out_wire_1_2(vertical_tile_23_15_to_tile_24_15_2),
		.out_wire_1_3(vertical_tile_23_15_to_tile_24_15_3),
		.in_wire_1_0(vertical_tile_24_15_to_tile_23_15_0),
		.in_wire_1_1(vertical_tile_24_15_to_tile_23_15_1),
		.in_wire_1_2(vertical_tile_24_15_to_tile_23_15_2),
		.in_wire_1_3(vertical_tile_24_15_to_tile_23_15_3),
		.out_wire_2_0(horizontal_tile_23_15_to_tile_23_14_0),
		.out_wire_2_1(horizontal_tile_23_15_to_tile_23_14_1),
		.out_wire_2_2(horizontal_tile_23_15_to_tile_23_14_2),
		.out_wire_2_3(horizontal_tile_23_15_to_tile_23_14_3),
		.in_wire_2_0(horizontal_tile_23_14_to_tile_23_15_0),
		.in_wire_2_1(horizontal_tile_23_14_to_tile_23_15_1),
		.in_wire_2_2(horizontal_tile_23_14_to_tile_23_15_2),
		.in_wire_2_3(horizontal_tile_23_14_to_tile_23_15_3),
		.out_wire_0_0(horizontal_tile_23_15_to_tile_23_16_0),
		.out_wire_0_1(horizontal_tile_23_15_to_tile_23_16_1),
		.out_wire_0_2(horizontal_tile_23_15_to_tile_23_16_2),
		.out_wire_0_3(horizontal_tile_23_15_to_tile_23_16_3),
		.in_wire_0_0(horizontal_tile_23_16_to_tile_23_15_0),
		.in_wire_0_1(horizontal_tile_23_16_to_tile_23_15_1),
		.in_wire_0_2(horizontal_tile_23_16_to_tile_23_15_2),
		.in_wire_0_3(horizontal_tile_23_16_to_tile_23_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(752)
	);

	pe_tile pe_tile_23_16(
		.out_wire_3_0(vertical_tile_23_16_to_tile_22_16_0),
		.out_wire_3_1(vertical_tile_23_16_to_tile_22_16_1),
		.out_wire_3_2(vertical_tile_23_16_to_tile_22_16_2),
		.out_wire_3_3(vertical_tile_23_16_to_tile_22_16_3),
		.in_wire_3_0(vertical_tile_22_16_to_tile_23_16_0),
		.in_wire_3_1(vertical_tile_22_16_to_tile_23_16_1),
		.in_wire_3_2(vertical_tile_22_16_to_tile_23_16_2),
		.in_wire_3_3(vertical_tile_22_16_to_tile_23_16_3),
		.out_wire_1_0(vertical_tile_23_16_to_tile_24_16_0),
		.out_wire_1_1(vertical_tile_23_16_to_tile_24_16_1),
		.out_wire_1_2(vertical_tile_23_16_to_tile_24_16_2),
		.out_wire_1_3(vertical_tile_23_16_to_tile_24_16_3),
		.in_wire_1_0(vertical_tile_24_16_to_tile_23_16_0),
		.in_wire_1_1(vertical_tile_24_16_to_tile_23_16_1),
		.in_wire_1_2(vertical_tile_24_16_to_tile_23_16_2),
		.in_wire_1_3(vertical_tile_24_16_to_tile_23_16_3),
		.out_wire_2_0(horizontal_tile_23_16_to_tile_23_15_0),
		.out_wire_2_1(horizontal_tile_23_16_to_tile_23_15_1),
		.out_wire_2_2(horizontal_tile_23_16_to_tile_23_15_2),
		.out_wire_2_3(horizontal_tile_23_16_to_tile_23_15_3),
		.in_wire_2_0(horizontal_tile_23_15_to_tile_23_16_0),
		.in_wire_2_1(horizontal_tile_23_15_to_tile_23_16_1),
		.in_wire_2_2(horizontal_tile_23_15_to_tile_23_16_2),
		.in_wire_2_3(horizontal_tile_23_15_to_tile_23_16_3),
		.out_wire_0_0(horizontal_tile_23_16_to_tile_23_17_0),
		.out_wire_0_1(horizontal_tile_23_16_to_tile_23_17_1),
		.out_wire_0_2(horizontal_tile_23_16_to_tile_23_17_2),
		.out_wire_0_3(horizontal_tile_23_16_to_tile_23_17_3),
		.in_wire_0_0(horizontal_tile_23_17_to_tile_23_16_0),
		.in_wire_0_1(horizontal_tile_23_17_to_tile_23_16_1),
		.in_wire_0_2(horizontal_tile_23_17_to_tile_23_16_2),
		.in_wire_0_3(horizontal_tile_23_17_to_tile_23_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(753)
	);

	pe_tile pe_tile_23_17(
		.out_wire_3_0(vertical_tile_23_17_to_tile_22_17_0),
		.out_wire_3_1(vertical_tile_23_17_to_tile_22_17_1),
		.out_wire_3_2(vertical_tile_23_17_to_tile_22_17_2),
		.out_wire_3_3(vertical_tile_23_17_to_tile_22_17_3),
		.in_wire_3_0(vertical_tile_22_17_to_tile_23_17_0),
		.in_wire_3_1(vertical_tile_22_17_to_tile_23_17_1),
		.in_wire_3_2(vertical_tile_22_17_to_tile_23_17_2),
		.in_wire_3_3(vertical_tile_22_17_to_tile_23_17_3),
		.out_wire_1_0(vertical_tile_23_17_to_tile_24_17_0),
		.out_wire_1_1(vertical_tile_23_17_to_tile_24_17_1),
		.out_wire_1_2(vertical_tile_23_17_to_tile_24_17_2),
		.out_wire_1_3(vertical_tile_23_17_to_tile_24_17_3),
		.in_wire_1_0(vertical_tile_24_17_to_tile_23_17_0),
		.in_wire_1_1(vertical_tile_24_17_to_tile_23_17_1),
		.in_wire_1_2(vertical_tile_24_17_to_tile_23_17_2),
		.in_wire_1_3(vertical_tile_24_17_to_tile_23_17_3),
		.out_wire_2_0(horizontal_tile_23_17_to_tile_23_16_0),
		.out_wire_2_1(horizontal_tile_23_17_to_tile_23_16_1),
		.out_wire_2_2(horizontal_tile_23_17_to_tile_23_16_2),
		.out_wire_2_3(horizontal_tile_23_17_to_tile_23_16_3),
		.in_wire_2_0(horizontal_tile_23_16_to_tile_23_17_0),
		.in_wire_2_1(horizontal_tile_23_16_to_tile_23_17_1),
		.in_wire_2_2(horizontal_tile_23_16_to_tile_23_17_2),
		.in_wire_2_3(horizontal_tile_23_16_to_tile_23_17_3),
		.out_wire_0_0(horizontal_tile_23_17_to_tile_23_18_0),
		.out_wire_0_1(horizontal_tile_23_17_to_tile_23_18_1),
		.out_wire_0_2(horizontal_tile_23_17_to_tile_23_18_2),
		.out_wire_0_3(horizontal_tile_23_17_to_tile_23_18_3),
		.in_wire_0_0(horizontal_tile_23_18_to_tile_23_17_0),
		.in_wire_0_1(horizontal_tile_23_18_to_tile_23_17_1),
		.in_wire_0_2(horizontal_tile_23_18_to_tile_23_17_2),
		.in_wire_0_3(horizontal_tile_23_18_to_tile_23_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(754)
	);

	pe_tile pe_tile_23_18(
		.out_wire_3_0(vertical_tile_23_18_to_tile_22_18_0),
		.out_wire_3_1(vertical_tile_23_18_to_tile_22_18_1),
		.out_wire_3_2(vertical_tile_23_18_to_tile_22_18_2),
		.out_wire_3_3(vertical_tile_23_18_to_tile_22_18_3),
		.in_wire_3_0(vertical_tile_22_18_to_tile_23_18_0),
		.in_wire_3_1(vertical_tile_22_18_to_tile_23_18_1),
		.in_wire_3_2(vertical_tile_22_18_to_tile_23_18_2),
		.in_wire_3_3(vertical_tile_22_18_to_tile_23_18_3),
		.out_wire_1_0(vertical_tile_23_18_to_tile_24_18_0),
		.out_wire_1_1(vertical_tile_23_18_to_tile_24_18_1),
		.out_wire_1_2(vertical_tile_23_18_to_tile_24_18_2),
		.out_wire_1_3(vertical_tile_23_18_to_tile_24_18_3),
		.in_wire_1_0(vertical_tile_24_18_to_tile_23_18_0),
		.in_wire_1_1(vertical_tile_24_18_to_tile_23_18_1),
		.in_wire_1_2(vertical_tile_24_18_to_tile_23_18_2),
		.in_wire_1_3(vertical_tile_24_18_to_tile_23_18_3),
		.out_wire_2_0(horizontal_tile_23_18_to_tile_23_17_0),
		.out_wire_2_1(horizontal_tile_23_18_to_tile_23_17_1),
		.out_wire_2_2(horizontal_tile_23_18_to_tile_23_17_2),
		.out_wire_2_3(horizontal_tile_23_18_to_tile_23_17_3),
		.in_wire_2_0(horizontal_tile_23_17_to_tile_23_18_0),
		.in_wire_2_1(horizontal_tile_23_17_to_tile_23_18_1),
		.in_wire_2_2(horizontal_tile_23_17_to_tile_23_18_2),
		.in_wire_2_3(horizontal_tile_23_17_to_tile_23_18_3),
		.out_wire_0_0(horizontal_tile_23_18_to_tile_23_19_0),
		.out_wire_0_1(horizontal_tile_23_18_to_tile_23_19_1),
		.out_wire_0_2(horizontal_tile_23_18_to_tile_23_19_2),
		.out_wire_0_3(horizontal_tile_23_18_to_tile_23_19_3),
		.in_wire_0_0(horizontal_tile_23_19_to_tile_23_18_0),
		.in_wire_0_1(horizontal_tile_23_19_to_tile_23_18_1),
		.in_wire_0_2(horizontal_tile_23_19_to_tile_23_18_2),
		.in_wire_0_3(horizontal_tile_23_19_to_tile_23_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(755)
	);

	pe_tile pe_tile_23_19(
		.out_wire_3_0(vertical_tile_23_19_to_tile_22_19_0),
		.out_wire_3_1(vertical_tile_23_19_to_tile_22_19_1),
		.out_wire_3_2(vertical_tile_23_19_to_tile_22_19_2),
		.out_wire_3_3(vertical_tile_23_19_to_tile_22_19_3),
		.in_wire_3_0(vertical_tile_22_19_to_tile_23_19_0),
		.in_wire_3_1(vertical_tile_22_19_to_tile_23_19_1),
		.in_wire_3_2(vertical_tile_22_19_to_tile_23_19_2),
		.in_wire_3_3(vertical_tile_22_19_to_tile_23_19_3),
		.out_wire_1_0(vertical_tile_23_19_to_tile_24_19_0),
		.out_wire_1_1(vertical_tile_23_19_to_tile_24_19_1),
		.out_wire_1_2(vertical_tile_23_19_to_tile_24_19_2),
		.out_wire_1_3(vertical_tile_23_19_to_tile_24_19_3),
		.in_wire_1_0(vertical_tile_24_19_to_tile_23_19_0),
		.in_wire_1_1(vertical_tile_24_19_to_tile_23_19_1),
		.in_wire_1_2(vertical_tile_24_19_to_tile_23_19_2),
		.in_wire_1_3(vertical_tile_24_19_to_tile_23_19_3),
		.out_wire_2_0(horizontal_tile_23_19_to_tile_23_18_0),
		.out_wire_2_1(horizontal_tile_23_19_to_tile_23_18_1),
		.out_wire_2_2(horizontal_tile_23_19_to_tile_23_18_2),
		.out_wire_2_3(horizontal_tile_23_19_to_tile_23_18_3),
		.in_wire_2_0(horizontal_tile_23_18_to_tile_23_19_0),
		.in_wire_2_1(horizontal_tile_23_18_to_tile_23_19_1),
		.in_wire_2_2(horizontal_tile_23_18_to_tile_23_19_2),
		.in_wire_2_3(horizontal_tile_23_18_to_tile_23_19_3),
		.out_wire_0_0(horizontal_tile_23_19_to_tile_23_20_0),
		.out_wire_0_1(horizontal_tile_23_19_to_tile_23_20_1),
		.out_wire_0_2(horizontal_tile_23_19_to_tile_23_20_2),
		.out_wire_0_3(horizontal_tile_23_19_to_tile_23_20_3),
		.in_wire_0_0(horizontal_tile_23_20_to_tile_23_19_0),
		.in_wire_0_1(horizontal_tile_23_20_to_tile_23_19_1),
		.in_wire_0_2(horizontal_tile_23_20_to_tile_23_19_2),
		.in_wire_0_3(horizontal_tile_23_20_to_tile_23_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(756)
	);

	pe_tile pe_tile_23_20(
		.out_wire_3_0(vertical_tile_23_20_to_tile_22_20_0),
		.out_wire_3_1(vertical_tile_23_20_to_tile_22_20_1),
		.out_wire_3_2(vertical_tile_23_20_to_tile_22_20_2),
		.out_wire_3_3(vertical_tile_23_20_to_tile_22_20_3),
		.in_wire_3_0(vertical_tile_22_20_to_tile_23_20_0),
		.in_wire_3_1(vertical_tile_22_20_to_tile_23_20_1),
		.in_wire_3_2(vertical_tile_22_20_to_tile_23_20_2),
		.in_wire_3_3(vertical_tile_22_20_to_tile_23_20_3),
		.out_wire_1_0(vertical_tile_23_20_to_tile_24_20_0),
		.out_wire_1_1(vertical_tile_23_20_to_tile_24_20_1),
		.out_wire_1_2(vertical_tile_23_20_to_tile_24_20_2),
		.out_wire_1_3(vertical_tile_23_20_to_tile_24_20_3),
		.in_wire_1_0(vertical_tile_24_20_to_tile_23_20_0),
		.in_wire_1_1(vertical_tile_24_20_to_tile_23_20_1),
		.in_wire_1_2(vertical_tile_24_20_to_tile_23_20_2),
		.in_wire_1_3(vertical_tile_24_20_to_tile_23_20_3),
		.out_wire_2_0(horizontal_tile_23_20_to_tile_23_19_0),
		.out_wire_2_1(horizontal_tile_23_20_to_tile_23_19_1),
		.out_wire_2_2(horizontal_tile_23_20_to_tile_23_19_2),
		.out_wire_2_3(horizontal_tile_23_20_to_tile_23_19_3),
		.in_wire_2_0(horizontal_tile_23_19_to_tile_23_20_0),
		.in_wire_2_1(horizontal_tile_23_19_to_tile_23_20_1),
		.in_wire_2_2(horizontal_tile_23_19_to_tile_23_20_2),
		.in_wire_2_3(horizontal_tile_23_19_to_tile_23_20_3),
		.out_wire_0_0(horizontal_tile_23_20_to_tile_23_21_0),
		.out_wire_0_1(horizontal_tile_23_20_to_tile_23_21_1),
		.out_wire_0_2(horizontal_tile_23_20_to_tile_23_21_2),
		.out_wire_0_3(horizontal_tile_23_20_to_tile_23_21_3),
		.in_wire_0_0(horizontal_tile_23_21_to_tile_23_20_0),
		.in_wire_0_1(horizontal_tile_23_21_to_tile_23_20_1),
		.in_wire_0_2(horizontal_tile_23_21_to_tile_23_20_2),
		.in_wire_0_3(horizontal_tile_23_21_to_tile_23_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(757)
	);

	pe_tile pe_tile_23_21(
		.out_wire_3_0(vertical_tile_23_21_to_tile_22_21_0),
		.out_wire_3_1(vertical_tile_23_21_to_tile_22_21_1),
		.out_wire_3_2(vertical_tile_23_21_to_tile_22_21_2),
		.out_wire_3_3(vertical_tile_23_21_to_tile_22_21_3),
		.in_wire_3_0(vertical_tile_22_21_to_tile_23_21_0),
		.in_wire_3_1(vertical_tile_22_21_to_tile_23_21_1),
		.in_wire_3_2(vertical_tile_22_21_to_tile_23_21_2),
		.in_wire_3_3(vertical_tile_22_21_to_tile_23_21_3),
		.out_wire_1_0(vertical_tile_23_21_to_tile_24_21_0),
		.out_wire_1_1(vertical_tile_23_21_to_tile_24_21_1),
		.out_wire_1_2(vertical_tile_23_21_to_tile_24_21_2),
		.out_wire_1_3(vertical_tile_23_21_to_tile_24_21_3),
		.in_wire_1_0(vertical_tile_24_21_to_tile_23_21_0),
		.in_wire_1_1(vertical_tile_24_21_to_tile_23_21_1),
		.in_wire_1_2(vertical_tile_24_21_to_tile_23_21_2),
		.in_wire_1_3(vertical_tile_24_21_to_tile_23_21_3),
		.out_wire_2_0(horizontal_tile_23_21_to_tile_23_20_0),
		.out_wire_2_1(horizontal_tile_23_21_to_tile_23_20_1),
		.out_wire_2_2(horizontal_tile_23_21_to_tile_23_20_2),
		.out_wire_2_3(horizontal_tile_23_21_to_tile_23_20_3),
		.in_wire_2_0(horizontal_tile_23_20_to_tile_23_21_0),
		.in_wire_2_1(horizontal_tile_23_20_to_tile_23_21_1),
		.in_wire_2_2(horizontal_tile_23_20_to_tile_23_21_2),
		.in_wire_2_3(horizontal_tile_23_20_to_tile_23_21_3),
		.out_wire_0_0(horizontal_tile_23_21_to_tile_23_22_0),
		.out_wire_0_1(horizontal_tile_23_21_to_tile_23_22_1),
		.out_wire_0_2(horizontal_tile_23_21_to_tile_23_22_2),
		.out_wire_0_3(horizontal_tile_23_21_to_tile_23_22_3),
		.in_wire_0_0(horizontal_tile_23_22_to_tile_23_21_0),
		.in_wire_0_1(horizontal_tile_23_22_to_tile_23_21_1),
		.in_wire_0_2(horizontal_tile_23_22_to_tile_23_21_2),
		.in_wire_0_3(horizontal_tile_23_22_to_tile_23_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(758)
	);

	pe_tile pe_tile_23_22(
		.out_wire_3_0(vertical_tile_23_22_to_tile_22_22_0),
		.out_wire_3_1(vertical_tile_23_22_to_tile_22_22_1),
		.out_wire_3_2(vertical_tile_23_22_to_tile_22_22_2),
		.out_wire_3_3(vertical_tile_23_22_to_tile_22_22_3),
		.in_wire_3_0(vertical_tile_22_22_to_tile_23_22_0),
		.in_wire_3_1(vertical_tile_22_22_to_tile_23_22_1),
		.in_wire_3_2(vertical_tile_22_22_to_tile_23_22_2),
		.in_wire_3_3(vertical_tile_22_22_to_tile_23_22_3),
		.out_wire_1_0(vertical_tile_23_22_to_tile_24_22_0),
		.out_wire_1_1(vertical_tile_23_22_to_tile_24_22_1),
		.out_wire_1_2(vertical_tile_23_22_to_tile_24_22_2),
		.out_wire_1_3(vertical_tile_23_22_to_tile_24_22_3),
		.in_wire_1_0(vertical_tile_24_22_to_tile_23_22_0),
		.in_wire_1_1(vertical_tile_24_22_to_tile_23_22_1),
		.in_wire_1_2(vertical_tile_24_22_to_tile_23_22_2),
		.in_wire_1_3(vertical_tile_24_22_to_tile_23_22_3),
		.out_wire_2_0(horizontal_tile_23_22_to_tile_23_21_0),
		.out_wire_2_1(horizontal_tile_23_22_to_tile_23_21_1),
		.out_wire_2_2(horizontal_tile_23_22_to_tile_23_21_2),
		.out_wire_2_3(horizontal_tile_23_22_to_tile_23_21_3),
		.in_wire_2_0(horizontal_tile_23_21_to_tile_23_22_0),
		.in_wire_2_1(horizontal_tile_23_21_to_tile_23_22_1),
		.in_wire_2_2(horizontal_tile_23_21_to_tile_23_22_2),
		.in_wire_2_3(horizontal_tile_23_21_to_tile_23_22_3),
		.out_wire_0_0(horizontal_tile_23_22_to_tile_23_23_0),
		.out_wire_0_1(horizontal_tile_23_22_to_tile_23_23_1),
		.out_wire_0_2(horizontal_tile_23_22_to_tile_23_23_2),
		.out_wire_0_3(horizontal_tile_23_22_to_tile_23_23_3),
		.in_wire_0_0(horizontal_tile_23_23_to_tile_23_22_0),
		.in_wire_0_1(horizontal_tile_23_23_to_tile_23_22_1),
		.in_wire_0_2(horizontal_tile_23_23_to_tile_23_22_2),
		.in_wire_0_3(horizontal_tile_23_23_to_tile_23_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(759)
	);

	pe_tile pe_tile_23_23(
		.out_wire_3_0(vertical_tile_23_23_to_tile_22_23_0),
		.out_wire_3_1(vertical_tile_23_23_to_tile_22_23_1),
		.out_wire_3_2(vertical_tile_23_23_to_tile_22_23_2),
		.out_wire_3_3(vertical_tile_23_23_to_tile_22_23_3),
		.in_wire_3_0(vertical_tile_22_23_to_tile_23_23_0),
		.in_wire_3_1(vertical_tile_22_23_to_tile_23_23_1),
		.in_wire_3_2(vertical_tile_22_23_to_tile_23_23_2),
		.in_wire_3_3(vertical_tile_22_23_to_tile_23_23_3),
		.out_wire_1_0(vertical_tile_23_23_to_tile_24_23_0),
		.out_wire_1_1(vertical_tile_23_23_to_tile_24_23_1),
		.out_wire_1_2(vertical_tile_23_23_to_tile_24_23_2),
		.out_wire_1_3(vertical_tile_23_23_to_tile_24_23_3),
		.in_wire_1_0(vertical_tile_24_23_to_tile_23_23_0),
		.in_wire_1_1(vertical_tile_24_23_to_tile_23_23_1),
		.in_wire_1_2(vertical_tile_24_23_to_tile_23_23_2),
		.in_wire_1_3(vertical_tile_24_23_to_tile_23_23_3),
		.out_wire_2_0(horizontal_tile_23_23_to_tile_23_22_0),
		.out_wire_2_1(horizontal_tile_23_23_to_tile_23_22_1),
		.out_wire_2_2(horizontal_tile_23_23_to_tile_23_22_2),
		.out_wire_2_3(horizontal_tile_23_23_to_tile_23_22_3),
		.in_wire_2_0(horizontal_tile_23_22_to_tile_23_23_0),
		.in_wire_2_1(horizontal_tile_23_22_to_tile_23_23_1),
		.in_wire_2_2(horizontal_tile_23_22_to_tile_23_23_2),
		.in_wire_2_3(horizontal_tile_23_22_to_tile_23_23_3),
		.out_wire_0_0(horizontal_tile_23_23_to_tile_23_24_0),
		.out_wire_0_1(horizontal_tile_23_23_to_tile_23_24_1),
		.out_wire_0_2(horizontal_tile_23_23_to_tile_23_24_2),
		.out_wire_0_3(horizontal_tile_23_23_to_tile_23_24_3),
		.in_wire_0_0(horizontal_tile_23_24_to_tile_23_23_0),
		.in_wire_0_1(horizontal_tile_23_24_to_tile_23_23_1),
		.in_wire_0_2(horizontal_tile_23_24_to_tile_23_23_2),
		.in_wire_0_3(horizontal_tile_23_24_to_tile_23_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(760)
	);

	pe_tile pe_tile_23_24(
		.out_wire_3_0(vertical_tile_23_24_to_tile_22_24_0),
		.out_wire_3_1(vertical_tile_23_24_to_tile_22_24_1),
		.out_wire_3_2(vertical_tile_23_24_to_tile_22_24_2),
		.out_wire_3_3(vertical_tile_23_24_to_tile_22_24_3),
		.in_wire_3_0(vertical_tile_22_24_to_tile_23_24_0),
		.in_wire_3_1(vertical_tile_22_24_to_tile_23_24_1),
		.in_wire_3_2(vertical_tile_22_24_to_tile_23_24_2),
		.in_wire_3_3(vertical_tile_22_24_to_tile_23_24_3),
		.out_wire_1_0(vertical_tile_23_24_to_tile_24_24_0),
		.out_wire_1_1(vertical_tile_23_24_to_tile_24_24_1),
		.out_wire_1_2(vertical_tile_23_24_to_tile_24_24_2),
		.out_wire_1_3(vertical_tile_23_24_to_tile_24_24_3),
		.in_wire_1_0(vertical_tile_24_24_to_tile_23_24_0),
		.in_wire_1_1(vertical_tile_24_24_to_tile_23_24_1),
		.in_wire_1_2(vertical_tile_24_24_to_tile_23_24_2),
		.in_wire_1_3(vertical_tile_24_24_to_tile_23_24_3),
		.out_wire_2_0(horizontal_tile_23_24_to_tile_23_23_0),
		.out_wire_2_1(horizontal_tile_23_24_to_tile_23_23_1),
		.out_wire_2_2(horizontal_tile_23_24_to_tile_23_23_2),
		.out_wire_2_3(horizontal_tile_23_24_to_tile_23_23_3),
		.in_wire_2_0(horizontal_tile_23_23_to_tile_23_24_0),
		.in_wire_2_1(horizontal_tile_23_23_to_tile_23_24_1),
		.in_wire_2_2(horizontal_tile_23_23_to_tile_23_24_2),
		.in_wire_2_3(horizontal_tile_23_23_to_tile_23_24_3),
		.out_wire_0_0(horizontal_tile_23_24_to_tile_23_25_0),
		.out_wire_0_1(horizontal_tile_23_24_to_tile_23_25_1),
		.out_wire_0_2(horizontal_tile_23_24_to_tile_23_25_2),
		.out_wire_0_3(horizontal_tile_23_24_to_tile_23_25_3),
		.in_wire_0_0(horizontal_tile_23_25_to_tile_23_24_0),
		.in_wire_0_1(horizontal_tile_23_25_to_tile_23_24_1),
		.in_wire_0_2(horizontal_tile_23_25_to_tile_23_24_2),
		.in_wire_0_3(horizontal_tile_23_25_to_tile_23_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(761)
	);

	pe_tile pe_tile_23_25(
		.out_wire_3_0(vertical_tile_23_25_to_tile_22_25_0),
		.out_wire_3_1(vertical_tile_23_25_to_tile_22_25_1),
		.out_wire_3_2(vertical_tile_23_25_to_tile_22_25_2),
		.out_wire_3_3(vertical_tile_23_25_to_tile_22_25_3),
		.in_wire_3_0(vertical_tile_22_25_to_tile_23_25_0),
		.in_wire_3_1(vertical_tile_22_25_to_tile_23_25_1),
		.in_wire_3_2(vertical_tile_22_25_to_tile_23_25_2),
		.in_wire_3_3(vertical_tile_22_25_to_tile_23_25_3),
		.out_wire_1_0(vertical_tile_23_25_to_tile_24_25_0),
		.out_wire_1_1(vertical_tile_23_25_to_tile_24_25_1),
		.out_wire_1_2(vertical_tile_23_25_to_tile_24_25_2),
		.out_wire_1_3(vertical_tile_23_25_to_tile_24_25_3),
		.in_wire_1_0(vertical_tile_24_25_to_tile_23_25_0),
		.in_wire_1_1(vertical_tile_24_25_to_tile_23_25_1),
		.in_wire_1_2(vertical_tile_24_25_to_tile_23_25_2),
		.in_wire_1_3(vertical_tile_24_25_to_tile_23_25_3),
		.out_wire_2_0(horizontal_tile_23_25_to_tile_23_24_0),
		.out_wire_2_1(horizontal_tile_23_25_to_tile_23_24_1),
		.out_wire_2_2(horizontal_tile_23_25_to_tile_23_24_2),
		.out_wire_2_3(horizontal_tile_23_25_to_tile_23_24_3),
		.in_wire_2_0(horizontal_tile_23_24_to_tile_23_25_0),
		.in_wire_2_1(horizontal_tile_23_24_to_tile_23_25_1),
		.in_wire_2_2(horizontal_tile_23_24_to_tile_23_25_2),
		.in_wire_2_3(horizontal_tile_23_24_to_tile_23_25_3),
		.out_wire_0_0(horizontal_tile_23_25_to_tile_23_26_0),
		.out_wire_0_1(horizontal_tile_23_25_to_tile_23_26_1),
		.out_wire_0_2(horizontal_tile_23_25_to_tile_23_26_2),
		.out_wire_0_3(horizontal_tile_23_25_to_tile_23_26_3),
		.in_wire_0_0(horizontal_tile_23_26_to_tile_23_25_0),
		.in_wire_0_1(horizontal_tile_23_26_to_tile_23_25_1),
		.in_wire_0_2(horizontal_tile_23_26_to_tile_23_25_2),
		.in_wire_0_3(horizontal_tile_23_26_to_tile_23_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(762)
	);

	pe_tile pe_tile_23_26(
		.out_wire_3_0(vertical_tile_23_26_to_tile_22_26_0),
		.out_wire_3_1(vertical_tile_23_26_to_tile_22_26_1),
		.out_wire_3_2(vertical_tile_23_26_to_tile_22_26_2),
		.out_wire_3_3(vertical_tile_23_26_to_tile_22_26_3),
		.in_wire_3_0(vertical_tile_22_26_to_tile_23_26_0),
		.in_wire_3_1(vertical_tile_22_26_to_tile_23_26_1),
		.in_wire_3_2(vertical_tile_22_26_to_tile_23_26_2),
		.in_wire_3_3(vertical_tile_22_26_to_tile_23_26_3),
		.out_wire_1_0(vertical_tile_23_26_to_tile_24_26_0),
		.out_wire_1_1(vertical_tile_23_26_to_tile_24_26_1),
		.out_wire_1_2(vertical_tile_23_26_to_tile_24_26_2),
		.out_wire_1_3(vertical_tile_23_26_to_tile_24_26_3),
		.in_wire_1_0(vertical_tile_24_26_to_tile_23_26_0),
		.in_wire_1_1(vertical_tile_24_26_to_tile_23_26_1),
		.in_wire_1_2(vertical_tile_24_26_to_tile_23_26_2),
		.in_wire_1_3(vertical_tile_24_26_to_tile_23_26_3),
		.out_wire_2_0(horizontal_tile_23_26_to_tile_23_25_0),
		.out_wire_2_1(horizontal_tile_23_26_to_tile_23_25_1),
		.out_wire_2_2(horizontal_tile_23_26_to_tile_23_25_2),
		.out_wire_2_3(horizontal_tile_23_26_to_tile_23_25_3),
		.in_wire_2_0(horizontal_tile_23_25_to_tile_23_26_0),
		.in_wire_2_1(horizontal_tile_23_25_to_tile_23_26_1),
		.in_wire_2_2(horizontal_tile_23_25_to_tile_23_26_2),
		.in_wire_2_3(horizontal_tile_23_25_to_tile_23_26_3),
		.out_wire_0_0(horizontal_tile_23_26_to_tile_23_27_0),
		.out_wire_0_1(horizontal_tile_23_26_to_tile_23_27_1),
		.out_wire_0_2(horizontal_tile_23_26_to_tile_23_27_2),
		.out_wire_0_3(horizontal_tile_23_26_to_tile_23_27_3),
		.in_wire_0_0(horizontal_tile_23_27_to_tile_23_26_0),
		.in_wire_0_1(horizontal_tile_23_27_to_tile_23_26_1),
		.in_wire_0_2(horizontal_tile_23_27_to_tile_23_26_2),
		.in_wire_0_3(horizontal_tile_23_27_to_tile_23_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(763)
	);

	pe_tile pe_tile_23_27(
		.out_wire_3_0(vertical_tile_23_27_to_tile_22_27_0),
		.out_wire_3_1(vertical_tile_23_27_to_tile_22_27_1),
		.out_wire_3_2(vertical_tile_23_27_to_tile_22_27_2),
		.out_wire_3_3(vertical_tile_23_27_to_tile_22_27_3),
		.in_wire_3_0(vertical_tile_22_27_to_tile_23_27_0),
		.in_wire_3_1(vertical_tile_22_27_to_tile_23_27_1),
		.in_wire_3_2(vertical_tile_22_27_to_tile_23_27_2),
		.in_wire_3_3(vertical_tile_22_27_to_tile_23_27_3),
		.out_wire_1_0(vertical_tile_23_27_to_tile_24_27_0),
		.out_wire_1_1(vertical_tile_23_27_to_tile_24_27_1),
		.out_wire_1_2(vertical_tile_23_27_to_tile_24_27_2),
		.out_wire_1_3(vertical_tile_23_27_to_tile_24_27_3),
		.in_wire_1_0(vertical_tile_24_27_to_tile_23_27_0),
		.in_wire_1_1(vertical_tile_24_27_to_tile_23_27_1),
		.in_wire_1_2(vertical_tile_24_27_to_tile_23_27_2),
		.in_wire_1_3(vertical_tile_24_27_to_tile_23_27_3),
		.out_wire_2_0(horizontal_tile_23_27_to_tile_23_26_0),
		.out_wire_2_1(horizontal_tile_23_27_to_tile_23_26_1),
		.out_wire_2_2(horizontal_tile_23_27_to_tile_23_26_2),
		.out_wire_2_3(horizontal_tile_23_27_to_tile_23_26_3),
		.in_wire_2_0(horizontal_tile_23_26_to_tile_23_27_0),
		.in_wire_2_1(horizontal_tile_23_26_to_tile_23_27_1),
		.in_wire_2_2(horizontal_tile_23_26_to_tile_23_27_2),
		.in_wire_2_3(horizontal_tile_23_26_to_tile_23_27_3),
		.out_wire_0_0(horizontal_tile_23_27_to_tile_23_28_0),
		.out_wire_0_1(horizontal_tile_23_27_to_tile_23_28_1),
		.out_wire_0_2(horizontal_tile_23_27_to_tile_23_28_2),
		.out_wire_0_3(horizontal_tile_23_27_to_tile_23_28_3),
		.in_wire_0_0(horizontal_tile_23_28_to_tile_23_27_0),
		.in_wire_0_1(horizontal_tile_23_28_to_tile_23_27_1),
		.in_wire_0_2(horizontal_tile_23_28_to_tile_23_27_2),
		.in_wire_0_3(horizontal_tile_23_28_to_tile_23_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(764)
	);

	pe_tile pe_tile_23_28(
		.out_wire_3_0(vertical_tile_23_28_to_tile_22_28_0),
		.out_wire_3_1(vertical_tile_23_28_to_tile_22_28_1),
		.out_wire_3_2(vertical_tile_23_28_to_tile_22_28_2),
		.out_wire_3_3(vertical_tile_23_28_to_tile_22_28_3),
		.in_wire_3_0(vertical_tile_22_28_to_tile_23_28_0),
		.in_wire_3_1(vertical_tile_22_28_to_tile_23_28_1),
		.in_wire_3_2(vertical_tile_22_28_to_tile_23_28_2),
		.in_wire_3_3(vertical_tile_22_28_to_tile_23_28_3),
		.out_wire_1_0(vertical_tile_23_28_to_tile_24_28_0),
		.out_wire_1_1(vertical_tile_23_28_to_tile_24_28_1),
		.out_wire_1_2(vertical_tile_23_28_to_tile_24_28_2),
		.out_wire_1_3(vertical_tile_23_28_to_tile_24_28_3),
		.in_wire_1_0(vertical_tile_24_28_to_tile_23_28_0),
		.in_wire_1_1(vertical_tile_24_28_to_tile_23_28_1),
		.in_wire_1_2(vertical_tile_24_28_to_tile_23_28_2),
		.in_wire_1_3(vertical_tile_24_28_to_tile_23_28_3),
		.out_wire_2_0(horizontal_tile_23_28_to_tile_23_27_0),
		.out_wire_2_1(horizontal_tile_23_28_to_tile_23_27_1),
		.out_wire_2_2(horizontal_tile_23_28_to_tile_23_27_2),
		.out_wire_2_3(horizontal_tile_23_28_to_tile_23_27_3),
		.in_wire_2_0(horizontal_tile_23_27_to_tile_23_28_0),
		.in_wire_2_1(horizontal_tile_23_27_to_tile_23_28_1),
		.in_wire_2_2(horizontal_tile_23_27_to_tile_23_28_2),
		.in_wire_2_3(horizontal_tile_23_27_to_tile_23_28_3),
		.out_wire_0_0(horizontal_tile_23_28_to_tile_23_29_0),
		.out_wire_0_1(horizontal_tile_23_28_to_tile_23_29_1),
		.out_wire_0_2(horizontal_tile_23_28_to_tile_23_29_2),
		.out_wire_0_3(horizontal_tile_23_28_to_tile_23_29_3),
		.in_wire_0_0(horizontal_tile_23_29_to_tile_23_28_0),
		.in_wire_0_1(horizontal_tile_23_29_to_tile_23_28_1),
		.in_wire_0_2(horizontal_tile_23_29_to_tile_23_28_2),
		.in_wire_0_3(horizontal_tile_23_29_to_tile_23_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(765)
	);

	pe_tile pe_tile_23_29(
		.out_wire_3_0(vertical_tile_23_29_to_tile_22_29_0),
		.out_wire_3_1(vertical_tile_23_29_to_tile_22_29_1),
		.out_wire_3_2(vertical_tile_23_29_to_tile_22_29_2),
		.out_wire_3_3(vertical_tile_23_29_to_tile_22_29_3),
		.in_wire_3_0(vertical_tile_22_29_to_tile_23_29_0),
		.in_wire_3_1(vertical_tile_22_29_to_tile_23_29_1),
		.in_wire_3_2(vertical_tile_22_29_to_tile_23_29_2),
		.in_wire_3_3(vertical_tile_22_29_to_tile_23_29_3),
		.out_wire_1_0(vertical_tile_23_29_to_tile_24_29_0),
		.out_wire_1_1(vertical_tile_23_29_to_tile_24_29_1),
		.out_wire_1_2(vertical_tile_23_29_to_tile_24_29_2),
		.out_wire_1_3(vertical_tile_23_29_to_tile_24_29_3),
		.in_wire_1_0(vertical_tile_24_29_to_tile_23_29_0),
		.in_wire_1_1(vertical_tile_24_29_to_tile_23_29_1),
		.in_wire_1_2(vertical_tile_24_29_to_tile_23_29_2),
		.in_wire_1_3(vertical_tile_24_29_to_tile_23_29_3),
		.out_wire_2_0(horizontal_tile_23_29_to_tile_23_28_0),
		.out_wire_2_1(horizontal_tile_23_29_to_tile_23_28_1),
		.out_wire_2_2(horizontal_tile_23_29_to_tile_23_28_2),
		.out_wire_2_3(horizontal_tile_23_29_to_tile_23_28_3),
		.in_wire_2_0(horizontal_tile_23_28_to_tile_23_29_0),
		.in_wire_2_1(horizontal_tile_23_28_to_tile_23_29_1),
		.in_wire_2_2(horizontal_tile_23_28_to_tile_23_29_2),
		.in_wire_2_3(horizontal_tile_23_28_to_tile_23_29_3),
		.out_wire_0_0(horizontal_tile_23_29_to_tile_23_30_0),
		.out_wire_0_1(horizontal_tile_23_29_to_tile_23_30_1),
		.out_wire_0_2(horizontal_tile_23_29_to_tile_23_30_2),
		.out_wire_0_3(horizontal_tile_23_29_to_tile_23_30_3),
		.in_wire_0_0(horizontal_tile_23_30_to_tile_23_29_0),
		.in_wire_0_1(horizontal_tile_23_30_to_tile_23_29_1),
		.in_wire_0_2(horizontal_tile_23_30_to_tile_23_29_2),
		.in_wire_0_3(horizontal_tile_23_30_to_tile_23_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(766)
	);

	pe_tile pe_tile_23_30(
		.out_wire_3_0(vertical_tile_23_30_to_tile_22_30_0),
		.out_wire_3_1(vertical_tile_23_30_to_tile_22_30_1),
		.out_wire_3_2(vertical_tile_23_30_to_tile_22_30_2),
		.out_wire_3_3(vertical_tile_23_30_to_tile_22_30_3),
		.in_wire_3_0(vertical_tile_22_30_to_tile_23_30_0),
		.in_wire_3_1(vertical_tile_22_30_to_tile_23_30_1),
		.in_wire_3_2(vertical_tile_22_30_to_tile_23_30_2),
		.in_wire_3_3(vertical_tile_22_30_to_tile_23_30_3),
		.out_wire_1_0(vertical_tile_23_30_to_tile_24_30_0),
		.out_wire_1_1(vertical_tile_23_30_to_tile_24_30_1),
		.out_wire_1_2(vertical_tile_23_30_to_tile_24_30_2),
		.out_wire_1_3(vertical_tile_23_30_to_tile_24_30_3),
		.in_wire_1_0(vertical_tile_24_30_to_tile_23_30_0),
		.in_wire_1_1(vertical_tile_24_30_to_tile_23_30_1),
		.in_wire_1_2(vertical_tile_24_30_to_tile_23_30_2),
		.in_wire_1_3(vertical_tile_24_30_to_tile_23_30_3),
		.out_wire_2_0(horizontal_tile_23_30_to_tile_23_29_0),
		.out_wire_2_1(horizontal_tile_23_30_to_tile_23_29_1),
		.out_wire_2_2(horizontal_tile_23_30_to_tile_23_29_2),
		.out_wire_2_3(horizontal_tile_23_30_to_tile_23_29_3),
		.in_wire_2_0(horizontal_tile_23_29_to_tile_23_30_0),
		.in_wire_2_1(horizontal_tile_23_29_to_tile_23_30_1),
		.in_wire_2_2(horizontal_tile_23_29_to_tile_23_30_2),
		.in_wire_2_3(horizontal_tile_23_29_to_tile_23_30_3),
		.out_wire_0_0(horizontal_tile_23_30_to_tile_23_31_0),
		.out_wire_0_1(horizontal_tile_23_30_to_tile_23_31_1),
		.out_wire_0_2(horizontal_tile_23_30_to_tile_23_31_2),
		.out_wire_0_3(horizontal_tile_23_30_to_tile_23_31_3),
		.in_wire_0_0(horizontal_tile_23_31_to_tile_23_30_0),
		.in_wire_0_1(horizontal_tile_23_31_to_tile_23_30_1),
		.in_wire_0_2(horizontal_tile_23_31_to_tile_23_30_2),
		.in_wire_0_3(horizontal_tile_23_31_to_tile_23_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(767)
	);

	pe_tile_right pe_tile_23_31(
		.out_wire_3_0(vertical_tile_23_31_to_tile_22_31_0),
		.out_wire_3_1(vertical_tile_23_31_to_tile_22_31_1),
		.out_wire_3_2(vertical_tile_23_31_to_tile_22_31_2),
		.out_wire_3_3(vertical_tile_23_31_to_tile_22_31_3),
		.in_wire_3_0(vertical_tile_22_31_to_tile_23_31_0),
		.in_wire_3_1(vertical_tile_22_31_to_tile_23_31_1),
		.in_wire_3_2(vertical_tile_22_31_to_tile_23_31_2),
		.in_wire_3_3(vertical_tile_22_31_to_tile_23_31_3),
		.out_wire_1_0(vertical_tile_23_31_to_tile_24_31_0),
		.out_wire_1_1(vertical_tile_23_31_to_tile_24_31_1),
		.out_wire_1_2(vertical_tile_23_31_to_tile_24_31_2),
		.out_wire_1_3(vertical_tile_23_31_to_tile_24_31_3),
		.in_wire_1_0(vertical_tile_24_31_to_tile_23_31_0),
		.in_wire_1_1(vertical_tile_24_31_to_tile_23_31_1),
		.in_wire_1_2(vertical_tile_24_31_to_tile_23_31_2),
		.in_wire_1_3(vertical_tile_24_31_to_tile_23_31_3),
		.out_wire_2_0(horizontal_tile_23_31_to_tile_23_30_0),
		.out_wire_2_1(horizontal_tile_23_31_to_tile_23_30_1),
		.out_wire_2_2(horizontal_tile_23_31_to_tile_23_30_2),
		.out_wire_2_3(horizontal_tile_23_31_to_tile_23_30_3),
		.in_wire_2_0(horizontal_tile_23_30_to_tile_23_31_0),
		.in_wire_2_1(horizontal_tile_23_30_to_tile_23_31_1),
		.in_wire_2_2(horizontal_tile_23_30_to_tile_23_31_2),
		.in_wire_2_3(horizontal_tile_23_30_to_tile_23_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(768)
	);

	pe_tile_left pe_tile_24_0(
		.out_wire_3_0(vertical_tile_24_0_to_tile_23_0_0),
		.out_wire_3_1(vertical_tile_24_0_to_tile_23_0_1),
		.out_wire_3_2(vertical_tile_24_0_to_tile_23_0_2),
		.out_wire_3_3(vertical_tile_24_0_to_tile_23_0_3),
		.in_wire_3_0(vertical_tile_23_0_to_tile_24_0_0),
		.in_wire_3_1(vertical_tile_23_0_to_tile_24_0_1),
		.in_wire_3_2(vertical_tile_23_0_to_tile_24_0_2),
		.in_wire_3_3(vertical_tile_23_0_to_tile_24_0_3),
		.out_wire_1_0(vertical_tile_24_0_to_tile_25_0_0),
		.out_wire_1_1(vertical_tile_24_0_to_tile_25_0_1),
		.out_wire_1_2(vertical_tile_24_0_to_tile_25_0_2),
		.out_wire_1_3(vertical_tile_24_0_to_tile_25_0_3),
		.in_wire_1_0(vertical_tile_25_0_to_tile_24_0_0),
		.in_wire_1_1(vertical_tile_25_0_to_tile_24_0_1),
		.in_wire_1_2(vertical_tile_25_0_to_tile_24_0_2),
		.in_wire_1_3(vertical_tile_25_0_to_tile_24_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_24_0_to_tile_24_1_0),
		.out_wire_0_1(horizontal_tile_24_0_to_tile_24_1_1),
		.out_wire_0_2(horizontal_tile_24_0_to_tile_24_1_2),
		.out_wire_0_3(horizontal_tile_24_0_to_tile_24_1_3),
		.in_wire_0_0(horizontal_tile_24_1_to_tile_24_0_0),
		.in_wire_0_1(horizontal_tile_24_1_to_tile_24_0_1),
		.in_wire_0_2(horizontal_tile_24_1_to_tile_24_0_2),
		.in_wire_0_3(horizontal_tile_24_1_to_tile_24_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(769)
	);

	pe_tile pe_tile_24_1(
		.out_wire_3_0(vertical_tile_24_1_to_tile_23_1_0),
		.out_wire_3_1(vertical_tile_24_1_to_tile_23_1_1),
		.out_wire_3_2(vertical_tile_24_1_to_tile_23_1_2),
		.out_wire_3_3(vertical_tile_24_1_to_tile_23_1_3),
		.in_wire_3_0(vertical_tile_23_1_to_tile_24_1_0),
		.in_wire_3_1(vertical_tile_23_1_to_tile_24_1_1),
		.in_wire_3_2(vertical_tile_23_1_to_tile_24_1_2),
		.in_wire_3_3(vertical_tile_23_1_to_tile_24_1_3),
		.out_wire_1_0(vertical_tile_24_1_to_tile_25_1_0),
		.out_wire_1_1(vertical_tile_24_1_to_tile_25_1_1),
		.out_wire_1_2(vertical_tile_24_1_to_tile_25_1_2),
		.out_wire_1_3(vertical_tile_24_1_to_tile_25_1_3),
		.in_wire_1_0(vertical_tile_25_1_to_tile_24_1_0),
		.in_wire_1_1(vertical_tile_25_1_to_tile_24_1_1),
		.in_wire_1_2(vertical_tile_25_1_to_tile_24_1_2),
		.in_wire_1_3(vertical_tile_25_1_to_tile_24_1_3),
		.out_wire_2_0(horizontal_tile_24_1_to_tile_24_0_0),
		.out_wire_2_1(horizontal_tile_24_1_to_tile_24_0_1),
		.out_wire_2_2(horizontal_tile_24_1_to_tile_24_0_2),
		.out_wire_2_3(horizontal_tile_24_1_to_tile_24_0_3),
		.in_wire_2_0(horizontal_tile_24_0_to_tile_24_1_0),
		.in_wire_2_1(horizontal_tile_24_0_to_tile_24_1_1),
		.in_wire_2_2(horizontal_tile_24_0_to_tile_24_1_2),
		.in_wire_2_3(horizontal_tile_24_0_to_tile_24_1_3),
		.out_wire_0_0(horizontal_tile_24_1_to_tile_24_2_0),
		.out_wire_0_1(horizontal_tile_24_1_to_tile_24_2_1),
		.out_wire_0_2(horizontal_tile_24_1_to_tile_24_2_2),
		.out_wire_0_3(horizontal_tile_24_1_to_tile_24_2_3),
		.in_wire_0_0(horizontal_tile_24_2_to_tile_24_1_0),
		.in_wire_0_1(horizontal_tile_24_2_to_tile_24_1_1),
		.in_wire_0_2(horizontal_tile_24_2_to_tile_24_1_2),
		.in_wire_0_3(horizontal_tile_24_2_to_tile_24_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(770)
	);

	pe_tile pe_tile_24_2(
		.out_wire_3_0(vertical_tile_24_2_to_tile_23_2_0),
		.out_wire_3_1(vertical_tile_24_2_to_tile_23_2_1),
		.out_wire_3_2(vertical_tile_24_2_to_tile_23_2_2),
		.out_wire_3_3(vertical_tile_24_2_to_tile_23_2_3),
		.in_wire_3_0(vertical_tile_23_2_to_tile_24_2_0),
		.in_wire_3_1(vertical_tile_23_2_to_tile_24_2_1),
		.in_wire_3_2(vertical_tile_23_2_to_tile_24_2_2),
		.in_wire_3_3(vertical_tile_23_2_to_tile_24_2_3),
		.out_wire_1_0(vertical_tile_24_2_to_tile_25_2_0),
		.out_wire_1_1(vertical_tile_24_2_to_tile_25_2_1),
		.out_wire_1_2(vertical_tile_24_2_to_tile_25_2_2),
		.out_wire_1_3(vertical_tile_24_2_to_tile_25_2_3),
		.in_wire_1_0(vertical_tile_25_2_to_tile_24_2_0),
		.in_wire_1_1(vertical_tile_25_2_to_tile_24_2_1),
		.in_wire_1_2(vertical_tile_25_2_to_tile_24_2_2),
		.in_wire_1_3(vertical_tile_25_2_to_tile_24_2_3),
		.out_wire_2_0(horizontal_tile_24_2_to_tile_24_1_0),
		.out_wire_2_1(horizontal_tile_24_2_to_tile_24_1_1),
		.out_wire_2_2(horizontal_tile_24_2_to_tile_24_1_2),
		.out_wire_2_3(horizontal_tile_24_2_to_tile_24_1_3),
		.in_wire_2_0(horizontal_tile_24_1_to_tile_24_2_0),
		.in_wire_2_1(horizontal_tile_24_1_to_tile_24_2_1),
		.in_wire_2_2(horizontal_tile_24_1_to_tile_24_2_2),
		.in_wire_2_3(horizontal_tile_24_1_to_tile_24_2_3),
		.out_wire_0_0(horizontal_tile_24_2_to_tile_24_3_0),
		.out_wire_0_1(horizontal_tile_24_2_to_tile_24_3_1),
		.out_wire_0_2(horizontal_tile_24_2_to_tile_24_3_2),
		.out_wire_0_3(horizontal_tile_24_2_to_tile_24_3_3),
		.in_wire_0_0(horizontal_tile_24_3_to_tile_24_2_0),
		.in_wire_0_1(horizontal_tile_24_3_to_tile_24_2_1),
		.in_wire_0_2(horizontal_tile_24_3_to_tile_24_2_2),
		.in_wire_0_3(horizontal_tile_24_3_to_tile_24_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(771)
	);

	pe_tile pe_tile_24_3(
		.out_wire_3_0(vertical_tile_24_3_to_tile_23_3_0),
		.out_wire_3_1(vertical_tile_24_3_to_tile_23_3_1),
		.out_wire_3_2(vertical_tile_24_3_to_tile_23_3_2),
		.out_wire_3_3(vertical_tile_24_3_to_tile_23_3_3),
		.in_wire_3_0(vertical_tile_23_3_to_tile_24_3_0),
		.in_wire_3_1(vertical_tile_23_3_to_tile_24_3_1),
		.in_wire_3_2(vertical_tile_23_3_to_tile_24_3_2),
		.in_wire_3_3(vertical_tile_23_3_to_tile_24_3_3),
		.out_wire_1_0(vertical_tile_24_3_to_tile_25_3_0),
		.out_wire_1_1(vertical_tile_24_3_to_tile_25_3_1),
		.out_wire_1_2(vertical_tile_24_3_to_tile_25_3_2),
		.out_wire_1_3(vertical_tile_24_3_to_tile_25_3_3),
		.in_wire_1_0(vertical_tile_25_3_to_tile_24_3_0),
		.in_wire_1_1(vertical_tile_25_3_to_tile_24_3_1),
		.in_wire_1_2(vertical_tile_25_3_to_tile_24_3_2),
		.in_wire_1_3(vertical_tile_25_3_to_tile_24_3_3),
		.out_wire_2_0(horizontal_tile_24_3_to_tile_24_2_0),
		.out_wire_2_1(horizontal_tile_24_3_to_tile_24_2_1),
		.out_wire_2_2(horizontal_tile_24_3_to_tile_24_2_2),
		.out_wire_2_3(horizontal_tile_24_3_to_tile_24_2_3),
		.in_wire_2_0(horizontal_tile_24_2_to_tile_24_3_0),
		.in_wire_2_1(horizontal_tile_24_2_to_tile_24_3_1),
		.in_wire_2_2(horizontal_tile_24_2_to_tile_24_3_2),
		.in_wire_2_3(horizontal_tile_24_2_to_tile_24_3_3),
		.out_wire_0_0(horizontal_tile_24_3_to_tile_24_4_0),
		.out_wire_0_1(horizontal_tile_24_3_to_tile_24_4_1),
		.out_wire_0_2(horizontal_tile_24_3_to_tile_24_4_2),
		.out_wire_0_3(horizontal_tile_24_3_to_tile_24_4_3),
		.in_wire_0_0(horizontal_tile_24_4_to_tile_24_3_0),
		.in_wire_0_1(horizontal_tile_24_4_to_tile_24_3_1),
		.in_wire_0_2(horizontal_tile_24_4_to_tile_24_3_2),
		.in_wire_0_3(horizontal_tile_24_4_to_tile_24_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(772)
	);

	pe_tile pe_tile_24_4(
		.out_wire_3_0(vertical_tile_24_4_to_tile_23_4_0),
		.out_wire_3_1(vertical_tile_24_4_to_tile_23_4_1),
		.out_wire_3_2(vertical_tile_24_4_to_tile_23_4_2),
		.out_wire_3_3(vertical_tile_24_4_to_tile_23_4_3),
		.in_wire_3_0(vertical_tile_23_4_to_tile_24_4_0),
		.in_wire_3_1(vertical_tile_23_4_to_tile_24_4_1),
		.in_wire_3_2(vertical_tile_23_4_to_tile_24_4_2),
		.in_wire_3_3(vertical_tile_23_4_to_tile_24_4_3),
		.out_wire_1_0(vertical_tile_24_4_to_tile_25_4_0),
		.out_wire_1_1(vertical_tile_24_4_to_tile_25_4_1),
		.out_wire_1_2(vertical_tile_24_4_to_tile_25_4_2),
		.out_wire_1_3(vertical_tile_24_4_to_tile_25_4_3),
		.in_wire_1_0(vertical_tile_25_4_to_tile_24_4_0),
		.in_wire_1_1(vertical_tile_25_4_to_tile_24_4_1),
		.in_wire_1_2(vertical_tile_25_4_to_tile_24_4_2),
		.in_wire_1_3(vertical_tile_25_4_to_tile_24_4_3),
		.out_wire_2_0(horizontal_tile_24_4_to_tile_24_3_0),
		.out_wire_2_1(horizontal_tile_24_4_to_tile_24_3_1),
		.out_wire_2_2(horizontal_tile_24_4_to_tile_24_3_2),
		.out_wire_2_3(horizontal_tile_24_4_to_tile_24_3_3),
		.in_wire_2_0(horizontal_tile_24_3_to_tile_24_4_0),
		.in_wire_2_1(horizontal_tile_24_3_to_tile_24_4_1),
		.in_wire_2_2(horizontal_tile_24_3_to_tile_24_4_2),
		.in_wire_2_3(horizontal_tile_24_3_to_tile_24_4_3),
		.out_wire_0_0(horizontal_tile_24_4_to_tile_24_5_0),
		.out_wire_0_1(horizontal_tile_24_4_to_tile_24_5_1),
		.out_wire_0_2(horizontal_tile_24_4_to_tile_24_5_2),
		.out_wire_0_3(horizontal_tile_24_4_to_tile_24_5_3),
		.in_wire_0_0(horizontal_tile_24_5_to_tile_24_4_0),
		.in_wire_0_1(horizontal_tile_24_5_to_tile_24_4_1),
		.in_wire_0_2(horizontal_tile_24_5_to_tile_24_4_2),
		.in_wire_0_3(horizontal_tile_24_5_to_tile_24_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(773)
	);

	pe_tile pe_tile_24_5(
		.out_wire_3_0(vertical_tile_24_5_to_tile_23_5_0),
		.out_wire_3_1(vertical_tile_24_5_to_tile_23_5_1),
		.out_wire_3_2(vertical_tile_24_5_to_tile_23_5_2),
		.out_wire_3_3(vertical_tile_24_5_to_tile_23_5_3),
		.in_wire_3_0(vertical_tile_23_5_to_tile_24_5_0),
		.in_wire_3_1(vertical_tile_23_5_to_tile_24_5_1),
		.in_wire_3_2(vertical_tile_23_5_to_tile_24_5_2),
		.in_wire_3_3(vertical_tile_23_5_to_tile_24_5_3),
		.out_wire_1_0(vertical_tile_24_5_to_tile_25_5_0),
		.out_wire_1_1(vertical_tile_24_5_to_tile_25_5_1),
		.out_wire_1_2(vertical_tile_24_5_to_tile_25_5_2),
		.out_wire_1_3(vertical_tile_24_5_to_tile_25_5_3),
		.in_wire_1_0(vertical_tile_25_5_to_tile_24_5_0),
		.in_wire_1_1(vertical_tile_25_5_to_tile_24_5_1),
		.in_wire_1_2(vertical_tile_25_5_to_tile_24_5_2),
		.in_wire_1_3(vertical_tile_25_5_to_tile_24_5_3),
		.out_wire_2_0(horizontal_tile_24_5_to_tile_24_4_0),
		.out_wire_2_1(horizontal_tile_24_5_to_tile_24_4_1),
		.out_wire_2_2(horizontal_tile_24_5_to_tile_24_4_2),
		.out_wire_2_3(horizontal_tile_24_5_to_tile_24_4_3),
		.in_wire_2_0(horizontal_tile_24_4_to_tile_24_5_0),
		.in_wire_2_1(horizontal_tile_24_4_to_tile_24_5_1),
		.in_wire_2_2(horizontal_tile_24_4_to_tile_24_5_2),
		.in_wire_2_3(horizontal_tile_24_4_to_tile_24_5_3),
		.out_wire_0_0(horizontal_tile_24_5_to_tile_24_6_0),
		.out_wire_0_1(horizontal_tile_24_5_to_tile_24_6_1),
		.out_wire_0_2(horizontal_tile_24_5_to_tile_24_6_2),
		.out_wire_0_3(horizontal_tile_24_5_to_tile_24_6_3),
		.in_wire_0_0(horizontal_tile_24_6_to_tile_24_5_0),
		.in_wire_0_1(horizontal_tile_24_6_to_tile_24_5_1),
		.in_wire_0_2(horizontal_tile_24_6_to_tile_24_5_2),
		.in_wire_0_3(horizontal_tile_24_6_to_tile_24_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(774)
	);

	pe_tile pe_tile_24_6(
		.out_wire_3_0(vertical_tile_24_6_to_tile_23_6_0),
		.out_wire_3_1(vertical_tile_24_6_to_tile_23_6_1),
		.out_wire_3_2(vertical_tile_24_6_to_tile_23_6_2),
		.out_wire_3_3(vertical_tile_24_6_to_tile_23_6_3),
		.in_wire_3_0(vertical_tile_23_6_to_tile_24_6_0),
		.in_wire_3_1(vertical_tile_23_6_to_tile_24_6_1),
		.in_wire_3_2(vertical_tile_23_6_to_tile_24_6_2),
		.in_wire_3_3(vertical_tile_23_6_to_tile_24_6_3),
		.out_wire_1_0(vertical_tile_24_6_to_tile_25_6_0),
		.out_wire_1_1(vertical_tile_24_6_to_tile_25_6_1),
		.out_wire_1_2(vertical_tile_24_6_to_tile_25_6_2),
		.out_wire_1_3(vertical_tile_24_6_to_tile_25_6_3),
		.in_wire_1_0(vertical_tile_25_6_to_tile_24_6_0),
		.in_wire_1_1(vertical_tile_25_6_to_tile_24_6_1),
		.in_wire_1_2(vertical_tile_25_6_to_tile_24_6_2),
		.in_wire_1_3(vertical_tile_25_6_to_tile_24_6_3),
		.out_wire_2_0(horizontal_tile_24_6_to_tile_24_5_0),
		.out_wire_2_1(horizontal_tile_24_6_to_tile_24_5_1),
		.out_wire_2_2(horizontal_tile_24_6_to_tile_24_5_2),
		.out_wire_2_3(horizontal_tile_24_6_to_tile_24_5_3),
		.in_wire_2_0(horizontal_tile_24_5_to_tile_24_6_0),
		.in_wire_2_1(horizontal_tile_24_5_to_tile_24_6_1),
		.in_wire_2_2(horizontal_tile_24_5_to_tile_24_6_2),
		.in_wire_2_3(horizontal_tile_24_5_to_tile_24_6_3),
		.out_wire_0_0(horizontal_tile_24_6_to_tile_24_7_0),
		.out_wire_0_1(horizontal_tile_24_6_to_tile_24_7_1),
		.out_wire_0_2(horizontal_tile_24_6_to_tile_24_7_2),
		.out_wire_0_3(horizontal_tile_24_6_to_tile_24_7_3),
		.in_wire_0_0(horizontal_tile_24_7_to_tile_24_6_0),
		.in_wire_0_1(horizontal_tile_24_7_to_tile_24_6_1),
		.in_wire_0_2(horizontal_tile_24_7_to_tile_24_6_2),
		.in_wire_0_3(horizontal_tile_24_7_to_tile_24_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(775)
	);

	pe_tile pe_tile_24_7(
		.out_wire_3_0(vertical_tile_24_7_to_tile_23_7_0),
		.out_wire_3_1(vertical_tile_24_7_to_tile_23_7_1),
		.out_wire_3_2(vertical_tile_24_7_to_tile_23_7_2),
		.out_wire_3_3(vertical_tile_24_7_to_tile_23_7_3),
		.in_wire_3_0(vertical_tile_23_7_to_tile_24_7_0),
		.in_wire_3_1(vertical_tile_23_7_to_tile_24_7_1),
		.in_wire_3_2(vertical_tile_23_7_to_tile_24_7_2),
		.in_wire_3_3(vertical_tile_23_7_to_tile_24_7_3),
		.out_wire_1_0(vertical_tile_24_7_to_tile_25_7_0),
		.out_wire_1_1(vertical_tile_24_7_to_tile_25_7_1),
		.out_wire_1_2(vertical_tile_24_7_to_tile_25_7_2),
		.out_wire_1_3(vertical_tile_24_7_to_tile_25_7_3),
		.in_wire_1_0(vertical_tile_25_7_to_tile_24_7_0),
		.in_wire_1_1(vertical_tile_25_7_to_tile_24_7_1),
		.in_wire_1_2(vertical_tile_25_7_to_tile_24_7_2),
		.in_wire_1_3(vertical_tile_25_7_to_tile_24_7_3),
		.out_wire_2_0(horizontal_tile_24_7_to_tile_24_6_0),
		.out_wire_2_1(horizontal_tile_24_7_to_tile_24_6_1),
		.out_wire_2_2(horizontal_tile_24_7_to_tile_24_6_2),
		.out_wire_2_3(horizontal_tile_24_7_to_tile_24_6_3),
		.in_wire_2_0(horizontal_tile_24_6_to_tile_24_7_0),
		.in_wire_2_1(horizontal_tile_24_6_to_tile_24_7_1),
		.in_wire_2_2(horizontal_tile_24_6_to_tile_24_7_2),
		.in_wire_2_3(horizontal_tile_24_6_to_tile_24_7_3),
		.out_wire_0_0(horizontal_tile_24_7_to_tile_24_8_0),
		.out_wire_0_1(horizontal_tile_24_7_to_tile_24_8_1),
		.out_wire_0_2(horizontal_tile_24_7_to_tile_24_8_2),
		.out_wire_0_3(horizontal_tile_24_7_to_tile_24_8_3),
		.in_wire_0_0(horizontal_tile_24_8_to_tile_24_7_0),
		.in_wire_0_1(horizontal_tile_24_8_to_tile_24_7_1),
		.in_wire_0_2(horizontal_tile_24_8_to_tile_24_7_2),
		.in_wire_0_3(horizontal_tile_24_8_to_tile_24_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(776)
	);

	pe_tile pe_tile_24_8(
		.out_wire_3_0(vertical_tile_24_8_to_tile_23_8_0),
		.out_wire_3_1(vertical_tile_24_8_to_tile_23_8_1),
		.out_wire_3_2(vertical_tile_24_8_to_tile_23_8_2),
		.out_wire_3_3(vertical_tile_24_8_to_tile_23_8_3),
		.in_wire_3_0(vertical_tile_23_8_to_tile_24_8_0),
		.in_wire_3_1(vertical_tile_23_8_to_tile_24_8_1),
		.in_wire_3_2(vertical_tile_23_8_to_tile_24_8_2),
		.in_wire_3_3(vertical_tile_23_8_to_tile_24_8_3),
		.out_wire_1_0(vertical_tile_24_8_to_tile_25_8_0),
		.out_wire_1_1(vertical_tile_24_8_to_tile_25_8_1),
		.out_wire_1_2(vertical_tile_24_8_to_tile_25_8_2),
		.out_wire_1_3(vertical_tile_24_8_to_tile_25_8_3),
		.in_wire_1_0(vertical_tile_25_8_to_tile_24_8_0),
		.in_wire_1_1(vertical_tile_25_8_to_tile_24_8_1),
		.in_wire_1_2(vertical_tile_25_8_to_tile_24_8_2),
		.in_wire_1_3(vertical_tile_25_8_to_tile_24_8_3),
		.out_wire_2_0(horizontal_tile_24_8_to_tile_24_7_0),
		.out_wire_2_1(horizontal_tile_24_8_to_tile_24_7_1),
		.out_wire_2_2(horizontal_tile_24_8_to_tile_24_7_2),
		.out_wire_2_3(horizontal_tile_24_8_to_tile_24_7_3),
		.in_wire_2_0(horizontal_tile_24_7_to_tile_24_8_0),
		.in_wire_2_1(horizontal_tile_24_7_to_tile_24_8_1),
		.in_wire_2_2(horizontal_tile_24_7_to_tile_24_8_2),
		.in_wire_2_3(horizontal_tile_24_7_to_tile_24_8_3),
		.out_wire_0_0(horizontal_tile_24_8_to_tile_24_9_0),
		.out_wire_0_1(horizontal_tile_24_8_to_tile_24_9_1),
		.out_wire_0_2(horizontal_tile_24_8_to_tile_24_9_2),
		.out_wire_0_3(horizontal_tile_24_8_to_tile_24_9_3),
		.in_wire_0_0(horizontal_tile_24_9_to_tile_24_8_0),
		.in_wire_0_1(horizontal_tile_24_9_to_tile_24_8_1),
		.in_wire_0_2(horizontal_tile_24_9_to_tile_24_8_2),
		.in_wire_0_3(horizontal_tile_24_9_to_tile_24_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(777)
	);

	pe_tile pe_tile_24_9(
		.out_wire_3_0(vertical_tile_24_9_to_tile_23_9_0),
		.out_wire_3_1(vertical_tile_24_9_to_tile_23_9_1),
		.out_wire_3_2(vertical_tile_24_9_to_tile_23_9_2),
		.out_wire_3_3(vertical_tile_24_9_to_tile_23_9_3),
		.in_wire_3_0(vertical_tile_23_9_to_tile_24_9_0),
		.in_wire_3_1(vertical_tile_23_9_to_tile_24_9_1),
		.in_wire_3_2(vertical_tile_23_9_to_tile_24_9_2),
		.in_wire_3_3(vertical_tile_23_9_to_tile_24_9_3),
		.out_wire_1_0(vertical_tile_24_9_to_tile_25_9_0),
		.out_wire_1_1(vertical_tile_24_9_to_tile_25_9_1),
		.out_wire_1_2(vertical_tile_24_9_to_tile_25_9_2),
		.out_wire_1_3(vertical_tile_24_9_to_tile_25_9_3),
		.in_wire_1_0(vertical_tile_25_9_to_tile_24_9_0),
		.in_wire_1_1(vertical_tile_25_9_to_tile_24_9_1),
		.in_wire_1_2(vertical_tile_25_9_to_tile_24_9_2),
		.in_wire_1_3(vertical_tile_25_9_to_tile_24_9_3),
		.out_wire_2_0(horizontal_tile_24_9_to_tile_24_8_0),
		.out_wire_2_1(horizontal_tile_24_9_to_tile_24_8_1),
		.out_wire_2_2(horizontal_tile_24_9_to_tile_24_8_2),
		.out_wire_2_3(horizontal_tile_24_9_to_tile_24_8_3),
		.in_wire_2_0(horizontal_tile_24_8_to_tile_24_9_0),
		.in_wire_2_1(horizontal_tile_24_8_to_tile_24_9_1),
		.in_wire_2_2(horizontal_tile_24_8_to_tile_24_9_2),
		.in_wire_2_3(horizontal_tile_24_8_to_tile_24_9_3),
		.out_wire_0_0(horizontal_tile_24_9_to_tile_24_10_0),
		.out_wire_0_1(horizontal_tile_24_9_to_tile_24_10_1),
		.out_wire_0_2(horizontal_tile_24_9_to_tile_24_10_2),
		.out_wire_0_3(horizontal_tile_24_9_to_tile_24_10_3),
		.in_wire_0_0(horizontal_tile_24_10_to_tile_24_9_0),
		.in_wire_0_1(horizontal_tile_24_10_to_tile_24_9_1),
		.in_wire_0_2(horizontal_tile_24_10_to_tile_24_9_2),
		.in_wire_0_3(horizontal_tile_24_10_to_tile_24_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(778)
	);

	pe_tile pe_tile_24_10(
		.out_wire_3_0(vertical_tile_24_10_to_tile_23_10_0),
		.out_wire_3_1(vertical_tile_24_10_to_tile_23_10_1),
		.out_wire_3_2(vertical_tile_24_10_to_tile_23_10_2),
		.out_wire_3_3(vertical_tile_24_10_to_tile_23_10_3),
		.in_wire_3_0(vertical_tile_23_10_to_tile_24_10_0),
		.in_wire_3_1(vertical_tile_23_10_to_tile_24_10_1),
		.in_wire_3_2(vertical_tile_23_10_to_tile_24_10_2),
		.in_wire_3_3(vertical_tile_23_10_to_tile_24_10_3),
		.out_wire_1_0(vertical_tile_24_10_to_tile_25_10_0),
		.out_wire_1_1(vertical_tile_24_10_to_tile_25_10_1),
		.out_wire_1_2(vertical_tile_24_10_to_tile_25_10_2),
		.out_wire_1_3(vertical_tile_24_10_to_tile_25_10_3),
		.in_wire_1_0(vertical_tile_25_10_to_tile_24_10_0),
		.in_wire_1_1(vertical_tile_25_10_to_tile_24_10_1),
		.in_wire_1_2(vertical_tile_25_10_to_tile_24_10_2),
		.in_wire_1_3(vertical_tile_25_10_to_tile_24_10_3),
		.out_wire_2_0(horizontal_tile_24_10_to_tile_24_9_0),
		.out_wire_2_1(horizontal_tile_24_10_to_tile_24_9_1),
		.out_wire_2_2(horizontal_tile_24_10_to_tile_24_9_2),
		.out_wire_2_3(horizontal_tile_24_10_to_tile_24_9_3),
		.in_wire_2_0(horizontal_tile_24_9_to_tile_24_10_0),
		.in_wire_2_1(horizontal_tile_24_9_to_tile_24_10_1),
		.in_wire_2_2(horizontal_tile_24_9_to_tile_24_10_2),
		.in_wire_2_3(horizontal_tile_24_9_to_tile_24_10_3),
		.out_wire_0_0(horizontal_tile_24_10_to_tile_24_11_0),
		.out_wire_0_1(horizontal_tile_24_10_to_tile_24_11_1),
		.out_wire_0_2(horizontal_tile_24_10_to_tile_24_11_2),
		.out_wire_0_3(horizontal_tile_24_10_to_tile_24_11_3),
		.in_wire_0_0(horizontal_tile_24_11_to_tile_24_10_0),
		.in_wire_0_1(horizontal_tile_24_11_to_tile_24_10_1),
		.in_wire_0_2(horizontal_tile_24_11_to_tile_24_10_2),
		.in_wire_0_3(horizontal_tile_24_11_to_tile_24_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(779)
	);

	pe_tile pe_tile_24_11(
		.out_wire_3_0(vertical_tile_24_11_to_tile_23_11_0),
		.out_wire_3_1(vertical_tile_24_11_to_tile_23_11_1),
		.out_wire_3_2(vertical_tile_24_11_to_tile_23_11_2),
		.out_wire_3_3(vertical_tile_24_11_to_tile_23_11_3),
		.in_wire_3_0(vertical_tile_23_11_to_tile_24_11_0),
		.in_wire_3_1(vertical_tile_23_11_to_tile_24_11_1),
		.in_wire_3_2(vertical_tile_23_11_to_tile_24_11_2),
		.in_wire_3_3(vertical_tile_23_11_to_tile_24_11_3),
		.out_wire_1_0(vertical_tile_24_11_to_tile_25_11_0),
		.out_wire_1_1(vertical_tile_24_11_to_tile_25_11_1),
		.out_wire_1_2(vertical_tile_24_11_to_tile_25_11_2),
		.out_wire_1_3(vertical_tile_24_11_to_tile_25_11_3),
		.in_wire_1_0(vertical_tile_25_11_to_tile_24_11_0),
		.in_wire_1_1(vertical_tile_25_11_to_tile_24_11_1),
		.in_wire_1_2(vertical_tile_25_11_to_tile_24_11_2),
		.in_wire_1_3(vertical_tile_25_11_to_tile_24_11_3),
		.out_wire_2_0(horizontal_tile_24_11_to_tile_24_10_0),
		.out_wire_2_1(horizontal_tile_24_11_to_tile_24_10_1),
		.out_wire_2_2(horizontal_tile_24_11_to_tile_24_10_2),
		.out_wire_2_3(horizontal_tile_24_11_to_tile_24_10_3),
		.in_wire_2_0(horizontal_tile_24_10_to_tile_24_11_0),
		.in_wire_2_1(horizontal_tile_24_10_to_tile_24_11_1),
		.in_wire_2_2(horizontal_tile_24_10_to_tile_24_11_2),
		.in_wire_2_3(horizontal_tile_24_10_to_tile_24_11_3),
		.out_wire_0_0(horizontal_tile_24_11_to_tile_24_12_0),
		.out_wire_0_1(horizontal_tile_24_11_to_tile_24_12_1),
		.out_wire_0_2(horizontal_tile_24_11_to_tile_24_12_2),
		.out_wire_0_3(horizontal_tile_24_11_to_tile_24_12_3),
		.in_wire_0_0(horizontal_tile_24_12_to_tile_24_11_0),
		.in_wire_0_1(horizontal_tile_24_12_to_tile_24_11_1),
		.in_wire_0_2(horizontal_tile_24_12_to_tile_24_11_2),
		.in_wire_0_3(horizontal_tile_24_12_to_tile_24_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(780)
	);

	pe_tile pe_tile_24_12(
		.out_wire_3_0(vertical_tile_24_12_to_tile_23_12_0),
		.out_wire_3_1(vertical_tile_24_12_to_tile_23_12_1),
		.out_wire_3_2(vertical_tile_24_12_to_tile_23_12_2),
		.out_wire_3_3(vertical_tile_24_12_to_tile_23_12_3),
		.in_wire_3_0(vertical_tile_23_12_to_tile_24_12_0),
		.in_wire_3_1(vertical_tile_23_12_to_tile_24_12_1),
		.in_wire_3_2(vertical_tile_23_12_to_tile_24_12_2),
		.in_wire_3_3(vertical_tile_23_12_to_tile_24_12_3),
		.out_wire_1_0(vertical_tile_24_12_to_tile_25_12_0),
		.out_wire_1_1(vertical_tile_24_12_to_tile_25_12_1),
		.out_wire_1_2(vertical_tile_24_12_to_tile_25_12_2),
		.out_wire_1_3(vertical_tile_24_12_to_tile_25_12_3),
		.in_wire_1_0(vertical_tile_25_12_to_tile_24_12_0),
		.in_wire_1_1(vertical_tile_25_12_to_tile_24_12_1),
		.in_wire_1_2(vertical_tile_25_12_to_tile_24_12_2),
		.in_wire_1_3(vertical_tile_25_12_to_tile_24_12_3),
		.out_wire_2_0(horizontal_tile_24_12_to_tile_24_11_0),
		.out_wire_2_1(horizontal_tile_24_12_to_tile_24_11_1),
		.out_wire_2_2(horizontal_tile_24_12_to_tile_24_11_2),
		.out_wire_2_3(horizontal_tile_24_12_to_tile_24_11_3),
		.in_wire_2_0(horizontal_tile_24_11_to_tile_24_12_0),
		.in_wire_2_1(horizontal_tile_24_11_to_tile_24_12_1),
		.in_wire_2_2(horizontal_tile_24_11_to_tile_24_12_2),
		.in_wire_2_3(horizontal_tile_24_11_to_tile_24_12_3),
		.out_wire_0_0(horizontal_tile_24_12_to_tile_24_13_0),
		.out_wire_0_1(horizontal_tile_24_12_to_tile_24_13_1),
		.out_wire_0_2(horizontal_tile_24_12_to_tile_24_13_2),
		.out_wire_0_3(horizontal_tile_24_12_to_tile_24_13_3),
		.in_wire_0_0(horizontal_tile_24_13_to_tile_24_12_0),
		.in_wire_0_1(horizontal_tile_24_13_to_tile_24_12_1),
		.in_wire_0_2(horizontal_tile_24_13_to_tile_24_12_2),
		.in_wire_0_3(horizontal_tile_24_13_to_tile_24_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(781)
	);

	pe_tile pe_tile_24_13(
		.out_wire_3_0(vertical_tile_24_13_to_tile_23_13_0),
		.out_wire_3_1(vertical_tile_24_13_to_tile_23_13_1),
		.out_wire_3_2(vertical_tile_24_13_to_tile_23_13_2),
		.out_wire_3_3(vertical_tile_24_13_to_tile_23_13_3),
		.in_wire_3_0(vertical_tile_23_13_to_tile_24_13_0),
		.in_wire_3_1(vertical_tile_23_13_to_tile_24_13_1),
		.in_wire_3_2(vertical_tile_23_13_to_tile_24_13_2),
		.in_wire_3_3(vertical_tile_23_13_to_tile_24_13_3),
		.out_wire_1_0(vertical_tile_24_13_to_tile_25_13_0),
		.out_wire_1_1(vertical_tile_24_13_to_tile_25_13_1),
		.out_wire_1_2(vertical_tile_24_13_to_tile_25_13_2),
		.out_wire_1_3(vertical_tile_24_13_to_tile_25_13_3),
		.in_wire_1_0(vertical_tile_25_13_to_tile_24_13_0),
		.in_wire_1_1(vertical_tile_25_13_to_tile_24_13_1),
		.in_wire_1_2(vertical_tile_25_13_to_tile_24_13_2),
		.in_wire_1_3(vertical_tile_25_13_to_tile_24_13_3),
		.out_wire_2_0(horizontal_tile_24_13_to_tile_24_12_0),
		.out_wire_2_1(horizontal_tile_24_13_to_tile_24_12_1),
		.out_wire_2_2(horizontal_tile_24_13_to_tile_24_12_2),
		.out_wire_2_3(horizontal_tile_24_13_to_tile_24_12_3),
		.in_wire_2_0(horizontal_tile_24_12_to_tile_24_13_0),
		.in_wire_2_1(horizontal_tile_24_12_to_tile_24_13_1),
		.in_wire_2_2(horizontal_tile_24_12_to_tile_24_13_2),
		.in_wire_2_3(horizontal_tile_24_12_to_tile_24_13_3),
		.out_wire_0_0(horizontal_tile_24_13_to_tile_24_14_0),
		.out_wire_0_1(horizontal_tile_24_13_to_tile_24_14_1),
		.out_wire_0_2(horizontal_tile_24_13_to_tile_24_14_2),
		.out_wire_0_3(horizontal_tile_24_13_to_tile_24_14_3),
		.in_wire_0_0(horizontal_tile_24_14_to_tile_24_13_0),
		.in_wire_0_1(horizontal_tile_24_14_to_tile_24_13_1),
		.in_wire_0_2(horizontal_tile_24_14_to_tile_24_13_2),
		.in_wire_0_3(horizontal_tile_24_14_to_tile_24_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(782)
	);

	pe_tile pe_tile_24_14(
		.out_wire_3_0(vertical_tile_24_14_to_tile_23_14_0),
		.out_wire_3_1(vertical_tile_24_14_to_tile_23_14_1),
		.out_wire_3_2(vertical_tile_24_14_to_tile_23_14_2),
		.out_wire_3_3(vertical_tile_24_14_to_tile_23_14_3),
		.in_wire_3_0(vertical_tile_23_14_to_tile_24_14_0),
		.in_wire_3_1(vertical_tile_23_14_to_tile_24_14_1),
		.in_wire_3_2(vertical_tile_23_14_to_tile_24_14_2),
		.in_wire_3_3(vertical_tile_23_14_to_tile_24_14_3),
		.out_wire_1_0(vertical_tile_24_14_to_tile_25_14_0),
		.out_wire_1_1(vertical_tile_24_14_to_tile_25_14_1),
		.out_wire_1_2(vertical_tile_24_14_to_tile_25_14_2),
		.out_wire_1_3(vertical_tile_24_14_to_tile_25_14_3),
		.in_wire_1_0(vertical_tile_25_14_to_tile_24_14_0),
		.in_wire_1_1(vertical_tile_25_14_to_tile_24_14_1),
		.in_wire_1_2(vertical_tile_25_14_to_tile_24_14_2),
		.in_wire_1_3(vertical_tile_25_14_to_tile_24_14_3),
		.out_wire_2_0(horizontal_tile_24_14_to_tile_24_13_0),
		.out_wire_2_1(horizontal_tile_24_14_to_tile_24_13_1),
		.out_wire_2_2(horizontal_tile_24_14_to_tile_24_13_2),
		.out_wire_2_3(horizontal_tile_24_14_to_tile_24_13_3),
		.in_wire_2_0(horizontal_tile_24_13_to_tile_24_14_0),
		.in_wire_2_1(horizontal_tile_24_13_to_tile_24_14_1),
		.in_wire_2_2(horizontal_tile_24_13_to_tile_24_14_2),
		.in_wire_2_3(horizontal_tile_24_13_to_tile_24_14_3),
		.out_wire_0_0(horizontal_tile_24_14_to_tile_24_15_0),
		.out_wire_0_1(horizontal_tile_24_14_to_tile_24_15_1),
		.out_wire_0_2(horizontal_tile_24_14_to_tile_24_15_2),
		.out_wire_0_3(horizontal_tile_24_14_to_tile_24_15_3),
		.in_wire_0_0(horizontal_tile_24_15_to_tile_24_14_0),
		.in_wire_0_1(horizontal_tile_24_15_to_tile_24_14_1),
		.in_wire_0_2(horizontal_tile_24_15_to_tile_24_14_2),
		.in_wire_0_3(horizontal_tile_24_15_to_tile_24_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(783)
	);

	pe_tile pe_tile_24_15(
		.out_wire_3_0(vertical_tile_24_15_to_tile_23_15_0),
		.out_wire_3_1(vertical_tile_24_15_to_tile_23_15_1),
		.out_wire_3_2(vertical_tile_24_15_to_tile_23_15_2),
		.out_wire_3_3(vertical_tile_24_15_to_tile_23_15_3),
		.in_wire_3_0(vertical_tile_23_15_to_tile_24_15_0),
		.in_wire_3_1(vertical_tile_23_15_to_tile_24_15_1),
		.in_wire_3_2(vertical_tile_23_15_to_tile_24_15_2),
		.in_wire_3_3(vertical_tile_23_15_to_tile_24_15_3),
		.out_wire_1_0(vertical_tile_24_15_to_tile_25_15_0),
		.out_wire_1_1(vertical_tile_24_15_to_tile_25_15_1),
		.out_wire_1_2(vertical_tile_24_15_to_tile_25_15_2),
		.out_wire_1_3(vertical_tile_24_15_to_tile_25_15_3),
		.in_wire_1_0(vertical_tile_25_15_to_tile_24_15_0),
		.in_wire_1_1(vertical_tile_25_15_to_tile_24_15_1),
		.in_wire_1_2(vertical_tile_25_15_to_tile_24_15_2),
		.in_wire_1_3(vertical_tile_25_15_to_tile_24_15_3),
		.out_wire_2_0(horizontal_tile_24_15_to_tile_24_14_0),
		.out_wire_2_1(horizontal_tile_24_15_to_tile_24_14_1),
		.out_wire_2_2(horizontal_tile_24_15_to_tile_24_14_2),
		.out_wire_2_3(horizontal_tile_24_15_to_tile_24_14_3),
		.in_wire_2_0(horizontal_tile_24_14_to_tile_24_15_0),
		.in_wire_2_1(horizontal_tile_24_14_to_tile_24_15_1),
		.in_wire_2_2(horizontal_tile_24_14_to_tile_24_15_2),
		.in_wire_2_3(horizontal_tile_24_14_to_tile_24_15_3),
		.out_wire_0_0(horizontal_tile_24_15_to_tile_24_16_0),
		.out_wire_0_1(horizontal_tile_24_15_to_tile_24_16_1),
		.out_wire_0_2(horizontal_tile_24_15_to_tile_24_16_2),
		.out_wire_0_3(horizontal_tile_24_15_to_tile_24_16_3),
		.in_wire_0_0(horizontal_tile_24_16_to_tile_24_15_0),
		.in_wire_0_1(horizontal_tile_24_16_to_tile_24_15_1),
		.in_wire_0_2(horizontal_tile_24_16_to_tile_24_15_2),
		.in_wire_0_3(horizontal_tile_24_16_to_tile_24_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(784)
	);

	pe_tile pe_tile_24_16(
		.out_wire_3_0(vertical_tile_24_16_to_tile_23_16_0),
		.out_wire_3_1(vertical_tile_24_16_to_tile_23_16_1),
		.out_wire_3_2(vertical_tile_24_16_to_tile_23_16_2),
		.out_wire_3_3(vertical_tile_24_16_to_tile_23_16_3),
		.in_wire_3_0(vertical_tile_23_16_to_tile_24_16_0),
		.in_wire_3_1(vertical_tile_23_16_to_tile_24_16_1),
		.in_wire_3_2(vertical_tile_23_16_to_tile_24_16_2),
		.in_wire_3_3(vertical_tile_23_16_to_tile_24_16_3),
		.out_wire_1_0(vertical_tile_24_16_to_tile_25_16_0),
		.out_wire_1_1(vertical_tile_24_16_to_tile_25_16_1),
		.out_wire_1_2(vertical_tile_24_16_to_tile_25_16_2),
		.out_wire_1_3(vertical_tile_24_16_to_tile_25_16_3),
		.in_wire_1_0(vertical_tile_25_16_to_tile_24_16_0),
		.in_wire_1_1(vertical_tile_25_16_to_tile_24_16_1),
		.in_wire_1_2(vertical_tile_25_16_to_tile_24_16_2),
		.in_wire_1_3(vertical_tile_25_16_to_tile_24_16_3),
		.out_wire_2_0(horizontal_tile_24_16_to_tile_24_15_0),
		.out_wire_2_1(horizontal_tile_24_16_to_tile_24_15_1),
		.out_wire_2_2(horizontal_tile_24_16_to_tile_24_15_2),
		.out_wire_2_3(horizontal_tile_24_16_to_tile_24_15_3),
		.in_wire_2_0(horizontal_tile_24_15_to_tile_24_16_0),
		.in_wire_2_1(horizontal_tile_24_15_to_tile_24_16_1),
		.in_wire_2_2(horizontal_tile_24_15_to_tile_24_16_2),
		.in_wire_2_3(horizontal_tile_24_15_to_tile_24_16_3),
		.out_wire_0_0(horizontal_tile_24_16_to_tile_24_17_0),
		.out_wire_0_1(horizontal_tile_24_16_to_tile_24_17_1),
		.out_wire_0_2(horizontal_tile_24_16_to_tile_24_17_2),
		.out_wire_0_3(horizontal_tile_24_16_to_tile_24_17_3),
		.in_wire_0_0(horizontal_tile_24_17_to_tile_24_16_0),
		.in_wire_0_1(horizontal_tile_24_17_to_tile_24_16_1),
		.in_wire_0_2(horizontal_tile_24_17_to_tile_24_16_2),
		.in_wire_0_3(horizontal_tile_24_17_to_tile_24_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(785)
	);

	pe_tile pe_tile_24_17(
		.out_wire_3_0(vertical_tile_24_17_to_tile_23_17_0),
		.out_wire_3_1(vertical_tile_24_17_to_tile_23_17_1),
		.out_wire_3_2(vertical_tile_24_17_to_tile_23_17_2),
		.out_wire_3_3(vertical_tile_24_17_to_tile_23_17_3),
		.in_wire_3_0(vertical_tile_23_17_to_tile_24_17_0),
		.in_wire_3_1(vertical_tile_23_17_to_tile_24_17_1),
		.in_wire_3_2(vertical_tile_23_17_to_tile_24_17_2),
		.in_wire_3_3(vertical_tile_23_17_to_tile_24_17_3),
		.out_wire_1_0(vertical_tile_24_17_to_tile_25_17_0),
		.out_wire_1_1(vertical_tile_24_17_to_tile_25_17_1),
		.out_wire_1_2(vertical_tile_24_17_to_tile_25_17_2),
		.out_wire_1_3(vertical_tile_24_17_to_tile_25_17_3),
		.in_wire_1_0(vertical_tile_25_17_to_tile_24_17_0),
		.in_wire_1_1(vertical_tile_25_17_to_tile_24_17_1),
		.in_wire_1_2(vertical_tile_25_17_to_tile_24_17_2),
		.in_wire_1_3(vertical_tile_25_17_to_tile_24_17_3),
		.out_wire_2_0(horizontal_tile_24_17_to_tile_24_16_0),
		.out_wire_2_1(horizontal_tile_24_17_to_tile_24_16_1),
		.out_wire_2_2(horizontal_tile_24_17_to_tile_24_16_2),
		.out_wire_2_3(horizontal_tile_24_17_to_tile_24_16_3),
		.in_wire_2_0(horizontal_tile_24_16_to_tile_24_17_0),
		.in_wire_2_1(horizontal_tile_24_16_to_tile_24_17_1),
		.in_wire_2_2(horizontal_tile_24_16_to_tile_24_17_2),
		.in_wire_2_3(horizontal_tile_24_16_to_tile_24_17_3),
		.out_wire_0_0(horizontal_tile_24_17_to_tile_24_18_0),
		.out_wire_0_1(horizontal_tile_24_17_to_tile_24_18_1),
		.out_wire_0_2(horizontal_tile_24_17_to_tile_24_18_2),
		.out_wire_0_3(horizontal_tile_24_17_to_tile_24_18_3),
		.in_wire_0_0(horizontal_tile_24_18_to_tile_24_17_0),
		.in_wire_0_1(horizontal_tile_24_18_to_tile_24_17_1),
		.in_wire_0_2(horizontal_tile_24_18_to_tile_24_17_2),
		.in_wire_0_3(horizontal_tile_24_18_to_tile_24_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(786)
	);

	pe_tile pe_tile_24_18(
		.out_wire_3_0(vertical_tile_24_18_to_tile_23_18_0),
		.out_wire_3_1(vertical_tile_24_18_to_tile_23_18_1),
		.out_wire_3_2(vertical_tile_24_18_to_tile_23_18_2),
		.out_wire_3_3(vertical_tile_24_18_to_tile_23_18_3),
		.in_wire_3_0(vertical_tile_23_18_to_tile_24_18_0),
		.in_wire_3_1(vertical_tile_23_18_to_tile_24_18_1),
		.in_wire_3_2(vertical_tile_23_18_to_tile_24_18_2),
		.in_wire_3_3(vertical_tile_23_18_to_tile_24_18_3),
		.out_wire_1_0(vertical_tile_24_18_to_tile_25_18_0),
		.out_wire_1_1(vertical_tile_24_18_to_tile_25_18_1),
		.out_wire_1_2(vertical_tile_24_18_to_tile_25_18_2),
		.out_wire_1_3(vertical_tile_24_18_to_tile_25_18_3),
		.in_wire_1_0(vertical_tile_25_18_to_tile_24_18_0),
		.in_wire_1_1(vertical_tile_25_18_to_tile_24_18_1),
		.in_wire_1_2(vertical_tile_25_18_to_tile_24_18_2),
		.in_wire_1_3(vertical_tile_25_18_to_tile_24_18_3),
		.out_wire_2_0(horizontal_tile_24_18_to_tile_24_17_0),
		.out_wire_2_1(horizontal_tile_24_18_to_tile_24_17_1),
		.out_wire_2_2(horizontal_tile_24_18_to_tile_24_17_2),
		.out_wire_2_3(horizontal_tile_24_18_to_tile_24_17_3),
		.in_wire_2_0(horizontal_tile_24_17_to_tile_24_18_0),
		.in_wire_2_1(horizontal_tile_24_17_to_tile_24_18_1),
		.in_wire_2_2(horizontal_tile_24_17_to_tile_24_18_2),
		.in_wire_2_3(horizontal_tile_24_17_to_tile_24_18_3),
		.out_wire_0_0(horizontal_tile_24_18_to_tile_24_19_0),
		.out_wire_0_1(horizontal_tile_24_18_to_tile_24_19_1),
		.out_wire_0_2(horizontal_tile_24_18_to_tile_24_19_2),
		.out_wire_0_3(horizontal_tile_24_18_to_tile_24_19_3),
		.in_wire_0_0(horizontal_tile_24_19_to_tile_24_18_0),
		.in_wire_0_1(horizontal_tile_24_19_to_tile_24_18_1),
		.in_wire_0_2(horizontal_tile_24_19_to_tile_24_18_2),
		.in_wire_0_3(horizontal_tile_24_19_to_tile_24_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(787)
	);

	pe_tile pe_tile_24_19(
		.out_wire_3_0(vertical_tile_24_19_to_tile_23_19_0),
		.out_wire_3_1(vertical_tile_24_19_to_tile_23_19_1),
		.out_wire_3_2(vertical_tile_24_19_to_tile_23_19_2),
		.out_wire_3_3(vertical_tile_24_19_to_tile_23_19_3),
		.in_wire_3_0(vertical_tile_23_19_to_tile_24_19_0),
		.in_wire_3_1(vertical_tile_23_19_to_tile_24_19_1),
		.in_wire_3_2(vertical_tile_23_19_to_tile_24_19_2),
		.in_wire_3_3(vertical_tile_23_19_to_tile_24_19_3),
		.out_wire_1_0(vertical_tile_24_19_to_tile_25_19_0),
		.out_wire_1_1(vertical_tile_24_19_to_tile_25_19_1),
		.out_wire_1_2(vertical_tile_24_19_to_tile_25_19_2),
		.out_wire_1_3(vertical_tile_24_19_to_tile_25_19_3),
		.in_wire_1_0(vertical_tile_25_19_to_tile_24_19_0),
		.in_wire_1_1(vertical_tile_25_19_to_tile_24_19_1),
		.in_wire_1_2(vertical_tile_25_19_to_tile_24_19_2),
		.in_wire_1_3(vertical_tile_25_19_to_tile_24_19_3),
		.out_wire_2_0(horizontal_tile_24_19_to_tile_24_18_0),
		.out_wire_2_1(horizontal_tile_24_19_to_tile_24_18_1),
		.out_wire_2_2(horizontal_tile_24_19_to_tile_24_18_2),
		.out_wire_2_3(horizontal_tile_24_19_to_tile_24_18_3),
		.in_wire_2_0(horizontal_tile_24_18_to_tile_24_19_0),
		.in_wire_2_1(horizontal_tile_24_18_to_tile_24_19_1),
		.in_wire_2_2(horizontal_tile_24_18_to_tile_24_19_2),
		.in_wire_2_3(horizontal_tile_24_18_to_tile_24_19_3),
		.out_wire_0_0(horizontal_tile_24_19_to_tile_24_20_0),
		.out_wire_0_1(horizontal_tile_24_19_to_tile_24_20_1),
		.out_wire_0_2(horizontal_tile_24_19_to_tile_24_20_2),
		.out_wire_0_3(horizontal_tile_24_19_to_tile_24_20_3),
		.in_wire_0_0(horizontal_tile_24_20_to_tile_24_19_0),
		.in_wire_0_1(horizontal_tile_24_20_to_tile_24_19_1),
		.in_wire_0_2(horizontal_tile_24_20_to_tile_24_19_2),
		.in_wire_0_3(horizontal_tile_24_20_to_tile_24_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(788)
	);

	pe_tile pe_tile_24_20(
		.out_wire_3_0(vertical_tile_24_20_to_tile_23_20_0),
		.out_wire_3_1(vertical_tile_24_20_to_tile_23_20_1),
		.out_wire_3_2(vertical_tile_24_20_to_tile_23_20_2),
		.out_wire_3_3(vertical_tile_24_20_to_tile_23_20_3),
		.in_wire_3_0(vertical_tile_23_20_to_tile_24_20_0),
		.in_wire_3_1(vertical_tile_23_20_to_tile_24_20_1),
		.in_wire_3_2(vertical_tile_23_20_to_tile_24_20_2),
		.in_wire_3_3(vertical_tile_23_20_to_tile_24_20_3),
		.out_wire_1_0(vertical_tile_24_20_to_tile_25_20_0),
		.out_wire_1_1(vertical_tile_24_20_to_tile_25_20_1),
		.out_wire_1_2(vertical_tile_24_20_to_tile_25_20_2),
		.out_wire_1_3(vertical_tile_24_20_to_tile_25_20_3),
		.in_wire_1_0(vertical_tile_25_20_to_tile_24_20_0),
		.in_wire_1_1(vertical_tile_25_20_to_tile_24_20_1),
		.in_wire_1_2(vertical_tile_25_20_to_tile_24_20_2),
		.in_wire_1_3(vertical_tile_25_20_to_tile_24_20_3),
		.out_wire_2_0(horizontal_tile_24_20_to_tile_24_19_0),
		.out_wire_2_1(horizontal_tile_24_20_to_tile_24_19_1),
		.out_wire_2_2(horizontal_tile_24_20_to_tile_24_19_2),
		.out_wire_2_3(horizontal_tile_24_20_to_tile_24_19_3),
		.in_wire_2_0(horizontal_tile_24_19_to_tile_24_20_0),
		.in_wire_2_1(horizontal_tile_24_19_to_tile_24_20_1),
		.in_wire_2_2(horizontal_tile_24_19_to_tile_24_20_2),
		.in_wire_2_3(horizontal_tile_24_19_to_tile_24_20_3),
		.out_wire_0_0(horizontal_tile_24_20_to_tile_24_21_0),
		.out_wire_0_1(horizontal_tile_24_20_to_tile_24_21_1),
		.out_wire_0_2(horizontal_tile_24_20_to_tile_24_21_2),
		.out_wire_0_3(horizontal_tile_24_20_to_tile_24_21_3),
		.in_wire_0_0(horizontal_tile_24_21_to_tile_24_20_0),
		.in_wire_0_1(horizontal_tile_24_21_to_tile_24_20_1),
		.in_wire_0_2(horizontal_tile_24_21_to_tile_24_20_2),
		.in_wire_0_3(horizontal_tile_24_21_to_tile_24_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(789)
	);

	pe_tile pe_tile_24_21(
		.out_wire_3_0(vertical_tile_24_21_to_tile_23_21_0),
		.out_wire_3_1(vertical_tile_24_21_to_tile_23_21_1),
		.out_wire_3_2(vertical_tile_24_21_to_tile_23_21_2),
		.out_wire_3_3(vertical_tile_24_21_to_tile_23_21_3),
		.in_wire_3_0(vertical_tile_23_21_to_tile_24_21_0),
		.in_wire_3_1(vertical_tile_23_21_to_tile_24_21_1),
		.in_wire_3_2(vertical_tile_23_21_to_tile_24_21_2),
		.in_wire_3_3(vertical_tile_23_21_to_tile_24_21_3),
		.out_wire_1_0(vertical_tile_24_21_to_tile_25_21_0),
		.out_wire_1_1(vertical_tile_24_21_to_tile_25_21_1),
		.out_wire_1_2(vertical_tile_24_21_to_tile_25_21_2),
		.out_wire_1_3(vertical_tile_24_21_to_tile_25_21_3),
		.in_wire_1_0(vertical_tile_25_21_to_tile_24_21_0),
		.in_wire_1_1(vertical_tile_25_21_to_tile_24_21_1),
		.in_wire_1_2(vertical_tile_25_21_to_tile_24_21_2),
		.in_wire_1_3(vertical_tile_25_21_to_tile_24_21_3),
		.out_wire_2_0(horizontal_tile_24_21_to_tile_24_20_0),
		.out_wire_2_1(horizontal_tile_24_21_to_tile_24_20_1),
		.out_wire_2_2(horizontal_tile_24_21_to_tile_24_20_2),
		.out_wire_2_3(horizontal_tile_24_21_to_tile_24_20_3),
		.in_wire_2_0(horizontal_tile_24_20_to_tile_24_21_0),
		.in_wire_2_1(horizontal_tile_24_20_to_tile_24_21_1),
		.in_wire_2_2(horizontal_tile_24_20_to_tile_24_21_2),
		.in_wire_2_3(horizontal_tile_24_20_to_tile_24_21_3),
		.out_wire_0_0(horizontal_tile_24_21_to_tile_24_22_0),
		.out_wire_0_1(horizontal_tile_24_21_to_tile_24_22_1),
		.out_wire_0_2(horizontal_tile_24_21_to_tile_24_22_2),
		.out_wire_0_3(horizontal_tile_24_21_to_tile_24_22_3),
		.in_wire_0_0(horizontal_tile_24_22_to_tile_24_21_0),
		.in_wire_0_1(horizontal_tile_24_22_to_tile_24_21_1),
		.in_wire_0_2(horizontal_tile_24_22_to_tile_24_21_2),
		.in_wire_0_3(horizontal_tile_24_22_to_tile_24_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(790)
	);

	pe_tile pe_tile_24_22(
		.out_wire_3_0(vertical_tile_24_22_to_tile_23_22_0),
		.out_wire_3_1(vertical_tile_24_22_to_tile_23_22_1),
		.out_wire_3_2(vertical_tile_24_22_to_tile_23_22_2),
		.out_wire_3_3(vertical_tile_24_22_to_tile_23_22_3),
		.in_wire_3_0(vertical_tile_23_22_to_tile_24_22_0),
		.in_wire_3_1(vertical_tile_23_22_to_tile_24_22_1),
		.in_wire_3_2(vertical_tile_23_22_to_tile_24_22_2),
		.in_wire_3_3(vertical_tile_23_22_to_tile_24_22_3),
		.out_wire_1_0(vertical_tile_24_22_to_tile_25_22_0),
		.out_wire_1_1(vertical_tile_24_22_to_tile_25_22_1),
		.out_wire_1_2(vertical_tile_24_22_to_tile_25_22_2),
		.out_wire_1_3(vertical_tile_24_22_to_tile_25_22_3),
		.in_wire_1_0(vertical_tile_25_22_to_tile_24_22_0),
		.in_wire_1_1(vertical_tile_25_22_to_tile_24_22_1),
		.in_wire_1_2(vertical_tile_25_22_to_tile_24_22_2),
		.in_wire_1_3(vertical_tile_25_22_to_tile_24_22_3),
		.out_wire_2_0(horizontal_tile_24_22_to_tile_24_21_0),
		.out_wire_2_1(horizontal_tile_24_22_to_tile_24_21_1),
		.out_wire_2_2(horizontal_tile_24_22_to_tile_24_21_2),
		.out_wire_2_3(horizontal_tile_24_22_to_tile_24_21_3),
		.in_wire_2_0(horizontal_tile_24_21_to_tile_24_22_0),
		.in_wire_2_1(horizontal_tile_24_21_to_tile_24_22_1),
		.in_wire_2_2(horizontal_tile_24_21_to_tile_24_22_2),
		.in_wire_2_3(horizontal_tile_24_21_to_tile_24_22_3),
		.out_wire_0_0(horizontal_tile_24_22_to_tile_24_23_0),
		.out_wire_0_1(horizontal_tile_24_22_to_tile_24_23_1),
		.out_wire_0_2(horizontal_tile_24_22_to_tile_24_23_2),
		.out_wire_0_3(horizontal_tile_24_22_to_tile_24_23_3),
		.in_wire_0_0(horizontal_tile_24_23_to_tile_24_22_0),
		.in_wire_0_1(horizontal_tile_24_23_to_tile_24_22_1),
		.in_wire_0_2(horizontal_tile_24_23_to_tile_24_22_2),
		.in_wire_0_3(horizontal_tile_24_23_to_tile_24_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(791)
	);

	pe_tile pe_tile_24_23(
		.out_wire_3_0(vertical_tile_24_23_to_tile_23_23_0),
		.out_wire_3_1(vertical_tile_24_23_to_tile_23_23_1),
		.out_wire_3_2(vertical_tile_24_23_to_tile_23_23_2),
		.out_wire_3_3(vertical_tile_24_23_to_tile_23_23_3),
		.in_wire_3_0(vertical_tile_23_23_to_tile_24_23_0),
		.in_wire_3_1(vertical_tile_23_23_to_tile_24_23_1),
		.in_wire_3_2(vertical_tile_23_23_to_tile_24_23_2),
		.in_wire_3_3(vertical_tile_23_23_to_tile_24_23_3),
		.out_wire_1_0(vertical_tile_24_23_to_tile_25_23_0),
		.out_wire_1_1(vertical_tile_24_23_to_tile_25_23_1),
		.out_wire_1_2(vertical_tile_24_23_to_tile_25_23_2),
		.out_wire_1_3(vertical_tile_24_23_to_tile_25_23_3),
		.in_wire_1_0(vertical_tile_25_23_to_tile_24_23_0),
		.in_wire_1_1(vertical_tile_25_23_to_tile_24_23_1),
		.in_wire_1_2(vertical_tile_25_23_to_tile_24_23_2),
		.in_wire_1_3(vertical_tile_25_23_to_tile_24_23_3),
		.out_wire_2_0(horizontal_tile_24_23_to_tile_24_22_0),
		.out_wire_2_1(horizontal_tile_24_23_to_tile_24_22_1),
		.out_wire_2_2(horizontal_tile_24_23_to_tile_24_22_2),
		.out_wire_2_3(horizontal_tile_24_23_to_tile_24_22_3),
		.in_wire_2_0(horizontal_tile_24_22_to_tile_24_23_0),
		.in_wire_2_1(horizontal_tile_24_22_to_tile_24_23_1),
		.in_wire_2_2(horizontal_tile_24_22_to_tile_24_23_2),
		.in_wire_2_3(horizontal_tile_24_22_to_tile_24_23_3),
		.out_wire_0_0(horizontal_tile_24_23_to_tile_24_24_0),
		.out_wire_0_1(horizontal_tile_24_23_to_tile_24_24_1),
		.out_wire_0_2(horizontal_tile_24_23_to_tile_24_24_2),
		.out_wire_0_3(horizontal_tile_24_23_to_tile_24_24_3),
		.in_wire_0_0(horizontal_tile_24_24_to_tile_24_23_0),
		.in_wire_0_1(horizontal_tile_24_24_to_tile_24_23_1),
		.in_wire_0_2(horizontal_tile_24_24_to_tile_24_23_2),
		.in_wire_0_3(horizontal_tile_24_24_to_tile_24_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(792)
	);

	pe_tile pe_tile_24_24(
		.out_wire_3_0(vertical_tile_24_24_to_tile_23_24_0),
		.out_wire_3_1(vertical_tile_24_24_to_tile_23_24_1),
		.out_wire_3_2(vertical_tile_24_24_to_tile_23_24_2),
		.out_wire_3_3(vertical_tile_24_24_to_tile_23_24_3),
		.in_wire_3_0(vertical_tile_23_24_to_tile_24_24_0),
		.in_wire_3_1(vertical_tile_23_24_to_tile_24_24_1),
		.in_wire_3_2(vertical_tile_23_24_to_tile_24_24_2),
		.in_wire_3_3(vertical_tile_23_24_to_tile_24_24_3),
		.out_wire_1_0(vertical_tile_24_24_to_tile_25_24_0),
		.out_wire_1_1(vertical_tile_24_24_to_tile_25_24_1),
		.out_wire_1_2(vertical_tile_24_24_to_tile_25_24_2),
		.out_wire_1_3(vertical_tile_24_24_to_tile_25_24_3),
		.in_wire_1_0(vertical_tile_25_24_to_tile_24_24_0),
		.in_wire_1_1(vertical_tile_25_24_to_tile_24_24_1),
		.in_wire_1_2(vertical_tile_25_24_to_tile_24_24_2),
		.in_wire_1_3(vertical_tile_25_24_to_tile_24_24_3),
		.out_wire_2_0(horizontal_tile_24_24_to_tile_24_23_0),
		.out_wire_2_1(horizontal_tile_24_24_to_tile_24_23_1),
		.out_wire_2_2(horizontal_tile_24_24_to_tile_24_23_2),
		.out_wire_2_3(horizontal_tile_24_24_to_tile_24_23_3),
		.in_wire_2_0(horizontal_tile_24_23_to_tile_24_24_0),
		.in_wire_2_1(horizontal_tile_24_23_to_tile_24_24_1),
		.in_wire_2_2(horizontal_tile_24_23_to_tile_24_24_2),
		.in_wire_2_3(horizontal_tile_24_23_to_tile_24_24_3),
		.out_wire_0_0(horizontal_tile_24_24_to_tile_24_25_0),
		.out_wire_0_1(horizontal_tile_24_24_to_tile_24_25_1),
		.out_wire_0_2(horizontal_tile_24_24_to_tile_24_25_2),
		.out_wire_0_3(horizontal_tile_24_24_to_tile_24_25_3),
		.in_wire_0_0(horizontal_tile_24_25_to_tile_24_24_0),
		.in_wire_0_1(horizontal_tile_24_25_to_tile_24_24_1),
		.in_wire_0_2(horizontal_tile_24_25_to_tile_24_24_2),
		.in_wire_0_3(horizontal_tile_24_25_to_tile_24_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(793)
	);

	pe_tile pe_tile_24_25(
		.out_wire_3_0(vertical_tile_24_25_to_tile_23_25_0),
		.out_wire_3_1(vertical_tile_24_25_to_tile_23_25_1),
		.out_wire_3_2(vertical_tile_24_25_to_tile_23_25_2),
		.out_wire_3_3(vertical_tile_24_25_to_tile_23_25_3),
		.in_wire_3_0(vertical_tile_23_25_to_tile_24_25_0),
		.in_wire_3_1(vertical_tile_23_25_to_tile_24_25_1),
		.in_wire_3_2(vertical_tile_23_25_to_tile_24_25_2),
		.in_wire_3_3(vertical_tile_23_25_to_tile_24_25_3),
		.out_wire_1_0(vertical_tile_24_25_to_tile_25_25_0),
		.out_wire_1_1(vertical_tile_24_25_to_tile_25_25_1),
		.out_wire_1_2(vertical_tile_24_25_to_tile_25_25_2),
		.out_wire_1_3(vertical_tile_24_25_to_tile_25_25_3),
		.in_wire_1_0(vertical_tile_25_25_to_tile_24_25_0),
		.in_wire_1_1(vertical_tile_25_25_to_tile_24_25_1),
		.in_wire_1_2(vertical_tile_25_25_to_tile_24_25_2),
		.in_wire_1_3(vertical_tile_25_25_to_tile_24_25_3),
		.out_wire_2_0(horizontal_tile_24_25_to_tile_24_24_0),
		.out_wire_2_1(horizontal_tile_24_25_to_tile_24_24_1),
		.out_wire_2_2(horizontal_tile_24_25_to_tile_24_24_2),
		.out_wire_2_3(horizontal_tile_24_25_to_tile_24_24_3),
		.in_wire_2_0(horizontal_tile_24_24_to_tile_24_25_0),
		.in_wire_2_1(horizontal_tile_24_24_to_tile_24_25_1),
		.in_wire_2_2(horizontal_tile_24_24_to_tile_24_25_2),
		.in_wire_2_3(horizontal_tile_24_24_to_tile_24_25_3),
		.out_wire_0_0(horizontal_tile_24_25_to_tile_24_26_0),
		.out_wire_0_1(horizontal_tile_24_25_to_tile_24_26_1),
		.out_wire_0_2(horizontal_tile_24_25_to_tile_24_26_2),
		.out_wire_0_3(horizontal_tile_24_25_to_tile_24_26_3),
		.in_wire_0_0(horizontal_tile_24_26_to_tile_24_25_0),
		.in_wire_0_1(horizontal_tile_24_26_to_tile_24_25_1),
		.in_wire_0_2(horizontal_tile_24_26_to_tile_24_25_2),
		.in_wire_0_3(horizontal_tile_24_26_to_tile_24_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(794)
	);

	pe_tile pe_tile_24_26(
		.out_wire_3_0(vertical_tile_24_26_to_tile_23_26_0),
		.out_wire_3_1(vertical_tile_24_26_to_tile_23_26_1),
		.out_wire_3_2(vertical_tile_24_26_to_tile_23_26_2),
		.out_wire_3_3(vertical_tile_24_26_to_tile_23_26_3),
		.in_wire_3_0(vertical_tile_23_26_to_tile_24_26_0),
		.in_wire_3_1(vertical_tile_23_26_to_tile_24_26_1),
		.in_wire_3_2(vertical_tile_23_26_to_tile_24_26_2),
		.in_wire_3_3(vertical_tile_23_26_to_tile_24_26_3),
		.out_wire_1_0(vertical_tile_24_26_to_tile_25_26_0),
		.out_wire_1_1(vertical_tile_24_26_to_tile_25_26_1),
		.out_wire_1_2(vertical_tile_24_26_to_tile_25_26_2),
		.out_wire_1_3(vertical_tile_24_26_to_tile_25_26_3),
		.in_wire_1_0(vertical_tile_25_26_to_tile_24_26_0),
		.in_wire_1_1(vertical_tile_25_26_to_tile_24_26_1),
		.in_wire_1_2(vertical_tile_25_26_to_tile_24_26_2),
		.in_wire_1_3(vertical_tile_25_26_to_tile_24_26_3),
		.out_wire_2_0(horizontal_tile_24_26_to_tile_24_25_0),
		.out_wire_2_1(horizontal_tile_24_26_to_tile_24_25_1),
		.out_wire_2_2(horizontal_tile_24_26_to_tile_24_25_2),
		.out_wire_2_3(horizontal_tile_24_26_to_tile_24_25_3),
		.in_wire_2_0(horizontal_tile_24_25_to_tile_24_26_0),
		.in_wire_2_1(horizontal_tile_24_25_to_tile_24_26_1),
		.in_wire_2_2(horizontal_tile_24_25_to_tile_24_26_2),
		.in_wire_2_3(horizontal_tile_24_25_to_tile_24_26_3),
		.out_wire_0_0(horizontal_tile_24_26_to_tile_24_27_0),
		.out_wire_0_1(horizontal_tile_24_26_to_tile_24_27_1),
		.out_wire_0_2(horizontal_tile_24_26_to_tile_24_27_2),
		.out_wire_0_3(horizontal_tile_24_26_to_tile_24_27_3),
		.in_wire_0_0(horizontal_tile_24_27_to_tile_24_26_0),
		.in_wire_0_1(horizontal_tile_24_27_to_tile_24_26_1),
		.in_wire_0_2(horizontal_tile_24_27_to_tile_24_26_2),
		.in_wire_0_3(horizontal_tile_24_27_to_tile_24_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(795)
	);

	pe_tile pe_tile_24_27(
		.out_wire_3_0(vertical_tile_24_27_to_tile_23_27_0),
		.out_wire_3_1(vertical_tile_24_27_to_tile_23_27_1),
		.out_wire_3_2(vertical_tile_24_27_to_tile_23_27_2),
		.out_wire_3_3(vertical_tile_24_27_to_tile_23_27_3),
		.in_wire_3_0(vertical_tile_23_27_to_tile_24_27_0),
		.in_wire_3_1(vertical_tile_23_27_to_tile_24_27_1),
		.in_wire_3_2(vertical_tile_23_27_to_tile_24_27_2),
		.in_wire_3_3(vertical_tile_23_27_to_tile_24_27_3),
		.out_wire_1_0(vertical_tile_24_27_to_tile_25_27_0),
		.out_wire_1_1(vertical_tile_24_27_to_tile_25_27_1),
		.out_wire_1_2(vertical_tile_24_27_to_tile_25_27_2),
		.out_wire_1_3(vertical_tile_24_27_to_tile_25_27_3),
		.in_wire_1_0(vertical_tile_25_27_to_tile_24_27_0),
		.in_wire_1_1(vertical_tile_25_27_to_tile_24_27_1),
		.in_wire_1_2(vertical_tile_25_27_to_tile_24_27_2),
		.in_wire_1_3(vertical_tile_25_27_to_tile_24_27_3),
		.out_wire_2_0(horizontal_tile_24_27_to_tile_24_26_0),
		.out_wire_2_1(horizontal_tile_24_27_to_tile_24_26_1),
		.out_wire_2_2(horizontal_tile_24_27_to_tile_24_26_2),
		.out_wire_2_3(horizontal_tile_24_27_to_tile_24_26_3),
		.in_wire_2_0(horizontal_tile_24_26_to_tile_24_27_0),
		.in_wire_2_1(horizontal_tile_24_26_to_tile_24_27_1),
		.in_wire_2_2(horizontal_tile_24_26_to_tile_24_27_2),
		.in_wire_2_3(horizontal_tile_24_26_to_tile_24_27_3),
		.out_wire_0_0(horizontal_tile_24_27_to_tile_24_28_0),
		.out_wire_0_1(horizontal_tile_24_27_to_tile_24_28_1),
		.out_wire_0_2(horizontal_tile_24_27_to_tile_24_28_2),
		.out_wire_0_3(horizontal_tile_24_27_to_tile_24_28_3),
		.in_wire_0_0(horizontal_tile_24_28_to_tile_24_27_0),
		.in_wire_0_1(horizontal_tile_24_28_to_tile_24_27_1),
		.in_wire_0_2(horizontal_tile_24_28_to_tile_24_27_2),
		.in_wire_0_3(horizontal_tile_24_28_to_tile_24_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(796)
	);

	pe_tile pe_tile_24_28(
		.out_wire_3_0(vertical_tile_24_28_to_tile_23_28_0),
		.out_wire_3_1(vertical_tile_24_28_to_tile_23_28_1),
		.out_wire_3_2(vertical_tile_24_28_to_tile_23_28_2),
		.out_wire_3_3(vertical_tile_24_28_to_tile_23_28_3),
		.in_wire_3_0(vertical_tile_23_28_to_tile_24_28_0),
		.in_wire_3_1(vertical_tile_23_28_to_tile_24_28_1),
		.in_wire_3_2(vertical_tile_23_28_to_tile_24_28_2),
		.in_wire_3_3(vertical_tile_23_28_to_tile_24_28_3),
		.out_wire_1_0(vertical_tile_24_28_to_tile_25_28_0),
		.out_wire_1_1(vertical_tile_24_28_to_tile_25_28_1),
		.out_wire_1_2(vertical_tile_24_28_to_tile_25_28_2),
		.out_wire_1_3(vertical_tile_24_28_to_tile_25_28_3),
		.in_wire_1_0(vertical_tile_25_28_to_tile_24_28_0),
		.in_wire_1_1(vertical_tile_25_28_to_tile_24_28_1),
		.in_wire_1_2(vertical_tile_25_28_to_tile_24_28_2),
		.in_wire_1_3(vertical_tile_25_28_to_tile_24_28_3),
		.out_wire_2_0(horizontal_tile_24_28_to_tile_24_27_0),
		.out_wire_2_1(horizontal_tile_24_28_to_tile_24_27_1),
		.out_wire_2_2(horizontal_tile_24_28_to_tile_24_27_2),
		.out_wire_2_3(horizontal_tile_24_28_to_tile_24_27_3),
		.in_wire_2_0(horizontal_tile_24_27_to_tile_24_28_0),
		.in_wire_2_1(horizontal_tile_24_27_to_tile_24_28_1),
		.in_wire_2_2(horizontal_tile_24_27_to_tile_24_28_2),
		.in_wire_2_3(horizontal_tile_24_27_to_tile_24_28_3),
		.out_wire_0_0(horizontal_tile_24_28_to_tile_24_29_0),
		.out_wire_0_1(horizontal_tile_24_28_to_tile_24_29_1),
		.out_wire_0_2(horizontal_tile_24_28_to_tile_24_29_2),
		.out_wire_0_3(horizontal_tile_24_28_to_tile_24_29_3),
		.in_wire_0_0(horizontal_tile_24_29_to_tile_24_28_0),
		.in_wire_0_1(horizontal_tile_24_29_to_tile_24_28_1),
		.in_wire_0_2(horizontal_tile_24_29_to_tile_24_28_2),
		.in_wire_0_3(horizontal_tile_24_29_to_tile_24_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(797)
	);

	pe_tile pe_tile_24_29(
		.out_wire_3_0(vertical_tile_24_29_to_tile_23_29_0),
		.out_wire_3_1(vertical_tile_24_29_to_tile_23_29_1),
		.out_wire_3_2(vertical_tile_24_29_to_tile_23_29_2),
		.out_wire_3_3(vertical_tile_24_29_to_tile_23_29_3),
		.in_wire_3_0(vertical_tile_23_29_to_tile_24_29_0),
		.in_wire_3_1(vertical_tile_23_29_to_tile_24_29_1),
		.in_wire_3_2(vertical_tile_23_29_to_tile_24_29_2),
		.in_wire_3_3(vertical_tile_23_29_to_tile_24_29_3),
		.out_wire_1_0(vertical_tile_24_29_to_tile_25_29_0),
		.out_wire_1_1(vertical_tile_24_29_to_tile_25_29_1),
		.out_wire_1_2(vertical_tile_24_29_to_tile_25_29_2),
		.out_wire_1_3(vertical_tile_24_29_to_tile_25_29_3),
		.in_wire_1_0(vertical_tile_25_29_to_tile_24_29_0),
		.in_wire_1_1(vertical_tile_25_29_to_tile_24_29_1),
		.in_wire_1_2(vertical_tile_25_29_to_tile_24_29_2),
		.in_wire_1_3(vertical_tile_25_29_to_tile_24_29_3),
		.out_wire_2_0(horizontal_tile_24_29_to_tile_24_28_0),
		.out_wire_2_1(horizontal_tile_24_29_to_tile_24_28_1),
		.out_wire_2_2(horizontal_tile_24_29_to_tile_24_28_2),
		.out_wire_2_3(horizontal_tile_24_29_to_tile_24_28_3),
		.in_wire_2_0(horizontal_tile_24_28_to_tile_24_29_0),
		.in_wire_2_1(horizontal_tile_24_28_to_tile_24_29_1),
		.in_wire_2_2(horizontal_tile_24_28_to_tile_24_29_2),
		.in_wire_2_3(horizontal_tile_24_28_to_tile_24_29_3),
		.out_wire_0_0(horizontal_tile_24_29_to_tile_24_30_0),
		.out_wire_0_1(horizontal_tile_24_29_to_tile_24_30_1),
		.out_wire_0_2(horizontal_tile_24_29_to_tile_24_30_2),
		.out_wire_0_3(horizontal_tile_24_29_to_tile_24_30_3),
		.in_wire_0_0(horizontal_tile_24_30_to_tile_24_29_0),
		.in_wire_0_1(horizontal_tile_24_30_to_tile_24_29_1),
		.in_wire_0_2(horizontal_tile_24_30_to_tile_24_29_2),
		.in_wire_0_3(horizontal_tile_24_30_to_tile_24_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(798)
	);

	pe_tile pe_tile_24_30(
		.out_wire_3_0(vertical_tile_24_30_to_tile_23_30_0),
		.out_wire_3_1(vertical_tile_24_30_to_tile_23_30_1),
		.out_wire_3_2(vertical_tile_24_30_to_tile_23_30_2),
		.out_wire_3_3(vertical_tile_24_30_to_tile_23_30_3),
		.in_wire_3_0(vertical_tile_23_30_to_tile_24_30_0),
		.in_wire_3_1(vertical_tile_23_30_to_tile_24_30_1),
		.in_wire_3_2(vertical_tile_23_30_to_tile_24_30_2),
		.in_wire_3_3(vertical_tile_23_30_to_tile_24_30_3),
		.out_wire_1_0(vertical_tile_24_30_to_tile_25_30_0),
		.out_wire_1_1(vertical_tile_24_30_to_tile_25_30_1),
		.out_wire_1_2(vertical_tile_24_30_to_tile_25_30_2),
		.out_wire_1_3(vertical_tile_24_30_to_tile_25_30_3),
		.in_wire_1_0(vertical_tile_25_30_to_tile_24_30_0),
		.in_wire_1_1(vertical_tile_25_30_to_tile_24_30_1),
		.in_wire_1_2(vertical_tile_25_30_to_tile_24_30_2),
		.in_wire_1_3(vertical_tile_25_30_to_tile_24_30_3),
		.out_wire_2_0(horizontal_tile_24_30_to_tile_24_29_0),
		.out_wire_2_1(horizontal_tile_24_30_to_tile_24_29_1),
		.out_wire_2_2(horizontal_tile_24_30_to_tile_24_29_2),
		.out_wire_2_3(horizontal_tile_24_30_to_tile_24_29_3),
		.in_wire_2_0(horizontal_tile_24_29_to_tile_24_30_0),
		.in_wire_2_1(horizontal_tile_24_29_to_tile_24_30_1),
		.in_wire_2_2(horizontal_tile_24_29_to_tile_24_30_2),
		.in_wire_2_3(horizontal_tile_24_29_to_tile_24_30_3),
		.out_wire_0_0(horizontal_tile_24_30_to_tile_24_31_0),
		.out_wire_0_1(horizontal_tile_24_30_to_tile_24_31_1),
		.out_wire_0_2(horizontal_tile_24_30_to_tile_24_31_2),
		.out_wire_0_3(horizontal_tile_24_30_to_tile_24_31_3),
		.in_wire_0_0(horizontal_tile_24_31_to_tile_24_30_0),
		.in_wire_0_1(horizontal_tile_24_31_to_tile_24_30_1),
		.in_wire_0_2(horizontal_tile_24_31_to_tile_24_30_2),
		.in_wire_0_3(horizontal_tile_24_31_to_tile_24_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(799)
	);

	pe_tile_right pe_tile_24_31(
		.out_wire_3_0(vertical_tile_24_31_to_tile_23_31_0),
		.out_wire_3_1(vertical_tile_24_31_to_tile_23_31_1),
		.out_wire_3_2(vertical_tile_24_31_to_tile_23_31_2),
		.out_wire_3_3(vertical_tile_24_31_to_tile_23_31_3),
		.in_wire_3_0(vertical_tile_23_31_to_tile_24_31_0),
		.in_wire_3_1(vertical_tile_23_31_to_tile_24_31_1),
		.in_wire_3_2(vertical_tile_23_31_to_tile_24_31_2),
		.in_wire_3_3(vertical_tile_23_31_to_tile_24_31_3),
		.out_wire_1_0(vertical_tile_24_31_to_tile_25_31_0),
		.out_wire_1_1(vertical_tile_24_31_to_tile_25_31_1),
		.out_wire_1_2(vertical_tile_24_31_to_tile_25_31_2),
		.out_wire_1_3(vertical_tile_24_31_to_tile_25_31_3),
		.in_wire_1_0(vertical_tile_25_31_to_tile_24_31_0),
		.in_wire_1_1(vertical_tile_25_31_to_tile_24_31_1),
		.in_wire_1_2(vertical_tile_25_31_to_tile_24_31_2),
		.in_wire_1_3(vertical_tile_25_31_to_tile_24_31_3),
		.out_wire_2_0(horizontal_tile_24_31_to_tile_24_30_0),
		.out_wire_2_1(horizontal_tile_24_31_to_tile_24_30_1),
		.out_wire_2_2(horizontal_tile_24_31_to_tile_24_30_2),
		.out_wire_2_3(horizontal_tile_24_31_to_tile_24_30_3),
		.in_wire_2_0(horizontal_tile_24_30_to_tile_24_31_0),
		.in_wire_2_1(horizontal_tile_24_30_to_tile_24_31_1),
		.in_wire_2_2(horizontal_tile_24_30_to_tile_24_31_2),
		.in_wire_2_3(horizontal_tile_24_30_to_tile_24_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(800)
	);

	pe_tile_left pe_tile_25_0(
		.out_wire_3_0(vertical_tile_25_0_to_tile_24_0_0),
		.out_wire_3_1(vertical_tile_25_0_to_tile_24_0_1),
		.out_wire_3_2(vertical_tile_25_0_to_tile_24_0_2),
		.out_wire_3_3(vertical_tile_25_0_to_tile_24_0_3),
		.in_wire_3_0(vertical_tile_24_0_to_tile_25_0_0),
		.in_wire_3_1(vertical_tile_24_0_to_tile_25_0_1),
		.in_wire_3_2(vertical_tile_24_0_to_tile_25_0_2),
		.in_wire_3_3(vertical_tile_24_0_to_tile_25_0_3),
		.out_wire_1_0(vertical_tile_25_0_to_tile_26_0_0),
		.out_wire_1_1(vertical_tile_25_0_to_tile_26_0_1),
		.out_wire_1_2(vertical_tile_25_0_to_tile_26_0_2),
		.out_wire_1_3(vertical_tile_25_0_to_tile_26_0_3),
		.in_wire_1_0(vertical_tile_26_0_to_tile_25_0_0),
		.in_wire_1_1(vertical_tile_26_0_to_tile_25_0_1),
		.in_wire_1_2(vertical_tile_26_0_to_tile_25_0_2),
		.in_wire_1_3(vertical_tile_26_0_to_tile_25_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_25_0_to_tile_25_1_0),
		.out_wire_0_1(horizontal_tile_25_0_to_tile_25_1_1),
		.out_wire_0_2(horizontal_tile_25_0_to_tile_25_1_2),
		.out_wire_0_3(horizontal_tile_25_0_to_tile_25_1_3),
		.in_wire_0_0(horizontal_tile_25_1_to_tile_25_0_0),
		.in_wire_0_1(horizontal_tile_25_1_to_tile_25_0_1),
		.in_wire_0_2(horizontal_tile_25_1_to_tile_25_0_2),
		.in_wire_0_3(horizontal_tile_25_1_to_tile_25_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(801)
	);

	pe_tile pe_tile_25_1(
		.out_wire_3_0(vertical_tile_25_1_to_tile_24_1_0),
		.out_wire_3_1(vertical_tile_25_1_to_tile_24_1_1),
		.out_wire_3_2(vertical_tile_25_1_to_tile_24_1_2),
		.out_wire_3_3(vertical_tile_25_1_to_tile_24_1_3),
		.in_wire_3_0(vertical_tile_24_1_to_tile_25_1_0),
		.in_wire_3_1(vertical_tile_24_1_to_tile_25_1_1),
		.in_wire_3_2(vertical_tile_24_1_to_tile_25_1_2),
		.in_wire_3_3(vertical_tile_24_1_to_tile_25_1_3),
		.out_wire_1_0(vertical_tile_25_1_to_tile_26_1_0),
		.out_wire_1_1(vertical_tile_25_1_to_tile_26_1_1),
		.out_wire_1_2(vertical_tile_25_1_to_tile_26_1_2),
		.out_wire_1_3(vertical_tile_25_1_to_tile_26_1_3),
		.in_wire_1_0(vertical_tile_26_1_to_tile_25_1_0),
		.in_wire_1_1(vertical_tile_26_1_to_tile_25_1_1),
		.in_wire_1_2(vertical_tile_26_1_to_tile_25_1_2),
		.in_wire_1_3(vertical_tile_26_1_to_tile_25_1_3),
		.out_wire_2_0(horizontal_tile_25_1_to_tile_25_0_0),
		.out_wire_2_1(horizontal_tile_25_1_to_tile_25_0_1),
		.out_wire_2_2(horizontal_tile_25_1_to_tile_25_0_2),
		.out_wire_2_3(horizontal_tile_25_1_to_tile_25_0_3),
		.in_wire_2_0(horizontal_tile_25_0_to_tile_25_1_0),
		.in_wire_2_1(horizontal_tile_25_0_to_tile_25_1_1),
		.in_wire_2_2(horizontal_tile_25_0_to_tile_25_1_2),
		.in_wire_2_3(horizontal_tile_25_0_to_tile_25_1_3),
		.out_wire_0_0(horizontal_tile_25_1_to_tile_25_2_0),
		.out_wire_0_1(horizontal_tile_25_1_to_tile_25_2_1),
		.out_wire_0_2(horizontal_tile_25_1_to_tile_25_2_2),
		.out_wire_0_3(horizontal_tile_25_1_to_tile_25_2_3),
		.in_wire_0_0(horizontal_tile_25_2_to_tile_25_1_0),
		.in_wire_0_1(horizontal_tile_25_2_to_tile_25_1_1),
		.in_wire_0_2(horizontal_tile_25_2_to_tile_25_1_2),
		.in_wire_0_3(horizontal_tile_25_2_to_tile_25_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(802)
	);

	pe_tile pe_tile_25_2(
		.out_wire_3_0(vertical_tile_25_2_to_tile_24_2_0),
		.out_wire_3_1(vertical_tile_25_2_to_tile_24_2_1),
		.out_wire_3_2(vertical_tile_25_2_to_tile_24_2_2),
		.out_wire_3_3(vertical_tile_25_2_to_tile_24_2_3),
		.in_wire_3_0(vertical_tile_24_2_to_tile_25_2_0),
		.in_wire_3_1(vertical_tile_24_2_to_tile_25_2_1),
		.in_wire_3_2(vertical_tile_24_2_to_tile_25_2_2),
		.in_wire_3_3(vertical_tile_24_2_to_tile_25_2_3),
		.out_wire_1_0(vertical_tile_25_2_to_tile_26_2_0),
		.out_wire_1_1(vertical_tile_25_2_to_tile_26_2_1),
		.out_wire_1_2(vertical_tile_25_2_to_tile_26_2_2),
		.out_wire_1_3(vertical_tile_25_2_to_tile_26_2_3),
		.in_wire_1_0(vertical_tile_26_2_to_tile_25_2_0),
		.in_wire_1_1(vertical_tile_26_2_to_tile_25_2_1),
		.in_wire_1_2(vertical_tile_26_2_to_tile_25_2_2),
		.in_wire_1_3(vertical_tile_26_2_to_tile_25_2_3),
		.out_wire_2_0(horizontal_tile_25_2_to_tile_25_1_0),
		.out_wire_2_1(horizontal_tile_25_2_to_tile_25_1_1),
		.out_wire_2_2(horizontal_tile_25_2_to_tile_25_1_2),
		.out_wire_2_3(horizontal_tile_25_2_to_tile_25_1_3),
		.in_wire_2_0(horizontal_tile_25_1_to_tile_25_2_0),
		.in_wire_2_1(horizontal_tile_25_1_to_tile_25_2_1),
		.in_wire_2_2(horizontal_tile_25_1_to_tile_25_2_2),
		.in_wire_2_3(horizontal_tile_25_1_to_tile_25_2_3),
		.out_wire_0_0(horizontal_tile_25_2_to_tile_25_3_0),
		.out_wire_0_1(horizontal_tile_25_2_to_tile_25_3_1),
		.out_wire_0_2(horizontal_tile_25_2_to_tile_25_3_2),
		.out_wire_0_3(horizontal_tile_25_2_to_tile_25_3_3),
		.in_wire_0_0(horizontal_tile_25_3_to_tile_25_2_0),
		.in_wire_0_1(horizontal_tile_25_3_to_tile_25_2_1),
		.in_wire_0_2(horizontal_tile_25_3_to_tile_25_2_2),
		.in_wire_0_3(horizontal_tile_25_3_to_tile_25_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(803)
	);

	pe_tile pe_tile_25_3(
		.out_wire_3_0(vertical_tile_25_3_to_tile_24_3_0),
		.out_wire_3_1(vertical_tile_25_3_to_tile_24_3_1),
		.out_wire_3_2(vertical_tile_25_3_to_tile_24_3_2),
		.out_wire_3_3(vertical_tile_25_3_to_tile_24_3_3),
		.in_wire_3_0(vertical_tile_24_3_to_tile_25_3_0),
		.in_wire_3_1(vertical_tile_24_3_to_tile_25_3_1),
		.in_wire_3_2(vertical_tile_24_3_to_tile_25_3_2),
		.in_wire_3_3(vertical_tile_24_3_to_tile_25_3_3),
		.out_wire_1_0(vertical_tile_25_3_to_tile_26_3_0),
		.out_wire_1_1(vertical_tile_25_3_to_tile_26_3_1),
		.out_wire_1_2(vertical_tile_25_3_to_tile_26_3_2),
		.out_wire_1_3(vertical_tile_25_3_to_tile_26_3_3),
		.in_wire_1_0(vertical_tile_26_3_to_tile_25_3_0),
		.in_wire_1_1(vertical_tile_26_3_to_tile_25_3_1),
		.in_wire_1_2(vertical_tile_26_3_to_tile_25_3_2),
		.in_wire_1_3(vertical_tile_26_3_to_tile_25_3_3),
		.out_wire_2_0(horizontal_tile_25_3_to_tile_25_2_0),
		.out_wire_2_1(horizontal_tile_25_3_to_tile_25_2_1),
		.out_wire_2_2(horizontal_tile_25_3_to_tile_25_2_2),
		.out_wire_2_3(horizontal_tile_25_3_to_tile_25_2_3),
		.in_wire_2_0(horizontal_tile_25_2_to_tile_25_3_0),
		.in_wire_2_1(horizontal_tile_25_2_to_tile_25_3_1),
		.in_wire_2_2(horizontal_tile_25_2_to_tile_25_3_2),
		.in_wire_2_3(horizontal_tile_25_2_to_tile_25_3_3),
		.out_wire_0_0(horizontal_tile_25_3_to_tile_25_4_0),
		.out_wire_0_1(horizontal_tile_25_3_to_tile_25_4_1),
		.out_wire_0_2(horizontal_tile_25_3_to_tile_25_4_2),
		.out_wire_0_3(horizontal_tile_25_3_to_tile_25_4_3),
		.in_wire_0_0(horizontal_tile_25_4_to_tile_25_3_0),
		.in_wire_0_1(horizontal_tile_25_4_to_tile_25_3_1),
		.in_wire_0_2(horizontal_tile_25_4_to_tile_25_3_2),
		.in_wire_0_3(horizontal_tile_25_4_to_tile_25_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(804)
	);

	pe_tile pe_tile_25_4(
		.out_wire_3_0(vertical_tile_25_4_to_tile_24_4_0),
		.out_wire_3_1(vertical_tile_25_4_to_tile_24_4_1),
		.out_wire_3_2(vertical_tile_25_4_to_tile_24_4_2),
		.out_wire_3_3(vertical_tile_25_4_to_tile_24_4_3),
		.in_wire_3_0(vertical_tile_24_4_to_tile_25_4_0),
		.in_wire_3_1(vertical_tile_24_4_to_tile_25_4_1),
		.in_wire_3_2(vertical_tile_24_4_to_tile_25_4_2),
		.in_wire_3_3(vertical_tile_24_4_to_tile_25_4_3),
		.out_wire_1_0(vertical_tile_25_4_to_tile_26_4_0),
		.out_wire_1_1(vertical_tile_25_4_to_tile_26_4_1),
		.out_wire_1_2(vertical_tile_25_4_to_tile_26_4_2),
		.out_wire_1_3(vertical_tile_25_4_to_tile_26_4_3),
		.in_wire_1_0(vertical_tile_26_4_to_tile_25_4_0),
		.in_wire_1_1(vertical_tile_26_4_to_tile_25_4_1),
		.in_wire_1_2(vertical_tile_26_4_to_tile_25_4_2),
		.in_wire_1_3(vertical_tile_26_4_to_tile_25_4_3),
		.out_wire_2_0(horizontal_tile_25_4_to_tile_25_3_0),
		.out_wire_2_1(horizontal_tile_25_4_to_tile_25_3_1),
		.out_wire_2_2(horizontal_tile_25_4_to_tile_25_3_2),
		.out_wire_2_3(horizontal_tile_25_4_to_tile_25_3_3),
		.in_wire_2_0(horizontal_tile_25_3_to_tile_25_4_0),
		.in_wire_2_1(horizontal_tile_25_3_to_tile_25_4_1),
		.in_wire_2_2(horizontal_tile_25_3_to_tile_25_4_2),
		.in_wire_2_3(horizontal_tile_25_3_to_tile_25_4_3),
		.out_wire_0_0(horizontal_tile_25_4_to_tile_25_5_0),
		.out_wire_0_1(horizontal_tile_25_4_to_tile_25_5_1),
		.out_wire_0_2(horizontal_tile_25_4_to_tile_25_5_2),
		.out_wire_0_3(horizontal_tile_25_4_to_tile_25_5_3),
		.in_wire_0_0(horizontal_tile_25_5_to_tile_25_4_0),
		.in_wire_0_1(horizontal_tile_25_5_to_tile_25_4_1),
		.in_wire_0_2(horizontal_tile_25_5_to_tile_25_4_2),
		.in_wire_0_3(horizontal_tile_25_5_to_tile_25_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(805)
	);

	pe_tile pe_tile_25_5(
		.out_wire_3_0(vertical_tile_25_5_to_tile_24_5_0),
		.out_wire_3_1(vertical_tile_25_5_to_tile_24_5_1),
		.out_wire_3_2(vertical_tile_25_5_to_tile_24_5_2),
		.out_wire_3_3(vertical_tile_25_5_to_tile_24_5_3),
		.in_wire_3_0(vertical_tile_24_5_to_tile_25_5_0),
		.in_wire_3_1(vertical_tile_24_5_to_tile_25_5_1),
		.in_wire_3_2(vertical_tile_24_5_to_tile_25_5_2),
		.in_wire_3_3(vertical_tile_24_5_to_tile_25_5_3),
		.out_wire_1_0(vertical_tile_25_5_to_tile_26_5_0),
		.out_wire_1_1(vertical_tile_25_5_to_tile_26_5_1),
		.out_wire_1_2(vertical_tile_25_5_to_tile_26_5_2),
		.out_wire_1_3(vertical_tile_25_5_to_tile_26_5_3),
		.in_wire_1_0(vertical_tile_26_5_to_tile_25_5_0),
		.in_wire_1_1(vertical_tile_26_5_to_tile_25_5_1),
		.in_wire_1_2(vertical_tile_26_5_to_tile_25_5_2),
		.in_wire_1_3(vertical_tile_26_5_to_tile_25_5_3),
		.out_wire_2_0(horizontal_tile_25_5_to_tile_25_4_0),
		.out_wire_2_1(horizontal_tile_25_5_to_tile_25_4_1),
		.out_wire_2_2(horizontal_tile_25_5_to_tile_25_4_2),
		.out_wire_2_3(horizontal_tile_25_5_to_tile_25_4_3),
		.in_wire_2_0(horizontal_tile_25_4_to_tile_25_5_0),
		.in_wire_2_1(horizontal_tile_25_4_to_tile_25_5_1),
		.in_wire_2_2(horizontal_tile_25_4_to_tile_25_5_2),
		.in_wire_2_3(horizontal_tile_25_4_to_tile_25_5_3),
		.out_wire_0_0(horizontal_tile_25_5_to_tile_25_6_0),
		.out_wire_0_1(horizontal_tile_25_5_to_tile_25_6_1),
		.out_wire_0_2(horizontal_tile_25_5_to_tile_25_6_2),
		.out_wire_0_3(horizontal_tile_25_5_to_tile_25_6_3),
		.in_wire_0_0(horizontal_tile_25_6_to_tile_25_5_0),
		.in_wire_0_1(horizontal_tile_25_6_to_tile_25_5_1),
		.in_wire_0_2(horizontal_tile_25_6_to_tile_25_5_2),
		.in_wire_0_3(horizontal_tile_25_6_to_tile_25_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(806)
	);

	pe_tile pe_tile_25_6(
		.out_wire_3_0(vertical_tile_25_6_to_tile_24_6_0),
		.out_wire_3_1(vertical_tile_25_6_to_tile_24_6_1),
		.out_wire_3_2(vertical_tile_25_6_to_tile_24_6_2),
		.out_wire_3_3(vertical_tile_25_6_to_tile_24_6_3),
		.in_wire_3_0(vertical_tile_24_6_to_tile_25_6_0),
		.in_wire_3_1(vertical_tile_24_6_to_tile_25_6_1),
		.in_wire_3_2(vertical_tile_24_6_to_tile_25_6_2),
		.in_wire_3_3(vertical_tile_24_6_to_tile_25_6_3),
		.out_wire_1_0(vertical_tile_25_6_to_tile_26_6_0),
		.out_wire_1_1(vertical_tile_25_6_to_tile_26_6_1),
		.out_wire_1_2(vertical_tile_25_6_to_tile_26_6_2),
		.out_wire_1_3(vertical_tile_25_6_to_tile_26_6_3),
		.in_wire_1_0(vertical_tile_26_6_to_tile_25_6_0),
		.in_wire_1_1(vertical_tile_26_6_to_tile_25_6_1),
		.in_wire_1_2(vertical_tile_26_6_to_tile_25_6_2),
		.in_wire_1_3(vertical_tile_26_6_to_tile_25_6_3),
		.out_wire_2_0(horizontal_tile_25_6_to_tile_25_5_0),
		.out_wire_2_1(horizontal_tile_25_6_to_tile_25_5_1),
		.out_wire_2_2(horizontal_tile_25_6_to_tile_25_5_2),
		.out_wire_2_3(horizontal_tile_25_6_to_tile_25_5_3),
		.in_wire_2_0(horizontal_tile_25_5_to_tile_25_6_0),
		.in_wire_2_1(horizontal_tile_25_5_to_tile_25_6_1),
		.in_wire_2_2(horizontal_tile_25_5_to_tile_25_6_2),
		.in_wire_2_3(horizontal_tile_25_5_to_tile_25_6_3),
		.out_wire_0_0(horizontal_tile_25_6_to_tile_25_7_0),
		.out_wire_0_1(horizontal_tile_25_6_to_tile_25_7_1),
		.out_wire_0_2(horizontal_tile_25_6_to_tile_25_7_2),
		.out_wire_0_3(horizontal_tile_25_6_to_tile_25_7_3),
		.in_wire_0_0(horizontal_tile_25_7_to_tile_25_6_0),
		.in_wire_0_1(horizontal_tile_25_7_to_tile_25_6_1),
		.in_wire_0_2(horizontal_tile_25_7_to_tile_25_6_2),
		.in_wire_0_3(horizontal_tile_25_7_to_tile_25_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(807)
	);

	pe_tile pe_tile_25_7(
		.out_wire_3_0(vertical_tile_25_7_to_tile_24_7_0),
		.out_wire_3_1(vertical_tile_25_7_to_tile_24_7_1),
		.out_wire_3_2(vertical_tile_25_7_to_tile_24_7_2),
		.out_wire_3_3(vertical_tile_25_7_to_tile_24_7_3),
		.in_wire_3_0(vertical_tile_24_7_to_tile_25_7_0),
		.in_wire_3_1(vertical_tile_24_7_to_tile_25_7_1),
		.in_wire_3_2(vertical_tile_24_7_to_tile_25_7_2),
		.in_wire_3_3(vertical_tile_24_7_to_tile_25_7_3),
		.out_wire_1_0(vertical_tile_25_7_to_tile_26_7_0),
		.out_wire_1_1(vertical_tile_25_7_to_tile_26_7_1),
		.out_wire_1_2(vertical_tile_25_7_to_tile_26_7_2),
		.out_wire_1_3(vertical_tile_25_7_to_tile_26_7_3),
		.in_wire_1_0(vertical_tile_26_7_to_tile_25_7_0),
		.in_wire_1_1(vertical_tile_26_7_to_tile_25_7_1),
		.in_wire_1_2(vertical_tile_26_7_to_tile_25_7_2),
		.in_wire_1_3(vertical_tile_26_7_to_tile_25_7_3),
		.out_wire_2_0(horizontal_tile_25_7_to_tile_25_6_0),
		.out_wire_2_1(horizontal_tile_25_7_to_tile_25_6_1),
		.out_wire_2_2(horizontal_tile_25_7_to_tile_25_6_2),
		.out_wire_2_3(horizontal_tile_25_7_to_tile_25_6_3),
		.in_wire_2_0(horizontal_tile_25_6_to_tile_25_7_0),
		.in_wire_2_1(horizontal_tile_25_6_to_tile_25_7_1),
		.in_wire_2_2(horizontal_tile_25_6_to_tile_25_7_2),
		.in_wire_2_3(horizontal_tile_25_6_to_tile_25_7_3),
		.out_wire_0_0(horizontal_tile_25_7_to_tile_25_8_0),
		.out_wire_0_1(horizontal_tile_25_7_to_tile_25_8_1),
		.out_wire_0_2(horizontal_tile_25_7_to_tile_25_8_2),
		.out_wire_0_3(horizontal_tile_25_7_to_tile_25_8_3),
		.in_wire_0_0(horizontal_tile_25_8_to_tile_25_7_0),
		.in_wire_0_1(horizontal_tile_25_8_to_tile_25_7_1),
		.in_wire_0_2(horizontal_tile_25_8_to_tile_25_7_2),
		.in_wire_0_3(horizontal_tile_25_8_to_tile_25_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(808)
	);

	pe_tile pe_tile_25_8(
		.out_wire_3_0(vertical_tile_25_8_to_tile_24_8_0),
		.out_wire_3_1(vertical_tile_25_8_to_tile_24_8_1),
		.out_wire_3_2(vertical_tile_25_8_to_tile_24_8_2),
		.out_wire_3_3(vertical_tile_25_8_to_tile_24_8_3),
		.in_wire_3_0(vertical_tile_24_8_to_tile_25_8_0),
		.in_wire_3_1(vertical_tile_24_8_to_tile_25_8_1),
		.in_wire_3_2(vertical_tile_24_8_to_tile_25_8_2),
		.in_wire_3_3(vertical_tile_24_8_to_tile_25_8_3),
		.out_wire_1_0(vertical_tile_25_8_to_tile_26_8_0),
		.out_wire_1_1(vertical_tile_25_8_to_tile_26_8_1),
		.out_wire_1_2(vertical_tile_25_8_to_tile_26_8_2),
		.out_wire_1_3(vertical_tile_25_8_to_tile_26_8_3),
		.in_wire_1_0(vertical_tile_26_8_to_tile_25_8_0),
		.in_wire_1_1(vertical_tile_26_8_to_tile_25_8_1),
		.in_wire_1_2(vertical_tile_26_8_to_tile_25_8_2),
		.in_wire_1_3(vertical_tile_26_8_to_tile_25_8_3),
		.out_wire_2_0(horizontal_tile_25_8_to_tile_25_7_0),
		.out_wire_2_1(horizontal_tile_25_8_to_tile_25_7_1),
		.out_wire_2_2(horizontal_tile_25_8_to_tile_25_7_2),
		.out_wire_2_3(horizontal_tile_25_8_to_tile_25_7_3),
		.in_wire_2_0(horizontal_tile_25_7_to_tile_25_8_0),
		.in_wire_2_1(horizontal_tile_25_7_to_tile_25_8_1),
		.in_wire_2_2(horizontal_tile_25_7_to_tile_25_8_2),
		.in_wire_2_3(horizontal_tile_25_7_to_tile_25_8_3),
		.out_wire_0_0(horizontal_tile_25_8_to_tile_25_9_0),
		.out_wire_0_1(horizontal_tile_25_8_to_tile_25_9_1),
		.out_wire_0_2(horizontal_tile_25_8_to_tile_25_9_2),
		.out_wire_0_3(horizontal_tile_25_8_to_tile_25_9_3),
		.in_wire_0_0(horizontal_tile_25_9_to_tile_25_8_0),
		.in_wire_0_1(horizontal_tile_25_9_to_tile_25_8_1),
		.in_wire_0_2(horizontal_tile_25_9_to_tile_25_8_2),
		.in_wire_0_3(horizontal_tile_25_9_to_tile_25_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(809)
	);

	pe_tile pe_tile_25_9(
		.out_wire_3_0(vertical_tile_25_9_to_tile_24_9_0),
		.out_wire_3_1(vertical_tile_25_9_to_tile_24_9_1),
		.out_wire_3_2(vertical_tile_25_9_to_tile_24_9_2),
		.out_wire_3_3(vertical_tile_25_9_to_tile_24_9_3),
		.in_wire_3_0(vertical_tile_24_9_to_tile_25_9_0),
		.in_wire_3_1(vertical_tile_24_9_to_tile_25_9_1),
		.in_wire_3_2(vertical_tile_24_9_to_tile_25_9_2),
		.in_wire_3_3(vertical_tile_24_9_to_tile_25_9_3),
		.out_wire_1_0(vertical_tile_25_9_to_tile_26_9_0),
		.out_wire_1_1(vertical_tile_25_9_to_tile_26_9_1),
		.out_wire_1_2(vertical_tile_25_9_to_tile_26_9_2),
		.out_wire_1_3(vertical_tile_25_9_to_tile_26_9_3),
		.in_wire_1_0(vertical_tile_26_9_to_tile_25_9_0),
		.in_wire_1_1(vertical_tile_26_9_to_tile_25_9_1),
		.in_wire_1_2(vertical_tile_26_9_to_tile_25_9_2),
		.in_wire_1_3(vertical_tile_26_9_to_tile_25_9_3),
		.out_wire_2_0(horizontal_tile_25_9_to_tile_25_8_0),
		.out_wire_2_1(horizontal_tile_25_9_to_tile_25_8_1),
		.out_wire_2_2(horizontal_tile_25_9_to_tile_25_8_2),
		.out_wire_2_3(horizontal_tile_25_9_to_tile_25_8_3),
		.in_wire_2_0(horizontal_tile_25_8_to_tile_25_9_0),
		.in_wire_2_1(horizontal_tile_25_8_to_tile_25_9_1),
		.in_wire_2_2(horizontal_tile_25_8_to_tile_25_9_2),
		.in_wire_2_3(horizontal_tile_25_8_to_tile_25_9_3),
		.out_wire_0_0(horizontal_tile_25_9_to_tile_25_10_0),
		.out_wire_0_1(horizontal_tile_25_9_to_tile_25_10_1),
		.out_wire_0_2(horizontal_tile_25_9_to_tile_25_10_2),
		.out_wire_0_3(horizontal_tile_25_9_to_tile_25_10_3),
		.in_wire_0_0(horizontal_tile_25_10_to_tile_25_9_0),
		.in_wire_0_1(horizontal_tile_25_10_to_tile_25_9_1),
		.in_wire_0_2(horizontal_tile_25_10_to_tile_25_9_2),
		.in_wire_0_3(horizontal_tile_25_10_to_tile_25_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(810)
	);

	pe_tile pe_tile_25_10(
		.out_wire_3_0(vertical_tile_25_10_to_tile_24_10_0),
		.out_wire_3_1(vertical_tile_25_10_to_tile_24_10_1),
		.out_wire_3_2(vertical_tile_25_10_to_tile_24_10_2),
		.out_wire_3_3(vertical_tile_25_10_to_tile_24_10_3),
		.in_wire_3_0(vertical_tile_24_10_to_tile_25_10_0),
		.in_wire_3_1(vertical_tile_24_10_to_tile_25_10_1),
		.in_wire_3_2(vertical_tile_24_10_to_tile_25_10_2),
		.in_wire_3_3(vertical_tile_24_10_to_tile_25_10_3),
		.out_wire_1_0(vertical_tile_25_10_to_tile_26_10_0),
		.out_wire_1_1(vertical_tile_25_10_to_tile_26_10_1),
		.out_wire_1_2(vertical_tile_25_10_to_tile_26_10_2),
		.out_wire_1_3(vertical_tile_25_10_to_tile_26_10_3),
		.in_wire_1_0(vertical_tile_26_10_to_tile_25_10_0),
		.in_wire_1_1(vertical_tile_26_10_to_tile_25_10_1),
		.in_wire_1_2(vertical_tile_26_10_to_tile_25_10_2),
		.in_wire_1_3(vertical_tile_26_10_to_tile_25_10_3),
		.out_wire_2_0(horizontal_tile_25_10_to_tile_25_9_0),
		.out_wire_2_1(horizontal_tile_25_10_to_tile_25_9_1),
		.out_wire_2_2(horizontal_tile_25_10_to_tile_25_9_2),
		.out_wire_2_3(horizontal_tile_25_10_to_tile_25_9_3),
		.in_wire_2_0(horizontal_tile_25_9_to_tile_25_10_0),
		.in_wire_2_1(horizontal_tile_25_9_to_tile_25_10_1),
		.in_wire_2_2(horizontal_tile_25_9_to_tile_25_10_2),
		.in_wire_2_3(horizontal_tile_25_9_to_tile_25_10_3),
		.out_wire_0_0(horizontal_tile_25_10_to_tile_25_11_0),
		.out_wire_0_1(horizontal_tile_25_10_to_tile_25_11_1),
		.out_wire_0_2(horizontal_tile_25_10_to_tile_25_11_2),
		.out_wire_0_3(horizontal_tile_25_10_to_tile_25_11_3),
		.in_wire_0_0(horizontal_tile_25_11_to_tile_25_10_0),
		.in_wire_0_1(horizontal_tile_25_11_to_tile_25_10_1),
		.in_wire_0_2(horizontal_tile_25_11_to_tile_25_10_2),
		.in_wire_0_3(horizontal_tile_25_11_to_tile_25_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(811)
	);

	pe_tile pe_tile_25_11(
		.out_wire_3_0(vertical_tile_25_11_to_tile_24_11_0),
		.out_wire_3_1(vertical_tile_25_11_to_tile_24_11_1),
		.out_wire_3_2(vertical_tile_25_11_to_tile_24_11_2),
		.out_wire_3_3(vertical_tile_25_11_to_tile_24_11_3),
		.in_wire_3_0(vertical_tile_24_11_to_tile_25_11_0),
		.in_wire_3_1(vertical_tile_24_11_to_tile_25_11_1),
		.in_wire_3_2(vertical_tile_24_11_to_tile_25_11_2),
		.in_wire_3_3(vertical_tile_24_11_to_tile_25_11_3),
		.out_wire_1_0(vertical_tile_25_11_to_tile_26_11_0),
		.out_wire_1_1(vertical_tile_25_11_to_tile_26_11_1),
		.out_wire_1_2(vertical_tile_25_11_to_tile_26_11_2),
		.out_wire_1_3(vertical_tile_25_11_to_tile_26_11_3),
		.in_wire_1_0(vertical_tile_26_11_to_tile_25_11_0),
		.in_wire_1_1(vertical_tile_26_11_to_tile_25_11_1),
		.in_wire_1_2(vertical_tile_26_11_to_tile_25_11_2),
		.in_wire_1_3(vertical_tile_26_11_to_tile_25_11_3),
		.out_wire_2_0(horizontal_tile_25_11_to_tile_25_10_0),
		.out_wire_2_1(horizontal_tile_25_11_to_tile_25_10_1),
		.out_wire_2_2(horizontal_tile_25_11_to_tile_25_10_2),
		.out_wire_2_3(horizontal_tile_25_11_to_tile_25_10_3),
		.in_wire_2_0(horizontal_tile_25_10_to_tile_25_11_0),
		.in_wire_2_1(horizontal_tile_25_10_to_tile_25_11_1),
		.in_wire_2_2(horizontal_tile_25_10_to_tile_25_11_2),
		.in_wire_2_3(horizontal_tile_25_10_to_tile_25_11_3),
		.out_wire_0_0(horizontal_tile_25_11_to_tile_25_12_0),
		.out_wire_0_1(horizontal_tile_25_11_to_tile_25_12_1),
		.out_wire_0_2(horizontal_tile_25_11_to_tile_25_12_2),
		.out_wire_0_3(horizontal_tile_25_11_to_tile_25_12_3),
		.in_wire_0_0(horizontal_tile_25_12_to_tile_25_11_0),
		.in_wire_0_1(horizontal_tile_25_12_to_tile_25_11_1),
		.in_wire_0_2(horizontal_tile_25_12_to_tile_25_11_2),
		.in_wire_0_3(horizontal_tile_25_12_to_tile_25_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(812)
	);

	pe_tile pe_tile_25_12(
		.out_wire_3_0(vertical_tile_25_12_to_tile_24_12_0),
		.out_wire_3_1(vertical_tile_25_12_to_tile_24_12_1),
		.out_wire_3_2(vertical_tile_25_12_to_tile_24_12_2),
		.out_wire_3_3(vertical_tile_25_12_to_tile_24_12_3),
		.in_wire_3_0(vertical_tile_24_12_to_tile_25_12_0),
		.in_wire_3_1(vertical_tile_24_12_to_tile_25_12_1),
		.in_wire_3_2(vertical_tile_24_12_to_tile_25_12_2),
		.in_wire_3_3(vertical_tile_24_12_to_tile_25_12_3),
		.out_wire_1_0(vertical_tile_25_12_to_tile_26_12_0),
		.out_wire_1_1(vertical_tile_25_12_to_tile_26_12_1),
		.out_wire_1_2(vertical_tile_25_12_to_tile_26_12_2),
		.out_wire_1_3(vertical_tile_25_12_to_tile_26_12_3),
		.in_wire_1_0(vertical_tile_26_12_to_tile_25_12_0),
		.in_wire_1_1(vertical_tile_26_12_to_tile_25_12_1),
		.in_wire_1_2(vertical_tile_26_12_to_tile_25_12_2),
		.in_wire_1_3(vertical_tile_26_12_to_tile_25_12_3),
		.out_wire_2_0(horizontal_tile_25_12_to_tile_25_11_0),
		.out_wire_2_1(horizontal_tile_25_12_to_tile_25_11_1),
		.out_wire_2_2(horizontal_tile_25_12_to_tile_25_11_2),
		.out_wire_2_3(horizontal_tile_25_12_to_tile_25_11_3),
		.in_wire_2_0(horizontal_tile_25_11_to_tile_25_12_0),
		.in_wire_2_1(horizontal_tile_25_11_to_tile_25_12_1),
		.in_wire_2_2(horizontal_tile_25_11_to_tile_25_12_2),
		.in_wire_2_3(horizontal_tile_25_11_to_tile_25_12_3),
		.out_wire_0_0(horizontal_tile_25_12_to_tile_25_13_0),
		.out_wire_0_1(horizontal_tile_25_12_to_tile_25_13_1),
		.out_wire_0_2(horizontal_tile_25_12_to_tile_25_13_2),
		.out_wire_0_3(horizontal_tile_25_12_to_tile_25_13_3),
		.in_wire_0_0(horizontal_tile_25_13_to_tile_25_12_0),
		.in_wire_0_1(horizontal_tile_25_13_to_tile_25_12_1),
		.in_wire_0_2(horizontal_tile_25_13_to_tile_25_12_2),
		.in_wire_0_3(horizontal_tile_25_13_to_tile_25_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(813)
	);

	pe_tile pe_tile_25_13(
		.out_wire_3_0(vertical_tile_25_13_to_tile_24_13_0),
		.out_wire_3_1(vertical_tile_25_13_to_tile_24_13_1),
		.out_wire_3_2(vertical_tile_25_13_to_tile_24_13_2),
		.out_wire_3_3(vertical_tile_25_13_to_tile_24_13_3),
		.in_wire_3_0(vertical_tile_24_13_to_tile_25_13_0),
		.in_wire_3_1(vertical_tile_24_13_to_tile_25_13_1),
		.in_wire_3_2(vertical_tile_24_13_to_tile_25_13_2),
		.in_wire_3_3(vertical_tile_24_13_to_tile_25_13_3),
		.out_wire_1_0(vertical_tile_25_13_to_tile_26_13_0),
		.out_wire_1_1(vertical_tile_25_13_to_tile_26_13_1),
		.out_wire_1_2(vertical_tile_25_13_to_tile_26_13_2),
		.out_wire_1_3(vertical_tile_25_13_to_tile_26_13_3),
		.in_wire_1_0(vertical_tile_26_13_to_tile_25_13_0),
		.in_wire_1_1(vertical_tile_26_13_to_tile_25_13_1),
		.in_wire_1_2(vertical_tile_26_13_to_tile_25_13_2),
		.in_wire_1_3(vertical_tile_26_13_to_tile_25_13_3),
		.out_wire_2_0(horizontal_tile_25_13_to_tile_25_12_0),
		.out_wire_2_1(horizontal_tile_25_13_to_tile_25_12_1),
		.out_wire_2_2(horizontal_tile_25_13_to_tile_25_12_2),
		.out_wire_2_3(horizontal_tile_25_13_to_tile_25_12_3),
		.in_wire_2_0(horizontal_tile_25_12_to_tile_25_13_0),
		.in_wire_2_1(horizontal_tile_25_12_to_tile_25_13_1),
		.in_wire_2_2(horizontal_tile_25_12_to_tile_25_13_2),
		.in_wire_2_3(horizontal_tile_25_12_to_tile_25_13_3),
		.out_wire_0_0(horizontal_tile_25_13_to_tile_25_14_0),
		.out_wire_0_1(horizontal_tile_25_13_to_tile_25_14_1),
		.out_wire_0_2(horizontal_tile_25_13_to_tile_25_14_2),
		.out_wire_0_3(horizontal_tile_25_13_to_tile_25_14_3),
		.in_wire_0_0(horizontal_tile_25_14_to_tile_25_13_0),
		.in_wire_0_1(horizontal_tile_25_14_to_tile_25_13_1),
		.in_wire_0_2(horizontal_tile_25_14_to_tile_25_13_2),
		.in_wire_0_3(horizontal_tile_25_14_to_tile_25_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(814)
	);

	pe_tile pe_tile_25_14(
		.out_wire_3_0(vertical_tile_25_14_to_tile_24_14_0),
		.out_wire_3_1(vertical_tile_25_14_to_tile_24_14_1),
		.out_wire_3_2(vertical_tile_25_14_to_tile_24_14_2),
		.out_wire_3_3(vertical_tile_25_14_to_tile_24_14_3),
		.in_wire_3_0(vertical_tile_24_14_to_tile_25_14_0),
		.in_wire_3_1(vertical_tile_24_14_to_tile_25_14_1),
		.in_wire_3_2(vertical_tile_24_14_to_tile_25_14_2),
		.in_wire_3_3(vertical_tile_24_14_to_tile_25_14_3),
		.out_wire_1_0(vertical_tile_25_14_to_tile_26_14_0),
		.out_wire_1_1(vertical_tile_25_14_to_tile_26_14_1),
		.out_wire_1_2(vertical_tile_25_14_to_tile_26_14_2),
		.out_wire_1_3(vertical_tile_25_14_to_tile_26_14_3),
		.in_wire_1_0(vertical_tile_26_14_to_tile_25_14_0),
		.in_wire_1_1(vertical_tile_26_14_to_tile_25_14_1),
		.in_wire_1_2(vertical_tile_26_14_to_tile_25_14_2),
		.in_wire_1_3(vertical_tile_26_14_to_tile_25_14_3),
		.out_wire_2_0(horizontal_tile_25_14_to_tile_25_13_0),
		.out_wire_2_1(horizontal_tile_25_14_to_tile_25_13_1),
		.out_wire_2_2(horizontal_tile_25_14_to_tile_25_13_2),
		.out_wire_2_3(horizontal_tile_25_14_to_tile_25_13_3),
		.in_wire_2_0(horizontal_tile_25_13_to_tile_25_14_0),
		.in_wire_2_1(horizontal_tile_25_13_to_tile_25_14_1),
		.in_wire_2_2(horizontal_tile_25_13_to_tile_25_14_2),
		.in_wire_2_3(horizontal_tile_25_13_to_tile_25_14_3),
		.out_wire_0_0(horizontal_tile_25_14_to_tile_25_15_0),
		.out_wire_0_1(horizontal_tile_25_14_to_tile_25_15_1),
		.out_wire_0_2(horizontal_tile_25_14_to_tile_25_15_2),
		.out_wire_0_3(horizontal_tile_25_14_to_tile_25_15_3),
		.in_wire_0_0(horizontal_tile_25_15_to_tile_25_14_0),
		.in_wire_0_1(horizontal_tile_25_15_to_tile_25_14_1),
		.in_wire_0_2(horizontal_tile_25_15_to_tile_25_14_2),
		.in_wire_0_3(horizontal_tile_25_15_to_tile_25_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(815)
	);

	pe_tile pe_tile_25_15(
		.out_wire_3_0(vertical_tile_25_15_to_tile_24_15_0),
		.out_wire_3_1(vertical_tile_25_15_to_tile_24_15_1),
		.out_wire_3_2(vertical_tile_25_15_to_tile_24_15_2),
		.out_wire_3_3(vertical_tile_25_15_to_tile_24_15_3),
		.in_wire_3_0(vertical_tile_24_15_to_tile_25_15_0),
		.in_wire_3_1(vertical_tile_24_15_to_tile_25_15_1),
		.in_wire_3_2(vertical_tile_24_15_to_tile_25_15_2),
		.in_wire_3_3(vertical_tile_24_15_to_tile_25_15_3),
		.out_wire_1_0(vertical_tile_25_15_to_tile_26_15_0),
		.out_wire_1_1(vertical_tile_25_15_to_tile_26_15_1),
		.out_wire_1_2(vertical_tile_25_15_to_tile_26_15_2),
		.out_wire_1_3(vertical_tile_25_15_to_tile_26_15_3),
		.in_wire_1_0(vertical_tile_26_15_to_tile_25_15_0),
		.in_wire_1_1(vertical_tile_26_15_to_tile_25_15_1),
		.in_wire_1_2(vertical_tile_26_15_to_tile_25_15_2),
		.in_wire_1_3(vertical_tile_26_15_to_tile_25_15_3),
		.out_wire_2_0(horizontal_tile_25_15_to_tile_25_14_0),
		.out_wire_2_1(horizontal_tile_25_15_to_tile_25_14_1),
		.out_wire_2_2(horizontal_tile_25_15_to_tile_25_14_2),
		.out_wire_2_3(horizontal_tile_25_15_to_tile_25_14_3),
		.in_wire_2_0(horizontal_tile_25_14_to_tile_25_15_0),
		.in_wire_2_1(horizontal_tile_25_14_to_tile_25_15_1),
		.in_wire_2_2(horizontal_tile_25_14_to_tile_25_15_2),
		.in_wire_2_3(horizontal_tile_25_14_to_tile_25_15_3),
		.out_wire_0_0(horizontal_tile_25_15_to_tile_25_16_0),
		.out_wire_0_1(horizontal_tile_25_15_to_tile_25_16_1),
		.out_wire_0_2(horizontal_tile_25_15_to_tile_25_16_2),
		.out_wire_0_3(horizontal_tile_25_15_to_tile_25_16_3),
		.in_wire_0_0(horizontal_tile_25_16_to_tile_25_15_0),
		.in_wire_0_1(horizontal_tile_25_16_to_tile_25_15_1),
		.in_wire_0_2(horizontal_tile_25_16_to_tile_25_15_2),
		.in_wire_0_3(horizontal_tile_25_16_to_tile_25_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(816)
	);

	pe_tile pe_tile_25_16(
		.out_wire_3_0(vertical_tile_25_16_to_tile_24_16_0),
		.out_wire_3_1(vertical_tile_25_16_to_tile_24_16_1),
		.out_wire_3_2(vertical_tile_25_16_to_tile_24_16_2),
		.out_wire_3_3(vertical_tile_25_16_to_tile_24_16_3),
		.in_wire_3_0(vertical_tile_24_16_to_tile_25_16_0),
		.in_wire_3_1(vertical_tile_24_16_to_tile_25_16_1),
		.in_wire_3_2(vertical_tile_24_16_to_tile_25_16_2),
		.in_wire_3_3(vertical_tile_24_16_to_tile_25_16_3),
		.out_wire_1_0(vertical_tile_25_16_to_tile_26_16_0),
		.out_wire_1_1(vertical_tile_25_16_to_tile_26_16_1),
		.out_wire_1_2(vertical_tile_25_16_to_tile_26_16_2),
		.out_wire_1_3(vertical_tile_25_16_to_tile_26_16_3),
		.in_wire_1_0(vertical_tile_26_16_to_tile_25_16_0),
		.in_wire_1_1(vertical_tile_26_16_to_tile_25_16_1),
		.in_wire_1_2(vertical_tile_26_16_to_tile_25_16_2),
		.in_wire_1_3(vertical_tile_26_16_to_tile_25_16_3),
		.out_wire_2_0(horizontal_tile_25_16_to_tile_25_15_0),
		.out_wire_2_1(horizontal_tile_25_16_to_tile_25_15_1),
		.out_wire_2_2(horizontal_tile_25_16_to_tile_25_15_2),
		.out_wire_2_3(horizontal_tile_25_16_to_tile_25_15_3),
		.in_wire_2_0(horizontal_tile_25_15_to_tile_25_16_0),
		.in_wire_2_1(horizontal_tile_25_15_to_tile_25_16_1),
		.in_wire_2_2(horizontal_tile_25_15_to_tile_25_16_2),
		.in_wire_2_3(horizontal_tile_25_15_to_tile_25_16_3),
		.out_wire_0_0(horizontal_tile_25_16_to_tile_25_17_0),
		.out_wire_0_1(horizontal_tile_25_16_to_tile_25_17_1),
		.out_wire_0_2(horizontal_tile_25_16_to_tile_25_17_2),
		.out_wire_0_3(horizontal_tile_25_16_to_tile_25_17_3),
		.in_wire_0_0(horizontal_tile_25_17_to_tile_25_16_0),
		.in_wire_0_1(horizontal_tile_25_17_to_tile_25_16_1),
		.in_wire_0_2(horizontal_tile_25_17_to_tile_25_16_2),
		.in_wire_0_3(horizontal_tile_25_17_to_tile_25_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(817)
	);

	pe_tile pe_tile_25_17(
		.out_wire_3_0(vertical_tile_25_17_to_tile_24_17_0),
		.out_wire_3_1(vertical_tile_25_17_to_tile_24_17_1),
		.out_wire_3_2(vertical_tile_25_17_to_tile_24_17_2),
		.out_wire_3_3(vertical_tile_25_17_to_tile_24_17_3),
		.in_wire_3_0(vertical_tile_24_17_to_tile_25_17_0),
		.in_wire_3_1(vertical_tile_24_17_to_tile_25_17_1),
		.in_wire_3_2(vertical_tile_24_17_to_tile_25_17_2),
		.in_wire_3_3(vertical_tile_24_17_to_tile_25_17_3),
		.out_wire_1_0(vertical_tile_25_17_to_tile_26_17_0),
		.out_wire_1_1(vertical_tile_25_17_to_tile_26_17_1),
		.out_wire_1_2(vertical_tile_25_17_to_tile_26_17_2),
		.out_wire_1_3(vertical_tile_25_17_to_tile_26_17_3),
		.in_wire_1_0(vertical_tile_26_17_to_tile_25_17_0),
		.in_wire_1_1(vertical_tile_26_17_to_tile_25_17_1),
		.in_wire_1_2(vertical_tile_26_17_to_tile_25_17_2),
		.in_wire_1_3(vertical_tile_26_17_to_tile_25_17_3),
		.out_wire_2_0(horizontal_tile_25_17_to_tile_25_16_0),
		.out_wire_2_1(horizontal_tile_25_17_to_tile_25_16_1),
		.out_wire_2_2(horizontal_tile_25_17_to_tile_25_16_2),
		.out_wire_2_3(horizontal_tile_25_17_to_tile_25_16_3),
		.in_wire_2_0(horizontal_tile_25_16_to_tile_25_17_0),
		.in_wire_2_1(horizontal_tile_25_16_to_tile_25_17_1),
		.in_wire_2_2(horizontal_tile_25_16_to_tile_25_17_2),
		.in_wire_2_3(horizontal_tile_25_16_to_tile_25_17_3),
		.out_wire_0_0(horizontal_tile_25_17_to_tile_25_18_0),
		.out_wire_0_1(horizontal_tile_25_17_to_tile_25_18_1),
		.out_wire_0_2(horizontal_tile_25_17_to_tile_25_18_2),
		.out_wire_0_3(horizontal_tile_25_17_to_tile_25_18_3),
		.in_wire_0_0(horizontal_tile_25_18_to_tile_25_17_0),
		.in_wire_0_1(horizontal_tile_25_18_to_tile_25_17_1),
		.in_wire_0_2(horizontal_tile_25_18_to_tile_25_17_2),
		.in_wire_0_3(horizontal_tile_25_18_to_tile_25_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(818)
	);

	pe_tile pe_tile_25_18(
		.out_wire_3_0(vertical_tile_25_18_to_tile_24_18_0),
		.out_wire_3_1(vertical_tile_25_18_to_tile_24_18_1),
		.out_wire_3_2(vertical_tile_25_18_to_tile_24_18_2),
		.out_wire_3_3(vertical_tile_25_18_to_tile_24_18_3),
		.in_wire_3_0(vertical_tile_24_18_to_tile_25_18_0),
		.in_wire_3_1(vertical_tile_24_18_to_tile_25_18_1),
		.in_wire_3_2(vertical_tile_24_18_to_tile_25_18_2),
		.in_wire_3_3(vertical_tile_24_18_to_tile_25_18_3),
		.out_wire_1_0(vertical_tile_25_18_to_tile_26_18_0),
		.out_wire_1_1(vertical_tile_25_18_to_tile_26_18_1),
		.out_wire_1_2(vertical_tile_25_18_to_tile_26_18_2),
		.out_wire_1_3(vertical_tile_25_18_to_tile_26_18_3),
		.in_wire_1_0(vertical_tile_26_18_to_tile_25_18_0),
		.in_wire_1_1(vertical_tile_26_18_to_tile_25_18_1),
		.in_wire_1_2(vertical_tile_26_18_to_tile_25_18_2),
		.in_wire_1_3(vertical_tile_26_18_to_tile_25_18_3),
		.out_wire_2_0(horizontal_tile_25_18_to_tile_25_17_0),
		.out_wire_2_1(horizontal_tile_25_18_to_tile_25_17_1),
		.out_wire_2_2(horizontal_tile_25_18_to_tile_25_17_2),
		.out_wire_2_3(horizontal_tile_25_18_to_tile_25_17_3),
		.in_wire_2_0(horizontal_tile_25_17_to_tile_25_18_0),
		.in_wire_2_1(horizontal_tile_25_17_to_tile_25_18_1),
		.in_wire_2_2(horizontal_tile_25_17_to_tile_25_18_2),
		.in_wire_2_3(horizontal_tile_25_17_to_tile_25_18_3),
		.out_wire_0_0(horizontal_tile_25_18_to_tile_25_19_0),
		.out_wire_0_1(horizontal_tile_25_18_to_tile_25_19_1),
		.out_wire_0_2(horizontal_tile_25_18_to_tile_25_19_2),
		.out_wire_0_3(horizontal_tile_25_18_to_tile_25_19_3),
		.in_wire_0_0(horizontal_tile_25_19_to_tile_25_18_0),
		.in_wire_0_1(horizontal_tile_25_19_to_tile_25_18_1),
		.in_wire_0_2(horizontal_tile_25_19_to_tile_25_18_2),
		.in_wire_0_3(horizontal_tile_25_19_to_tile_25_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(819)
	);

	pe_tile pe_tile_25_19(
		.out_wire_3_0(vertical_tile_25_19_to_tile_24_19_0),
		.out_wire_3_1(vertical_tile_25_19_to_tile_24_19_1),
		.out_wire_3_2(vertical_tile_25_19_to_tile_24_19_2),
		.out_wire_3_3(vertical_tile_25_19_to_tile_24_19_3),
		.in_wire_3_0(vertical_tile_24_19_to_tile_25_19_0),
		.in_wire_3_1(vertical_tile_24_19_to_tile_25_19_1),
		.in_wire_3_2(vertical_tile_24_19_to_tile_25_19_2),
		.in_wire_3_3(vertical_tile_24_19_to_tile_25_19_3),
		.out_wire_1_0(vertical_tile_25_19_to_tile_26_19_0),
		.out_wire_1_1(vertical_tile_25_19_to_tile_26_19_1),
		.out_wire_1_2(vertical_tile_25_19_to_tile_26_19_2),
		.out_wire_1_3(vertical_tile_25_19_to_tile_26_19_3),
		.in_wire_1_0(vertical_tile_26_19_to_tile_25_19_0),
		.in_wire_1_1(vertical_tile_26_19_to_tile_25_19_1),
		.in_wire_1_2(vertical_tile_26_19_to_tile_25_19_2),
		.in_wire_1_3(vertical_tile_26_19_to_tile_25_19_3),
		.out_wire_2_0(horizontal_tile_25_19_to_tile_25_18_0),
		.out_wire_2_1(horizontal_tile_25_19_to_tile_25_18_1),
		.out_wire_2_2(horizontal_tile_25_19_to_tile_25_18_2),
		.out_wire_2_3(horizontal_tile_25_19_to_tile_25_18_3),
		.in_wire_2_0(horizontal_tile_25_18_to_tile_25_19_0),
		.in_wire_2_1(horizontal_tile_25_18_to_tile_25_19_1),
		.in_wire_2_2(horizontal_tile_25_18_to_tile_25_19_2),
		.in_wire_2_3(horizontal_tile_25_18_to_tile_25_19_3),
		.out_wire_0_0(horizontal_tile_25_19_to_tile_25_20_0),
		.out_wire_0_1(horizontal_tile_25_19_to_tile_25_20_1),
		.out_wire_0_2(horizontal_tile_25_19_to_tile_25_20_2),
		.out_wire_0_3(horizontal_tile_25_19_to_tile_25_20_3),
		.in_wire_0_0(horizontal_tile_25_20_to_tile_25_19_0),
		.in_wire_0_1(horizontal_tile_25_20_to_tile_25_19_1),
		.in_wire_0_2(horizontal_tile_25_20_to_tile_25_19_2),
		.in_wire_0_3(horizontal_tile_25_20_to_tile_25_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(820)
	);

	pe_tile pe_tile_25_20(
		.out_wire_3_0(vertical_tile_25_20_to_tile_24_20_0),
		.out_wire_3_1(vertical_tile_25_20_to_tile_24_20_1),
		.out_wire_3_2(vertical_tile_25_20_to_tile_24_20_2),
		.out_wire_3_3(vertical_tile_25_20_to_tile_24_20_3),
		.in_wire_3_0(vertical_tile_24_20_to_tile_25_20_0),
		.in_wire_3_1(vertical_tile_24_20_to_tile_25_20_1),
		.in_wire_3_2(vertical_tile_24_20_to_tile_25_20_2),
		.in_wire_3_3(vertical_tile_24_20_to_tile_25_20_3),
		.out_wire_1_0(vertical_tile_25_20_to_tile_26_20_0),
		.out_wire_1_1(vertical_tile_25_20_to_tile_26_20_1),
		.out_wire_1_2(vertical_tile_25_20_to_tile_26_20_2),
		.out_wire_1_3(vertical_tile_25_20_to_tile_26_20_3),
		.in_wire_1_0(vertical_tile_26_20_to_tile_25_20_0),
		.in_wire_1_1(vertical_tile_26_20_to_tile_25_20_1),
		.in_wire_1_2(vertical_tile_26_20_to_tile_25_20_2),
		.in_wire_1_3(vertical_tile_26_20_to_tile_25_20_3),
		.out_wire_2_0(horizontal_tile_25_20_to_tile_25_19_0),
		.out_wire_2_1(horizontal_tile_25_20_to_tile_25_19_1),
		.out_wire_2_2(horizontal_tile_25_20_to_tile_25_19_2),
		.out_wire_2_3(horizontal_tile_25_20_to_tile_25_19_3),
		.in_wire_2_0(horizontal_tile_25_19_to_tile_25_20_0),
		.in_wire_2_1(horizontal_tile_25_19_to_tile_25_20_1),
		.in_wire_2_2(horizontal_tile_25_19_to_tile_25_20_2),
		.in_wire_2_3(horizontal_tile_25_19_to_tile_25_20_3),
		.out_wire_0_0(horizontal_tile_25_20_to_tile_25_21_0),
		.out_wire_0_1(horizontal_tile_25_20_to_tile_25_21_1),
		.out_wire_0_2(horizontal_tile_25_20_to_tile_25_21_2),
		.out_wire_0_3(horizontal_tile_25_20_to_tile_25_21_3),
		.in_wire_0_0(horizontal_tile_25_21_to_tile_25_20_0),
		.in_wire_0_1(horizontal_tile_25_21_to_tile_25_20_1),
		.in_wire_0_2(horizontal_tile_25_21_to_tile_25_20_2),
		.in_wire_0_3(horizontal_tile_25_21_to_tile_25_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(821)
	);

	pe_tile pe_tile_25_21(
		.out_wire_3_0(vertical_tile_25_21_to_tile_24_21_0),
		.out_wire_3_1(vertical_tile_25_21_to_tile_24_21_1),
		.out_wire_3_2(vertical_tile_25_21_to_tile_24_21_2),
		.out_wire_3_3(vertical_tile_25_21_to_tile_24_21_3),
		.in_wire_3_0(vertical_tile_24_21_to_tile_25_21_0),
		.in_wire_3_1(vertical_tile_24_21_to_tile_25_21_1),
		.in_wire_3_2(vertical_tile_24_21_to_tile_25_21_2),
		.in_wire_3_3(vertical_tile_24_21_to_tile_25_21_3),
		.out_wire_1_0(vertical_tile_25_21_to_tile_26_21_0),
		.out_wire_1_1(vertical_tile_25_21_to_tile_26_21_1),
		.out_wire_1_2(vertical_tile_25_21_to_tile_26_21_2),
		.out_wire_1_3(vertical_tile_25_21_to_tile_26_21_3),
		.in_wire_1_0(vertical_tile_26_21_to_tile_25_21_0),
		.in_wire_1_1(vertical_tile_26_21_to_tile_25_21_1),
		.in_wire_1_2(vertical_tile_26_21_to_tile_25_21_2),
		.in_wire_1_3(vertical_tile_26_21_to_tile_25_21_3),
		.out_wire_2_0(horizontal_tile_25_21_to_tile_25_20_0),
		.out_wire_2_1(horizontal_tile_25_21_to_tile_25_20_1),
		.out_wire_2_2(horizontal_tile_25_21_to_tile_25_20_2),
		.out_wire_2_3(horizontal_tile_25_21_to_tile_25_20_3),
		.in_wire_2_0(horizontal_tile_25_20_to_tile_25_21_0),
		.in_wire_2_1(horizontal_tile_25_20_to_tile_25_21_1),
		.in_wire_2_2(horizontal_tile_25_20_to_tile_25_21_2),
		.in_wire_2_3(horizontal_tile_25_20_to_tile_25_21_3),
		.out_wire_0_0(horizontal_tile_25_21_to_tile_25_22_0),
		.out_wire_0_1(horizontal_tile_25_21_to_tile_25_22_1),
		.out_wire_0_2(horizontal_tile_25_21_to_tile_25_22_2),
		.out_wire_0_3(horizontal_tile_25_21_to_tile_25_22_3),
		.in_wire_0_0(horizontal_tile_25_22_to_tile_25_21_0),
		.in_wire_0_1(horizontal_tile_25_22_to_tile_25_21_1),
		.in_wire_0_2(horizontal_tile_25_22_to_tile_25_21_2),
		.in_wire_0_3(horizontal_tile_25_22_to_tile_25_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(822)
	);

	pe_tile pe_tile_25_22(
		.out_wire_3_0(vertical_tile_25_22_to_tile_24_22_0),
		.out_wire_3_1(vertical_tile_25_22_to_tile_24_22_1),
		.out_wire_3_2(vertical_tile_25_22_to_tile_24_22_2),
		.out_wire_3_3(vertical_tile_25_22_to_tile_24_22_3),
		.in_wire_3_0(vertical_tile_24_22_to_tile_25_22_0),
		.in_wire_3_1(vertical_tile_24_22_to_tile_25_22_1),
		.in_wire_3_2(vertical_tile_24_22_to_tile_25_22_2),
		.in_wire_3_3(vertical_tile_24_22_to_tile_25_22_3),
		.out_wire_1_0(vertical_tile_25_22_to_tile_26_22_0),
		.out_wire_1_1(vertical_tile_25_22_to_tile_26_22_1),
		.out_wire_1_2(vertical_tile_25_22_to_tile_26_22_2),
		.out_wire_1_3(vertical_tile_25_22_to_tile_26_22_3),
		.in_wire_1_0(vertical_tile_26_22_to_tile_25_22_0),
		.in_wire_1_1(vertical_tile_26_22_to_tile_25_22_1),
		.in_wire_1_2(vertical_tile_26_22_to_tile_25_22_2),
		.in_wire_1_3(vertical_tile_26_22_to_tile_25_22_3),
		.out_wire_2_0(horizontal_tile_25_22_to_tile_25_21_0),
		.out_wire_2_1(horizontal_tile_25_22_to_tile_25_21_1),
		.out_wire_2_2(horizontal_tile_25_22_to_tile_25_21_2),
		.out_wire_2_3(horizontal_tile_25_22_to_tile_25_21_3),
		.in_wire_2_0(horizontal_tile_25_21_to_tile_25_22_0),
		.in_wire_2_1(horizontal_tile_25_21_to_tile_25_22_1),
		.in_wire_2_2(horizontal_tile_25_21_to_tile_25_22_2),
		.in_wire_2_3(horizontal_tile_25_21_to_tile_25_22_3),
		.out_wire_0_0(horizontal_tile_25_22_to_tile_25_23_0),
		.out_wire_0_1(horizontal_tile_25_22_to_tile_25_23_1),
		.out_wire_0_2(horizontal_tile_25_22_to_tile_25_23_2),
		.out_wire_0_3(horizontal_tile_25_22_to_tile_25_23_3),
		.in_wire_0_0(horizontal_tile_25_23_to_tile_25_22_0),
		.in_wire_0_1(horizontal_tile_25_23_to_tile_25_22_1),
		.in_wire_0_2(horizontal_tile_25_23_to_tile_25_22_2),
		.in_wire_0_3(horizontal_tile_25_23_to_tile_25_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(823)
	);

	pe_tile pe_tile_25_23(
		.out_wire_3_0(vertical_tile_25_23_to_tile_24_23_0),
		.out_wire_3_1(vertical_tile_25_23_to_tile_24_23_1),
		.out_wire_3_2(vertical_tile_25_23_to_tile_24_23_2),
		.out_wire_3_3(vertical_tile_25_23_to_tile_24_23_3),
		.in_wire_3_0(vertical_tile_24_23_to_tile_25_23_0),
		.in_wire_3_1(vertical_tile_24_23_to_tile_25_23_1),
		.in_wire_3_2(vertical_tile_24_23_to_tile_25_23_2),
		.in_wire_3_3(vertical_tile_24_23_to_tile_25_23_3),
		.out_wire_1_0(vertical_tile_25_23_to_tile_26_23_0),
		.out_wire_1_1(vertical_tile_25_23_to_tile_26_23_1),
		.out_wire_1_2(vertical_tile_25_23_to_tile_26_23_2),
		.out_wire_1_3(vertical_tile_25_23_to_tile_26_23_3),
		.in_wire_1_0(vertical_tile_26_23_to_tile_25_23_0),
		.in_wire_1_1(vertical_tile_26_23_to_tile_25_23_1),
		.in_wire_1_2(vertical_tile_26_23_to_tile_25_23_2),
		.in_wire_1_3(vertical_tile_26_23_to_tile_25_23_3),
		.out_wire_2_0(horizontal_tile_25_23_to_tile_25_22_0),
		.out_wire_2_1(horizontal_tile_25_23_to_tile_25_22_1),
		.out_wire_2_2(horizontal_tile_25_23_to_tile_25_22_2),
		.out_wire_2_3(horizontal_tile_25_23_to_tile_25_22_3),
		.in_wire_2_0(horizontal_tile_25_22_to_tile_25_23_0),
		.in_wire_2_1(horizontal_tile_25_22_to_tile_25_23_1),
		.in_wire_2_2(horizontal_tile_25_22_to_tile_25_23_2),
		.in_wire_2_3(horizontal_tile_25_22_to_tile_25_23_3),
		.out_wire_0_0(horizontal_tile_25_23_to_tile_25_24_0),
		.out_wire_0_1(horizontal_tile_25_23_to_tile_25_24_1),
		.out_wire_0_2(horizontal_tile_25_23_to_tile_25_24_2),
		.out_wire_0_3(horizontal_tile_25_23_to_tile_25_24_3),
		.in_wire_0_0(horizontal_tile_25_24_to_tile_25_23_0),
		.in_wire_0_1(horizontal_tile_25_24_to_tile_25_23_1),
		.in_wire_0_2(horizontal_tile_25_24_to_tile_25_23_2),
		.in_wire_0_3(horizontal_tile_25_24_to_tile_25_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(824)
	);

	pe_tile pe_tile_25_24(
		.out_wire_3_0(vertical_tile_25_24_to_tile_24_24_0),
		.out_wire_3_1(vertical_tile_25_24_to_tile_24_24_1),
		.out_wire_3_2(vertical_tile_25_24_to_tile_24_24_2),
		.out_wire_3_3(vertical_tile_25_24_to_tile_24_24_3),
		.in_wire_3_0(vertical_tile_24_24_to_tile_25_24_0),
		.in_wire_3_1(vertical_tile_24_24_to_tile_25_24_1),
		.in_wire_3_2(vertical_tile_24_24_to_tile_25_24_2),
		.in_wire_3_3(vertical_tile_24_24_to_tile_25_24_3),
		.out_wire_1_0(vertical_tile_25_24_to_tile_26_24_0),
		.out_wire_1_1(vertical_tile_25_24_to_tile_26_24_1),
		.out_wire_1_2(vertical_tile_25_24_to_tile_26_24_2),
		.out_wire_1_3(vertical_tile_25_24_to_tile_26_24_3),
		.in_wire_1_0(vertical_tile_26_24_to_tile_25_24_0),
		.in_wire_1_1(vertical_tile_26_24_to_tile_25_24_1),
		.in_wire_1_2(vertical_tile_26_24_to_tile_25_24_2),
		.in_wire_1_3(vertical_tile_26_24_to_tile_25_24_3),
		.out_wire_2_0(horizontal_tile_25_24_to_tile_25_23_0),
		.out_wire_2_1(horizontal_tile_25_24_to_tile_25_23_1),
		.out_wire_2_2(horizontal_tile_25_24_to_tile_25_23_2),
		.out_wire_2_3(horizontal_tile_25_24_to_tile_25_23_3),
		.in_wire_2_0(horizontal_tile_25_23_to_tile_25_24_0),
		.in_wire_2_1(horizontal_tile_25_23_to_tile_25_24_1),
		.in_wire_2_2(horizontal_tile_25_23_to_tile_25_24_2),
		.in_wire_2_3(horizontal_tile_25_23_to_tile_25_24_3),
		.out_wire_0_0(horizontal_tile_25_24_to_tile_25_25_0),
		.out_wire_0_1(horizontal_tile_25_24_to_tile_25_25_1),
		.out_wire_0_2(horizontal_tile_25_24_to_tile_25_25_2),
		.out_wire_0_3(horizontal_tile_25_24_to_tile_25_25_3),
		.in_wire_0_0(horizontal_tile_25_25_to_tile_25_24_0),
		.in_wire_0_1(horizontal_tile_25_25_to_tile_25_24_1),
		.in_wire_0_2(horizontal_tile_25_25_to_tile_25_24_2),
		.in_wire_0_3(horizontal_tile_25_25_to_tile_25_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(825)
	);

	pe_tile pe_tile_25_25(
		.out_wire_3_0(vertical_tile_25_25_to_tile_24_25_0),
		.out_wire_3_1(vertical_tile_25_25_to_tile_24_25_1),
		.out_wire_3_2(vertical_tile_25_25_to_tile_24_25_2),
		.out_wire_3_3(vertical_tile_25_25_to_tile_24_25_3),
		.in_wire_3_0(vertical_tile_24_25_to_tile_25_25_0),
		.in_wire_3_1(vertical_tile_24_25_to_tile_25_25_1),
		.in_wire_3_2(vertical_tile_24_25_to_tile_25_25_2),
		.in_wire_3_3(vertical_tile_24_25_to_tile_25_25_3),
		.out_wire_1_0(vertical_tile_25_25_to_tile_26_25_0),
		.out_wire_1_1(vertical_tile_25_25_to_tile_26_25_1),
		.out_wire_1_2(vertical_tile_25_25_to_tile_26_25_2),
		.out_wire_1_3(vertical_tile_25_25_to_tile_26_25_3),
		.in_wire_1_0(vertical_tile_26_25_to_tile_25_25_0),
		.in_wire_1_1(vertical_tile_26_25_to_tile_25_25_1),
		.in_wire_1_2(vertical_tile_26_25_to_tile_25_25_2),
		.in_wire_1_3(vertical_tile_26_25_to_tile_25_25_3),
		.out_wire_2_0(horizontal_tile_25_25_to_tile_25_24_0),
		.out_wire_2_1(horizontal_tile_25_25_to_tile_25_24_1),
		.out_wire_2_2(horizontal_tile_25_25_to_tile_25_24_2),
		.out_wire_2_3(horizontal_tile_25_25_to_tile_25_24_3),
		.in_wire_2_0(horizontal_tile_25_24_to_tile_25_25_0),
		.in_wire_2_1(horizontal_tile_25_24_to_tile_25_25_1),
		.in_wire_2_2(horizontal_tile_25_24_to_tile_25_25_2),
		.in_wire_2_3(horizontal_tile_25_24_to_tile_25_25_3),
		.out_wire_0_0(horizontal_tile_25_25_to_tile_25_26_0),
		.out_wire_0_1(horizontal_tile_25_25_to_tile_25_26_1),
		.out_wire_0_2(horizontal_tile_25_25_to_tile_25_26_2),
		.out_wire_0_3(horizontal_tile_25_25_to_tile_25_26_3),
		.in_wire_0_0(horizontal_tile_25_26_to_tile_25_25_0),
		.in_wire_0_1(horizontal_tile_25_26_to_tile_25_25_1),
		.in_wire_0_2(horizontal_tile_25_26_to_tile_25_25_2),
		.in_wire_0_3(horizontal_tile_25_26_to_tile_25_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(826)
	);

	pe_tile pe_tile_25_26(
		.out_wire_3_0(vertical_tile_25_26_to_tile_24_26_0),
		.out_wire_3_1(vertical_tile_25_26_to_tile_24_26_1),
		.out_wire_3_2(vertical_tile_25_26_to_tile_24_26_2),
		.out_wire_3_3(vertical_tile_25_26_to_tile_24_26_3),
		.in_wire_3_0(vertical_tile_24_26_to_tile_25_26_0),
		.in_wire_3_1(vertical_tile_24_26_to_tile_25_26_1),
		.in_wire_3_2(vertical_tile_24_26_to_tile_25_26_2),
		.in_wire_3_3(vertical_tile_24_26_to_tile_25_26_3),
		.out_wire_1_0(vertical_tile_25_26_to_tile_26_26_0),
		.out_wire_1_1(vertical_tile_25_26_to_tile_26_26_1),
		.out_wire_1_2(vertical_tile_25_26_to_tile_26_26_2),
		.out_wire_1_3(vertical_tile_25_26_to_tile_26_26_3),
		.in_wire_1_0(vertical_tile_26_26_to_tile_25_26_0),
		.in_wire_1_1(vertical_tile_26_26_to_tile_25_26_1),
		.in_wire_1_2(vertical_tile_26_26_to_tile_25_26_2),
		.in_wire_1_3(vertical_tile_26_26_to_tile_25_26_3),
		.out_wire_2_0(horizontal_tile_25_26_to_tile_25_25_0),
		.out_wire_2_1(horizontal_tile_25_26_to_tile_25_25_1),
		.out_wire_2_2(horizontal_tile_25_26_to_tile_25_25_2),
		.out_wire_2_3(horizontal_tile_25_26_to_tile_25_25_3),
		.in_wire_2_0(horizontal_tile_25_25_to_tile_25_26_0),
		.in_wire_2_1(horizontal_tile_25_25_to_tile_25_26_1),
		.in_wire_2_2(horizontal_tile_25_25_to_tile_25_26_2),
		.in_wire_2_3(horizontal_tile_25_25_to_tile_25_26_3),
		.out_wire_0_0(horizontal_tile_25_26_to_tile_25_27_0),
		.out_wire_0_1(horizontal_tile_25_26_to_tile_25_27_1),
		.out_wire_0_2(horizontal_tile_25_26_to_tile_25_27_2),
		.out_wire_0_3(horizontal_tile_25_26_to_tile_25_27_3),
		.in_wire_0_0(horizontal_tile_25_27_to_tile_25_26_0),
		.in_wire_0_1(horizontal_tile_25_27_to_tile_25_26_1),
		.in_wire_0_2(horizontal_tile_25_27_to_tile_25_26_2),
		.in_wire_0_3(horizontal_tile_25_27_to_tile_25_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(827)
	);

	pe_tile pe_tile_25_27(
		.out_wire_3_0(vertical_tile_25_27_to_tile_24_27_0),
		.out_wire_3_1(vertical_tile_25_27_to_tile_24_27_1),
		.out_wire_3_2(vertical_tile_25_27_to_tile_24_27_2),
		.out_wire_3_3(vertical_tile_25_27_to_tile_24_27_3),
		.in_wire_3_0(vertical_tile_24_27_to_tile_25_27_0),
		.in_wire_3_1(vertical_tile_24_27_to_tile_25_27_1),
		.in_wire_3_2(vertical_tile_24_27_to_tile_25_27_2),
		.in_wire_3_3(vertical_tile_24_27_to_tile_25_27_3),
		.out_wire_1_0(vertical_tile_25_27_to_tile_26_27_0),
		.out_wire_1_1(vertical_tile_25_27_to_tile_26_27_1),
		.out_wire_1_2(vertical_tile_25_27_to_tile_26_27_2),
		.out_wire_1_3(vertical_tile_25_27_to_tile_26_27_3),
		.in_wire_1_0(vertical_tile_26_27_to_tile_25_27_0),
		.in_wire_1_1(vertical_tile_26_27_to_tile_25_27_1),
		.in_wire_1_2(vertical_tile_26_27_to_tile_25_27_2),
		.in_wire_1_3(vertical_tile_26_27_to_tile_25_27_3),
		.out_wire_2_0(horizontal_tile_25_27_to_tile_25_26_0),
		.out_wire_2_1(horizontal_tile_25_27_to_tile_25_26_1),
		.out_wire_2_2(horizontal_tile_25_27_to_tile_25_26_2),
		.out_wire_2_3(horizontal_tile_25_27_to_tile_25_26_3),
		.in_wire_2_0(horizontal_tile_25_26_to_tile_25_27_0),
		.in_wire_2_1(horizontal_tile_25_26_to_tile_25_27_1),
		.in_wire_2_2(horizontal_tile_25_26_to_tile_25_27_2),
		.in_wire_2_3(horizontal_tile_25_26_to_tile_25_27_3),
		.out_wire_0_0(horizontal_tile_25_27_to_tile_25_28_0),
		.out_wire_0_1(horizontal_tile_25_27_to_tile_25_28_1),
		.out_wire_0_2(horizontal_tile_25_27_to_tile_25_28_2),
		.out_wire_0_3(horizontal_tile_25_27_to_tile_25_28_3),
		.in_wire_0_0(horizontal_tile_25_28_to_tile_25_27_0),
		.in_wire_0_1(horizontal_tile_25_28_to_tile_25_27_1),
		.in_wire_0_2(horizontal_tile_25_28_to_tile_25_27_2),
		.in_wire_0_3(horizontal_tile_25_28_to_tile_25_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(828)
	);

	pe_tile pe_tile_25_28(
		.out_wire_3_0(vertical_tile_25_28_to_tile_24_28_0),
		.out_wire_3_1(vertical_tile_25_28_to_tile_24_28_1),
		.out_wire_3_2(vertical_tile_25_28_to_tile_24_28_2),
		.out_wire_3_3(vertical_tile_25_28_to_tile_24_28_3),
		.in_wire_3_0(vertical_tile_24_28_to_tile_25_28_0),
		.in_wire_3_1(vertical_tile_24_28_to_tile_25_28_1),
		.in_wire_3_2(vertical_tile_24_28_to_tile_25_28_2),
		.in_wire_3_3(vertical_tile_24_28_to_tile_25_28_3),
		.out_wire_1_0(vertical_tile_25_28_to_tile_26_28_0),
		.out_wire_1_1(vertical_tile_25_28_to_tile_26_28_1),
		.out_wire_1_2(vertical_tile_25_28_to_tile_26_28_2),
		.out_wire_1_3(vertical_tile_25_28_to_tile_26_28_3),
		.in_wire_1_0(vertical_tile_26_28_to_tile_25_28_0),
		.in_wire_1_1(vertical_tile_26_28_to_tile_25_28_1),
		.in_wire_1_2(vertical_tile_26_28_to_tile_25_28_2),
		.in_wire_1_3(vertical_tile_26_28_to_tile_25_28_3),
		.out_wire_2_0(horizontal_tile_25_28_to_tile_25_27_0),
		.out_wire_2_1(horizontal_tile_25_28_to_tile_25_27_1),
		.out_wire_2_2(horizontal_tile_25_28_to_tile_25_27_2),
		.out_wire_2_3(horizontal_tile_25_28_to_tile_25_27_3),
		.in_wire_2_0(horizontal_tile_25_27_to_tile_25_28_0),
		.in_wire_2_1(horizontal_tile_25_27_to_tile_25_28_1),
		.in_wire_2_2(horizontal_tile_25_27_to_tile_25_28_2),
		.in_wire_2_3(horizontal_tile_25_27_to_tile_25_28_3),
		.out_wire_0_0(horizontal_tile_25_28_to_tile_25_29_0),
		.out_wire_0_1(horizontal_tile_25_28_to_tile_25_29_1),
		.out_wire_0_2(horizontal_tile_25_28_to_tile_25_29_2),
		.out_wire_0_3(horizontal_tile_25_28_to_tile_25_29_3),
		.in_wire_0_0(horizontal_tile_25_29_to_tile_25_28_0),
		.in_wire_0_1(horizontal_tile_25_29_to_tile_25_28_1),
		.in_wire_0_2(horizontal_tile_25_29_to_tile_25_28_2),
		.in_wire_0_3(horizontal_tile_25_29_to_tile_25_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(829)
	);

	pe_tile pe_tile_25_29(
		.out_wire_3_0(vertical_tile_25_29_to_tile_24_29_0),
		.out_wire_3_1(vertical_tile_25_29_to_tile_24_29_1),
		.out_wire_3_2(vertical_tile_25_29_to_tile_24_29_2),
		.out_wire_3_3(vertical_tile_25_29_to_tile_24_29_3),
		.in_wire_3_0(vertical_tile_24_29_to_tile_25_29_0),
		.in_wire_3_1(vertical_tile_24_29_to_tile_25_29_1),
		.in_wire_3_2(vertical_tile_24_29_to_tile_25_29_2),
		.in_wire_3_3(vertical_tile_24_29_to_tile_25_29_3),
		.out_wire_1_0(vertical_tile_25_29_to_tile_26_29_0),
		.out_wire_1_1(vertical_tile_25_29_to_tile_26_29_1),
		.out_wire_1_2(vertical_tile_25_29_to_tile_26_29_2),
		.out_wire_1_3(vertical_tile_25_29_to_tile_26_29_3),
		.in_wire_1_0(vertical_tile_26_29_to_tile_25_29_0),
		.in_wire_1_1(vertical_tile_26_29_to_tile_25_29_1),
		.in_wire_1_2(vertical_tile_26_29_to_tile_25_29_2),
		.in_wire_1_3(vertical_tile_26_29_to_tile_25_29_3),
		.out_wire_2_0(horizontal_tile_25_29_to_tile_25_28_0),
		.out_wire_2_1(horizontal_tile_25_29_to_tile_25_28_1),
		.out_wire_2_2(horizontal_tile_25_29_to_tile_25_28_2),
		.out_wire_2_3(horizontal_tile_25_29_to_tile_25_28_3),
		.in_wire_2_0(horizontal_tile_25_28_to_tile_25_29_0),
		.in_wire_2_1(horizontal_tile_25_28_to_tile_25_29_1),
		.in_wire_2_2(horizontal_tile_25_28_to_tile_25_29_2),
		.in_wire_2_3(horizontal_tile_25_28_to_tile_25_29_3),
		.out_wire_0_0(horizontal_tile_25_29_to_tile_25_30_0),
		.out_wire_0_1(horizontal_tile_25_29_to_tile_25_30_1),
		.out_wire_0_2(horizontal_tile_25_29_to_tile_25_30_2),
		.out_wire_0_3(horizontal_tile_25_29_to_tile_25_30_3),
		.in_wire_0_0(horizontal_tile_25_30_to_tile_25_29_0),
		.in_wire_0_1(horizontal_tile_25_30_to_tile_25_29_1),
		.in_wire_0_2(horizontal_tile_25_30_to_tile_25_29_2),
		.in_wire_0_3(horizontal_tile_25_30_to_tile_25_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(830)
	);

	pe_tile pe_tile_25_30(
		.out_wire_3_0(vertical_tile_25_30_to_tile_24_30_0),
		.out_wire_3_1(vertical_tile_25_30_to_tile_24_30_1),
		.out_wire_3_2(vertical_tile_25_30_to_tile_24_30_2),
		.out_wire_3_3(vertical_tile_25_30_to_tile_24_30_3),
		.in_wire_3_0(vertical_tile_24_30_to_tile_25_30_0),
		.in_wire_3_1(vertical_tile_24_30_to_tile_25_30_1),
		.in_wire_3_2(vertical_tile_24_30_to_tile_25_30_2),
		.in_wire_3_3(vertical_tile_24_30_to_tile_25_30_3),
		.out_wire_1_0(vertical_tile_25_30_to_tile_26_30_0),
		.out_wire_1_1(vertical_tile_25_30_to_tile_26_30_1),
		.out_wire_1_2(vertical_tile_25_30_to_tile_26_30_2),
		.out_wire_1_3(vertical_tile_25_30_to_tile_26_30_3),
		.in_wire_1_0(vertical_tile_26_30_to_tile_25_30_0),
		.in_wire_1_1(vertical_tile_26_30_to_tile_25_30_1),
		.in_wire_1_2(vertical_tile_26_30_to_tile_25_30_2),
		.in_wire_1_3(vertical_tile_26_30_to_tile_25_30_3),
		.out_wire_2_0(horizontal_tile_25_30_to_tile_25_29_0),
		.out_wire_2_1(horizontal_tile_25_30_to_tile_25_29_1),
		.out_wire_2_2(horizontal_tile_25_30_to_tile_25_29_2),
		.out_wire_2_3(horizontal_tile_25_30_to_tile_25_29_3),
		.in_wire_2_0(horizontal_tile_25_29_to_tile_25_30_0),
		.in_wire_2_1(horizontal_tile_25_29_to_tile_25_30_1),
		.in_wire_2_2(horizontal_tile_25_29_to_tile_25_30_2),
		.in_wire_2_3(horizontal_tile_25_29_to_tile_25_30_3),
		.out_wire_0_0(horizontal_tile_25_30_to_tile_25_31_0),
		.out_wire_0_1(horizontal_tile_25_30_to_tile_25_31_1),
		.out_wire_0_2(horizontal_tile_25_30_to_tile_25_31_2),
		.out_wire_0_3(horizontal_tile_25_30_to_tile_25_31_3),
		.in_wire_0_0(horizontal_tile_25_31_to_tile_25_30_0),
		.in_wire_0_1(horizontal_tile_25_31_to_tile_25_30_1),
		.in_wire_0_2(horizontal_tile_25_31_to_tile_25_30_2),
		.in_wire_0_3(horizontal_tile_25_31_to_tile_25_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(831)
	);

	pe_tile_right pe_tile_25_31(
		.out_wire_3_0(vertical_tile_25_31_to_tile_24_31_0),
		.out_wire_3_1(vertical_tile_25_31_to_tile_24_31_1),
		.out_wire_3_2(vertical_tile_25_31_to_tile_24_31_2),
		.out_wire_3_3(vertical_tile_25_31_to_tile_24_31_3),
		.in_wire_3_0(vertical_tile_24_31_to_tile_25_31_0),
		.in_wire_3_1(vertical_tile_24_31_to_tile_25_31_1),
		.in_wire_3_2(vertical_tile_24_31_to_tile_25_31_2),
		.in_wire_3_3(vertical_tile_24_31_to_tile_25_31_3),
		.out_wire_1_0(vertical_tile_25_31_to_tile_26_31_0),
		.out_wire_1_1(vertical_tile_25_31_to_tile_26_31_1),
		.out_wire_1_2(vertical_tile_25_31_to_tile_26_31_2),
		.out_wire_1_3(vertical_tile_25_31_to_tile_26_31_3),
		.in_wire_1_0(vertical_tile_26_31_to_tile_25_31_0),
		.in_wire_1_1(vertical_tile_26_31_to_tile_25_31_1),
		.in_wire_1_2(vertical_tile_26_31_to_tile_25_31_2),
		.in_wire_1_3(vertical_tile_26_31_to_tile_25_31_3),
		.out_wire_2_0(horizontal_tile_25_31_to_tile_25_30_0),
		.out_wire_2_1(horizontal_tile_25_31_to_tile_25_30_1),
		.out_wire_2_2(horizontal_tile_25_31_to_tile_25_30_2),
		.out_wire_2_3(horizontal_tile_25_31_to_tile_25_30_3),
		.in_wire_2_0(horizontal_tile_25_30_to_tile_25_31_0),
		.in_wire_2_1(horizontal_tile_25_30_to_tile_25_31_1),
		.in_wire_2_2(horizontal_tile_25_30_to_tile_25_31_2),
		.in_wire_2_3(horizontal_tile_25_30_to_tile_25_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(832)
	);

	pe_tile_left pe_tile_26_0(
		.out_wire_3_0(vertical_tile_26_0_to_tile_25_0_0),
		.out_wire_3_1(vertical_tile_26_0_to_tile_25_0_1),
		.out_wire_3_2(vertical_tile_26_0_to_tile_25_0_2),
		.out_wire_3_3(vertical_tile_26_0_to_tile_25_0_3),
		.in_wire_3_0(vertical_tile_25_0_to_tile_26_0_0),
		.in_wire_3_1(vertical_tile_25_0_to_tile_26_0_1),
		.in_wire_3_2(vertical_tile_25_0_to_tile_26_0_2),
		.in_wire_3_3(vertical_tile_25_0_to_tile_26_0_3),
		.out_wire_1_0(vertical_tile_26_0_to_tile_27_0_0),
		.out_wire_1_1(vertical_tile_26_0_to_tile_27_0_1),
		.out_wire_1_2(vertical_tile_26_0_to_tile_27_0_2),
		.out_wire_1_3(vertical_tile_26_0_to_tile_27_0_3),
		.in_wire_1_0(vertical_tile_27_0_to_tile_26_0_0),
		.in_wire_1_1(vertical_tile_27_0_to_tile_26_0_1),
		.in_wire_1_2(vertical_tile_27_0_to_tile_26_0_2),
		.in_wire_1_3(vertical_tile_27_0_to_tile_26_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_26_0_to_tile_26_1_0),
		.out_wire_0_1(horizontal_tile_26_0_to_tile_26_1_1),
		.out_wire_0_2(horizontal_tile_26_0_to_tile_26_1_2),
		.out_wire_0_3(horizontal_tile_26_0_to_tile_26_1_3),
		.in_wire_0_0(horizontal_tile_26_1_to_tile_26_0_0),
		.in_wire_0_1(horizontal_tile_26_1_to_tile_26_0_1),
		.in_wire_0_2(horizontal_tile_26_1_to_tile_26_0_2),
		.in_wire_0_3(horizontal_tile_26_1_to_tile_26_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(833)
	);

	pe_tile pe_tile_26_1(
		.out_wire_3_0(vertical_tile_26_1_to_tile_25_1_0),
		.out_wire_3_1(vertical_tile_26_1_to_tile_25_1_1),
		.out_wire_3_2(vertical_tile_26_1_to_tile_25_1_2),
		.out_wire_3_3(vertical_tile_26_1_to_tile_25_1_3),
		.in_wire_3_0(vertical_tile_25_1_to_tile_26_1_0),
		.in_wire_3_1(vertical_tile_25_1_to_tile_26_1_1),
		.in_wire_3_2(vertical_tile_25_1_to_tile_26_1_2),
		.in_wire_3_3(vertical_tile_25_1_to_tile_26_1_3),
		.out_wire_1_0(vertical_tile_26_1_to_tile_27_1_0),
		.out_wire_1_1(vertical_tile_26_1_to_tile_27_1_1),
		.out_wire_1_2(vertical_tile_26_1_to_tile_27_1_2),
		.out_wire_1_3(vertical_tile_26_1_to_tile_27_1_3),
		.in_wire_1_0(vertical_tile_27_1_to_tile_26_1_0),
		.in_wire_1_1(vertical_tile_27_1_to_tile_26_1_1),
		.in_wire_1_2(vertical_tile_27_1_to_tile_26_1_2),
		.in_wire_1_3(vertical_tile_27_1_to_tile_26_1_3),
		.out_wire_2_0(horizontal_tile_26_1_to_tile_26_0_0),
		.out_wire_2_1(horizontal_tile_26_1_to_tile_26_0_1),
		.out_wire_2_2(horizontal_tile_26_1_to_tile_26_0_2),
		.out_wire_2_3(horizontal_tile_26_1_to_tile_26_0_3),
		.in_wire_2_0(horizontal_tile_26_0_to_tile_26_1_0),
		.in_wire_2_1(horizontal_tile_26_0_to_tile_26_1_1),
		.in_wire_2_2(horizontal_tile_26_0_to_tile_26_1_2),
		.in_wire_2_3(horizontal_tile_26_0_to_tile_26_1_3),
		.out_wire_0_0(horizontal_tile_26_1_to_tile_26_2_0),
		.out_wire_0_1(horizontal_tile_26_1_to_tile_26_2_1),
		.out_wire_0_2(horizontal_tile_26_1_to_tile_26_2_2),
		.out_wire_0_3(horizontal_tile_26_1_to_tile_26_2_3),
		.in_wire_0_0(horizontal_tile_26_2_to_tile_26_1_0),
		.in_wire_0_1(horizontal_tile_26_2_to_tile_26_1_1),
		.in_wire_0_2(horizontal_tile_26_2_to_tile_26_1_2),
		.in_wire_0_3(horizontal_tile_26_2_to_tile_26_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(834)
	);

	pe_tile pe_tile_26_2(
		.out_wire_3_0(vertical_tile_26_2_to_tile_25_2_0),
		.out_wire_3_1(vertical_tile_26_2_to_tile_25_2_1),
		.out_wire_3_2(vertical_tile_26_2_to_tile_25_2_2),
		.out_wire_3_3(vertical_tile_26_2_to_tile_25_2_3),
		.in_wire_3_0(vertical_tile_25_2_to_tile_26_2_0),
		.in_wire_3_1(vertical_tile_25_2_to_tile_26_2_1),
		.in_wire_3_2(vertical_tile_25_2_to_tile_26_2_2),
		.in_wire_3_3(vertical_tile_25_2_to_tile_26_2_3),
		.out_wire_1_0(vertical_tile_26_2_to_tile_27_2_0),
		.out_wire_1_1(vertical_tile_26_2_to_tile_27_2_1),
		.out_wire_1_2(vertical_tile_26_2_to_tile_27_2_2),
		.out_wire_1_3(vertical_tile_26_2_to_tile_27_2_3),
		.in_wire_1_0(vertical_tile_27_2_to_tile_26_2_0),
		.in_wire_1_1(vertical_tile_27_2_to_tile_26_2_1),
		.in_wire_1_2(vertical_tile_27_2_to_tile_26_2_2),
		.in_wire_1_3(vertical_tile_27_2_to_tile_26_2_3),
		.out_wire_2_0(horizontal_tile_26_2_to_tile_26_1_0),
		.out_wire_2_1(horizontal_tile_26_2_to_tile_26_1_1),
		.out_wire_2_2(horizontal_tile_26_2_to_tile_26_1_2),
		.out_wire_2_3(horizontal_tile_26_2_to_tile_26_1_3),
		.in_wire_2_0(horizontal_tile_26_1_to_tile_26_2_0),
		.in_wire_2_1(horizontal_tile_26_1_to_tile_26_2_1),
		.in_wire_2_2(horizontal_tile_26_1_to_tile_26_2_2),
		.in_wire_2_3(horizontal_tile_26_1_to_tile_26_2_3),
		.out_wire_0_0(horizontal_tile_26_2_to_tile_26_3_0),
		.out_wire_0_1(horizontal_tile_26_2_to_tile_26_3_1),
		.out_wire_0_2(horizontal_tile_26_2_to_tile_26_3_2),
		.out_wire_0_3(horizontal_tile_26_2_to_tile_26_3_3),
		.in_wire_0_0(horizontal_tile_26_3_to_tile_26_2_0),
		.in_wire_0_1(horizontal_tile_26_3_to_tile_26_2_1),
		.in_wire_0_2(horizontal_tile_26_3_to_tile_26_2_2),
		.in_wire_0_3(horizontal_tile_26_3_to_tile_26_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(835)
	);

	pe_tile pe_tile_26_3(
		.out_wire_3_0(vertical_tile_26_3_to_tile_25_3_0),
		.out_wire_3_1(vertical_tile_26_3_to_tile_25_3_1),
		.out_wire_3_2(vertical_tile_26_3_to_tile_25_3_2),
		.out_wire_3_3(vertical_tile_26_3_to_tile_25_3_3),
		.in_wire_3_0(vertical_tile_25_3_to_tile_26_3_0),
		.in_wire_3_1(vertical_tile_25_3_to_tile_26_3_1),
		.in_wire_3_2(vertical_tile_25_3_to_tile_26_3_2),
		.in_wire_3_3(vertical_tile_25_3_to_tile_26_3_3),
		.out_wire_1_0(vertical_tile_26_3_to_tile_27_3_0),
		.out_wire_1_1(vertical_tile_26_3_to_tile_27_3_1),
		.out_wire_1_2(vertical_tile_26_3_to_tile_27_3_2),
		.out_wire_1_3(vertical_tile_26_3_to_tile_27_3_3),
		.in_wire_1_0(vertical_tile_27_3_to_tile_26_3_0),
		.in_wire_1_1(vertical_tile_27_3_to_tile_26_3_1),
		.in_wire_1_2(vertical_tile_27_3_to_tile_26_3_2),
		.in_wire_1_3(vertical_tile_27_3_to_tile_26_3_3),
		.out_wire_2_0(horizontal_tile_26_3_to_tile_26_2_0),
		.out_wire_2_1(horizontal_tile_26_3_to_tile_26_2_1),
		.out_wire_2_2(horizontal_tile_26_3_to_tile_26_2_2),
		.out_wire_2_3(horizontal_tile_26_3_to_tile_26_2_3),
		.in_wire_2_0(horizontal_tile_26_2_to_tile_26_3_0),
		.in_wire_2_1(horizontal_tile_26_2_to_tile_26_3_1),
		.in_wire_2_2(horizontal_tile_26_2_to_tile_26_3_2),
		.in_wire_2_3(horizontal_tile_26_2_to_tile_26_3_3),
		.out_wire_0_0(horizontal_tile_26_3_to_tile_26_4_0),
		.out_wire_0_1(horizontal_tile_26_3_to_tile_26_4_1),
		.out_wire_0_2(horizontal_tile_26_3_to_tile_26_4_2),
		.out_wire_0_3(horizontal_tile_26_3_to_tile_26_4_3),
		.in_wire_0_0(horizontal_tile_26_4_to_tile_26_3_0),
		.in_wire_0_1(horizontal_tile_26_4_to_tile_26_3_1),
		.in_wire_0_2(horizontal_tile_26_4_to_tile_26_3_2),
		.in_wire_0_3(horizontal_tile_26_4_to_tile_26_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(836)
	);

	pe_tile pe_tile_26_4(
		.out_wire_3_0(vertical_tile_26_4_to_tile_25_4_0),
		.out_wire_3_1(vertical_tile_26_4_to_tile_25_4_1),
		.out_wire_3_2(vertical_tile_26_4_to_tile_25_4_2),
		.out_wire_3_3(vertical_tile_26_4_to_tile_25_4_3),
		.in_wire_3_0(vertical_tile_25_4_to_tile_26_4_0),
		.in_wire_3_1(vertical_tile_25_4_to_tile_26_4_1),
		.in_wire_3_2(vertical_tile_25_4_to_tile_26_4_2),
		.in_wire_3_3(vertical_tile_25_4_to_tile_26_4_3),
		.out_wire_1_0(vertical_tile_26_4_to_tile_27_4_0),
		.out_wire_1_1(vertical_tile_26_4_to_tile_27_4_1),
		.out_wire_1_2(vertical_tile_26_4_to_tile_27_4_2),
		.out_wire_1_3(vertical_tile_26_4_to_tile_27_4_3),
		.in_wire_1_0(vertical_tile_27_4_to_tile_26_4_0),
		.in_wire_1_1(vertical_tile_27_4_to_tile_26_4_1),
		.in_wire_1_2(vertical_tile_27_4_to_tile_26_4_2),
		.in_wire_1_3(vertical_tile_27_4_to_tile_26_4_3),
		.out_wire_2_0(horizontal_tile_26_4_to_tile_26_3_0),
		.out_wire_2_1(horizontal_tile_26_4_to_tile_26_3_1),
		.out_wire_2_2(horizontal_tile_26_4_to_tile_26_3_2),
		.out_wire_2_3(horizontal_tile_26_4_to_tile_26_3_3),
		.in_wire_2_0(horizontal_tile_26_3_to_tile_26_4_0),
		.in_wire_2_1(horizontal_tile_26_3_to_tile_26_4_1),
		.in_wire_2_2(horizontal_tile_26_3_to_tile_26_4_2),
		.in_wire_2_3(horizontal_tile_26_3_to_tile_26_4_3),
		.out_wire_0_0(horizontal_tile_26_4_to_tile_26_5_0),
		.out_wire_0_1(horizontal_tile_26_4_to_tile_26_5_1),
		.out_wire_0_2(horizontal_tile_26_4_to_tile_26_5_2),
		.out_wire_0_3(horizontal_tile_26_4_to_tile_26_5_3),
		.in_wire_0_0(horizontal_tile_26_5_to_tile_26_4_0),
		.in_wire_0_1(horizontal_tile_26_5_to_tile_26_4_1),
		.in_wire_0_2(horizontal_tile_26_5_to_tile_26_4_2),
		.in_wire_0_3(horizontal_tile_26_5_to_tile_26_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(837)
	);

	pe_tile pe_tile_26_5(
		.out_wire_3_0(vertical_tile_26_5_to_tile_25_5_0),
		.out_wire_3_1(vertical_tile_26_5_to_tile_25_5_1),
		.out_wire_3_2(vertical_tile_26_5_to_tile_25_5_2),
		.out_wire_3_3(vertical_tile_26_5_to_tile_25_5_3),
		.in_wire_3_0(vertical_tile_25_5_to_tile_26_5_0),
		.in_wire_3_1(vertical_tile_25_5_to_tile_26_5_1),
		.in_wire_3_2(vertical_tile_25_5_to_tile_26_5_2),
		.in_wire_3_3(vertical_tile_25_5_to_tile_26_5_3),
		.out_wire_1_0(vertical_tile_26_5_to_tile_27_5_0),
		.out_wire_1_1(vertical_tile_26_5_to_tile_27_5_1),
		.out_wire_1_2(vertical_tile_26_5_to_tile_27_5_2),
		.out_wire_1_3(vertical_tile_26_5_to_tile_27_5_3),
		.in_wire_1_0(vertical_tile_27_5_to_tile_26_5_0),
		.in_wire_1_1(vertical_tile_27_5_to_tile_26_5_1),
		.in_wire_1_2(vertical_tile_27_5_to_tile_26_5_2),
		.in_wire_1_3(vertical_tile_27_5_to_tile_26_5_3),
		.out_wire_2_0(horizontal_tile_26_5_to_tile_26_4_0),
		.out_wire_2_1(horizontal_tile_26_5_to_tile_26_4_1),
		.out_wire_2_2(horizontal_tile_26_5_to_tile_26_4_2),
		.out_wire_2_3(horizontal_tile_26_5_to_tile_26_4_3),
		.in_wire_2_0(horizontal_tile_26_4_to_tile_26_5_0),
		.in_wire_2_1(horizontal_tile_26_4_to_tile_26_5_1),
		.in_wire_2_2(horizontal_tile_26_4_to_tile_26_5_2),
		.in_wire_2_3(horizontal_tile_26_4_to_tile_26_5_3),
		.out_wire_0_0(horizontal_tile_26_5_to_tile_26_6_0),
		.out_wire_0_1(horizontal_tile_26_5_to_tile_26_6_1),
		.out_wire_0_2(horizontal_tile_26_5_to_tile_26_6_2),
		.out_wire_0_3(horizontal_tile_26_5_to_tile_26_6_3),
		.in_wire_0_0(horizontal_tile_26_6_to_tile_26_5_0),
		.in_wire_0_1(horizontal_tile_26_6_to_tile_26_5_1),
		.in_wire_0_2(horizontal_tile_26_6_to_tile_26_5_2),
		.in_wire_0_3(horizontal_tile_26_6_to_tile_26_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(838)
	);

	pe_tile pe_tile_26_6(
		.out_wire_3_0(vertical_tile_26_6_to_tile_25_6_0),
		.out_wire_3_1(vertical_tile_26_6_to_tile_25_6_1),
		.out_wire_3_2(vertical_tile_26_6_to_tile_25_6_2),
		.out_wire_3_3(vertical_tile_26_6_to_tile_25_6_3),
		.in_wire_3_0(vertical_tile_25_6_to_tile_26_6_0),
		.in_wire_3_1(vertical_tile_25_6_to_tile_26_6_1),
		.in_wire_3_2(vertical_tile_25_6_to_tile_26_6_2),
		.in_wire_3_3(vertical_tile_25_6_to_tile_26_6_3),
		.out_wire_1_0(vertical_tile_26_6_to_tile_27_6_0),
		.out_wire_1_1(vertical_tile_26_6_to_tile_27_6_1),
		.out_wire_1_2(vertical_tile_26_6_to_tile_27_6_2),
		.out_wire_1_3(vertical_tile_26_6_to_tile_27_6_3),
		.in_wire_1_0(vertical_tile_27_6_to_tile_26_6_0),
		.in_wire_1_1(vertical_tile_27_6_to_tile_26_6_1),
		.in_wire_1_2(vertical_tile_27_6_to_tile_26_6_2),
		.in_wire_1_3(vertical_tile_27_6_to_tile_26_6_3),
		.out_wire_2_0(horizontal_tile_26_6_to_tile_26_5_0),
		.out_wire_2_1(horizontal_tile_26_6_to_tile_26_5_1),
		.out_wire_2_2(horizontal_tile_26_6_to_tile_26_5_2),
		.out_wire_2_3(horizontal_tile_26_6_to_tile_26_5_3),
		.in_wire_2_0(horizontal_tile_26_5_to_tile_26_6_0),
		.in_wire_2_1(horizontal_tile_26_5_to_tile_26_6_1),
		.in_wire_2_2(horizontal_tile_26_5_to_tile_26_6_2),
		.in_wire_2_3(horizontal_tile_26_5_to_tile_26_6_3),
		.out_wire_0_0(horizontal_tile_26_6_to_tile_26_7_0),
		.out_wire_0_1(horizontal_tile_26_6_to_tile_26_7_1),
		.out_wire_0_2(horizontal_tile_26_6_to_tile_26_7_2),
		.out_wire_0_3(horizontal_tile_26_6_to_tile_26_7_3),
		.in_wire_0_0(horizontal_tile_26_7_to_tile_26_6_0),
		.in_wire_0_1(horizontal_tile_26_7_to_tile_26_6_1),
		.in_wire_0_2(horizontal_tile_26_7_to_tile_26_6_2),
		.in_wire_0_3(horizontal_tile_26_7_to_tile_26_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(839)
	);

	pe_tile pe_tile_26_7(
		.out_wire_3_0(vertical_tile_26_7_to_tile_25_7_0),
		.out_wire_3_1(vertical_tile_26_7_to_tile_25_7_1),
		.out_wire_3_2(vertical_tile_26_7_to_tile_25_7_2),
		.out_wire_3_3(vertical_tile_26_7_to_tile_25_7_3),
		.in_wire_3_0(vertical_tile_25_7_to_tile_26_7_0),
		.in_wire_3_1(vertical_tile_25_7_to_tile_26_7_1),
		.in_wire_3_2(vertical_tile_25_7_to_tile_26_7_2),
		.in_wire_3_3(vertical_tile_25_7_to_tile_26_7_3),
		.out_wire_1_0(vertical_tile_26_7_to_tile_27_7_0),
		.out_wire_1_1(vertical_tile_26_7_to_tile_27_7_1),
		.out_wire_1_2(vertical_tile_26_7_to_tile_27_7_2),
		.out_wire_1_3(vertical_tile_26_7_to_tile_27_7_3),
		.in_wire_1_0(vertical_tile_27_7_to_tile_26_7_0),
		.in_wire_1_1(vertical_tile_27_7_to_tile_26_7_1),
		.in_wire_1_2(vertical_tile_27_7_to_tile_26_7_2),
		.in_wire_1_3(vertical_tile_27_7_to_tile_26_7_3),
		.out_wire_2_0(horizontal_tile_26_7_to_tile_26_6_0),
		.out_wire_2_1(horizontal_tile_26_7_to_tile_26_6_1),
		.out_wire_2_2(horizontal_tile_26_7_to_tile_26_6_2),
		.out_wire_2_3(horizontal_tile_26_7_to_tile_26_6_3),
		.in_wire_2_0(horizontal_tile_26_6_to_tile_26_7_0),
		.in_wire_2_1(horizontal_tile_26_6_to_tile_26_7_1),
		.in_wire_2_2(horizontal_tile_26_6_to_tile_26_7_2),
		.in_wire_2_3(horizontal_tile_26_6_to_tile_26_7_3),
		.out_wire_0_0(horizontal_tile_26_7_to_tile_26_8_0),
		.out_wire_0_1(horizontal_tile_26_7_to_tile_26_8_1),
		.out_wire_0_2(horizontal_tile_26_7_to_tile_26_8_2),
		.out_wire_0_3(horizontal_tile_26_7_to_tile_26_8_3),
		.in_wire_0_0(horizontal_tile_26_8_to_tile_26_7_0),
		.in_wire_0_1(horizontal_tile_26_8_to_tile_26_7_1),
		.in_wire_0_2(horizontal_tile_26_8_to_tile_26_7_2),
		.in_wire_0_3(horizontal_tile_26_8_to_tile_26_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(840)
	);

	pe_tile pe_tile_26_8(
		.out_wire_3_0(vertical_tile_26_8_to_tile_25_8_0),
		.out_wire_3_1(vertical_tile_26_8_to_tile_25_8_1),
		.out_wire_3_2(vertical_tile_26_8_to_tile_25_8_2),
		.out_wire_3_3(vertical_tile_26_8_to_tile_25_8_3),
		.in_wire_3_0(vertical_tile_25_8_to_tile_26_8_0),
		.in_wire_3_1(vertical_tile_25_8_to_tile_26_8_1),
		.in_wire_3_2(vertical_tile_25_8_to_tile_26_8_2),
		.in_wire_3_3(vertical_tile_25_8_to_tile_26_8_3),
		.out_wire_1_0(vertical_tile_26_8_to_tile_27_8_0),
		.out_wire_1_1(vertical_tile_26_8_to_tile_27_8_1),
		.out_wire_1_2(vertical_tile_26_8_to_tile_27_8_2),
		.out_wire_1_3(vertical_tile_26_8_to_tile_27_8_3),
		.in_wire_1_0(vertical_tile_27_8_to_tile_26_8_0),
		.in_wire_1_1(vertical_tile_27_8_to_tile_26_8_1),
		.in_wire_1_2(vertical_tile_27_8_to_tile_26_8_2),
		.in_wire_1_3(vertical_tile_27_8_to_tile_26_8_3),
		.out_wire_2_0(horizontal_tile_26_8_to_tile_26_7_0),
		.out_wire_2_1(horizontal_tile_26_8_to_tile_26_7_1),
		.out_wire_2_2(horizontal_tile_26_8_to_tile_26_7_2),
		.out_wire_2_3(horizontal_tile_26_8_to_tile_26_7_3),
		.in_wire_2_0(horizontal_tile_26_7_to_tile_26_8_0),
		.in_wire_2_1(horizontal_tile_26_7_to_tile_26_8_1),
		.in_wire_2_2(horizontal_tile_26_7_to_tile_26_8_2),
		.in_wire_2_3(horizontal_tile_26_7_to_tile_26_8_3),
		.out_wire_0_0(horizontal_tile_26_8_to_tile_26_9_0),
		.out_wire_0_1(horizontal_tile_26_8_to_tile_26_9_1),
		.out_wire_0_2(horizontal_tile_26_8_to_tile_26_9_2),
		.out_wire_0_3(horizontal_tile_26_8_to_tile_26_9_3),
		.in_wire_0_0(horizontal_tile_26_9_to_tile_26_8_0),
		.in_wire_0_1(horizontal_tile_26_9_to_tile_26_8_1),
		.in_wire_0_2(horizontal_tile_26_9_to_tile_26_8_2),
		.in_wire_0_3(horizontal_tile_26_9_to_tile_26_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(841)
	);

	pe_tile pe_tile_26_9(
		.out_wire_3_0(vertical_tile_26_9_to_tile_25_9_0),
		.out_wire_3_1(vertical_tile_26_9_to_tile_25_9_1),
		.out_wire_3_2(vertical_tile_26_9_to_tile_25_9_2),
		.out_wire_3_3(vertical_tile_26_9_to_tile_25_9_3),
		.in_wire_3_0(vertical_tile_25_9_to_tile_26_9_0),
		.in_wire_3_1(vertical_tile_25_9_to_tile_26_9_1),
		.in_wire_3_2(vertical_tile_25_9_to_tile_26_9_2),
		.in_wire_3_3(vertical_tile_25_9_to_tile_26_9_3),
		.out_wire_1_0(vertical_tile_26_9_to_tile_27_9_0),
		.out_wire_1_1(vertical_tile_26_9_to_tile_27_9_1),
		.out_wire_1_2(vertical_tile_26_9_to_tile_27_9_2),
		.out_wire_1_3(vertical_tile_26_9_to_tile_27_9_3),
		.in_wire_1_0(vertical_tile_27_9_to_tile_26_9_0),
		.in_wire_1_1(vertical_tile_27_9_to_tile_26_9_1),
		.in_wire_1_2(vertical_tile_27_9_to_tile_26_9_2),
		.in_wire_1_3(vertical_tile_27_9_to_tile_26_9_3),
		.out_wire_2_0(horizontal_tile_26_9_to_tile_26_8_0),
		.out_wire_2_1(horizontal_tile_26_9_to_tile_26_8_1),
		.out_wire_2_2(horizontal_tile_26_9_to_tile_26_8_2),
		.out_wire_2_3(horizontal_tile_26_9_to_tile_26_8_3),
		.in_wire_2_0(horizontal_tile_26_8_to_tile_26_9_0),
		.in_wire_2_1(horizontal_tile_26_8_to_tile_26_9_1),
		.in_wire_2_2(horizontal_tile_26_8_to_tile_26_9_2),
		.in_wire_2_3(horizontal_tile_26_8_to_tile_26_9_3),
		.out_wire_0_0(horizontal_tile_26_9_to_tile_26_10_0),
		.out_wire_0_1(horizontal_tile_26_9_to_tile_26_10_1),
		.out_wire_0_2(horizontal_tile_26_9_to_tile_26_10_2),
		.out_wire_0_3(horizontal_tile_26_9_to_tile_26_10_3),
		.in_wire_0_0(horizontal_tile_26_10_to_tile_26_9_0),
		.in_wire_0_1(horizontal_tile_26_10_to_tile_26_9_1),
		.in_wire_0_2(horizontal_tile_26_10_to_tile_26_9_2),
		.in_wire_0_3(horizontal_tile_26_10_to_tile_26_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(842)
	);

	pe_tile pe_tile_26_10(
		.out_wire_3_0(vertical_tile_26_10_to_tile_25_10_0),
		.out_wire_3_1(vertical_tile_26_10_to_tile_25_10_1),
		.out_wire_3_2(vertical_tile_26_10_to_tile_25_10_2),
		.out_wire_3_3(vertical_tile_26_10_to_tile_25_10_3),
		.in_wire_3_0(vertical_tile_25_10_to_tile_26_10_0),
		.in_wire_3_1(vertical_tile_25_10_to_tile_26_10_1),
		.in_wire_3_2(vertical_tile_25_10_to_tile_26_10_2),
		.in_wire_3_3(vertical_tile_25_10_to_tile_26_10_3),
		.out_wire_1_0(vertical_tile_26_10_to_tile_27_10_0),
		.out_wire_1_1(vertical_tile_26_10_to_tile_27_10_1),
		.out_wire_1_2(vertical_tile_26_10_to_tile_27_10_2),
		.out_wire_1_3(vertical_tile_26_10_to_tile_27_10_3),
		.in_wire_1_0(vertical_tile_27_10_to_tile_26_10_0),
		.in_wire_1_1(vertical_tile_27_10_to_tile_26_10_1),
		.in_wire_1_2(vertical_tile_27_10_to_tile_26_10_2),
		.in_wire_1_3(vertical_tile_27_10_to_tile_26_10_3),
		.out_wire_2_0(horizontal_tile_26_10_to_tile_26_9_0),
		.out_wire_2_1(horizontal_tile_26_10_to_tile_26_9_1),
		.out_wire_2_2(horizontal_tile_26_10_to_tile_26_9_2),
		.out_wire_2_3(horizontal_tile_26_10_to_tile_26_9_3),
		.in_wire_2_0(horizontal_tile_26_9_to_tile_26_10_0),
		.in_wire_2_1(horizontal_tile_26_9_to_tile_26_10_1),
		.in_wire_2_2(horizontal_tile_26_9_to_tile_26_10_2),
		.in_wire_2_3(horizontal_tile_26_9_to_tile_26_10_3),
		.out_wire_0_0(horizontal_tile_26_10_to_tile_26_11_0),
		.out_wire_0_1(horizontal_tile_26_10_to_tile_26_11_1),
		.out_wire_0_2(horizontal_tile_26_10_to_tile_26_11_2),
		.out_wire_0_3(horizontal_tile_26_10_to_tile_26_11_3),
		.in_wire_0_0(horizontal_tile_26_11_to_tile_26_10_0),
		.in_wire_0_1(horizontal_tile_26_11_to_tile_26_10_1),
		.in_wire_0_2(horizontal_tile_26_11_to_tile_26_10_2),
		.in_wire_0_3(horizontal_tile_26_11_to_tile_26_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(843)
	);

	pe_tile pe_tile_26_11(
		.out_wire_3_0(vertical_tile_26_11_to_tile_25_11_0),
		.out_wire_3_1(vertical_tile_26_11_to_tile_25_11_1),
		.out_wire_3_2(vertical_tile_26_11_to_tile_25_11_2),
		.out_wire_3_3(vertical_tile_26_11_to_tile_25_11_3),
		.in_wire_3_0(vertical_tile_25_11_to_tile_26_11_0),
		.in_wire_3_1(vertical_tile_25_11_to_tile_26_11_1),
		.in_wire_3_2(vertical_tile_25_11_to_tile_26_11_2),
		.in_wire_3_3(vertical_tile_25_11_to_tile_26_11_3),
		.out_wire_1_0(vertical_tile_26_11_to_tile_27_11_0),
		.out_wire_1_1(vertical_tile_26_11_to_tile_27_11_1),
		.out_wire_1_2(vertical_tile_26_11_to_tile_27_11_2),
		.out_wire_1_3(vertical_tile_26_11_to_tile_27_11_3),
		.in_wire_1_0(vertical_tile_27_11_to_tile_26_11_0),
		.in_wire_1_1(vertical_tile_27_11_to_tile_26_11_1),
		.in_wire_1_2(vertical_tile_27_11_to_tile_26_11_2),
		.in_wire_1_3(vertical_tile_27_11_to_tile_26_11_3),
		.out_wire_2_0(horizontal_tile_26_11_to_tile_26_10_0),
		.out_wire_2_1(horizontal_tile_26_11_to_tile_26_10_1),
		.out_wire_2_2(horizontal_tile_26_11_to_tile_26_10_2),
		.out_wire_2_3(horizontal_tile_26_11_to_tile_26_10_3),
		.in_wire_2_0(horizontal_tile_26_10_to_tile_26_11_0),
		.in_wire_2_1(horizontal_tile_26_10_to_tile_26_11_1),
		.in_wire_2_2(horizontal_tile_26_10_to_tile_26_11_2),
		.in_wire_2_3(horizontal_tile_26_10_to_tile_26_11_3),
		.out_wire_0_0(horizontal_tile_26_11_to_tile_26_12_0),
		.out_wire_0_1(horizontal_tile_26_11_to_tile_26_12_1),
		.out_wire_0_2(horizontal_tile_26_11_to_tile_26_12_2),
		.out_wire_0_3(horizontal_tile_26_11_to_tile_26_12_3),
		.in_wire_0_0(horizontal_tile_26_12_to_tile_26_11_0),
		.in_wire_0_1(horizontal_tile_26_12_to_tile_26_11_1),
		.in_wire_0_2(horizontal_tile_26_12_to_tile_26_11_2),
		.in_wire_0_3(horizontal_tile_26_12_to_tile_26_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(844)
	);

	pe_tile pe_tile_26_12(
		.out_wire_3_0(vertical_tile_26_12_to_tile_25_12_0),
		.out_wire_3_1(vertical_tile_26_12_to_tile_25_12_1),
		.out_wire_3_2(vertical_tile_26_12_to_tile_25_12_2),
		.out_wire_3_3(vertical_tile_26_12_to_tile_25_12_3),
		.in_wire_3_0(vertical_tile_25_12_to_tile_26_12_0),
		.in_wire_3_1(vertical_tile_25_12_to_tile_26_12_1),
		.in_wire_3_2(vertical_tile_25_12_to_tile_26_12_2),
		.in_wire_3_3(vertical_tile_25_12_to_tile_26_12_3),
		.out_wire_1_0(vertical_tile_26_12_to_tile_27_12_0),
		.out_wire_1_1(vertical_tile_26_12_to_tile_27_12_1),
		.out_wire_1_2(vertical_tile_26_12_to_tile_27_12_2),
		.out_wire_1_3(vertical_tile_26_12_to_tile_27_12_3),
		.in_wire_1_0(vertical_tile_27_12_to_tile_26_12_0),
		.in_wire_1_1(vertical_tile_27_12_to_tile_26_12_1),
		.in_wire_1_2(vertical_tile_27_12_to_tile_26_12_2),
		.in_wire_1_3(vertical_tile_27_12_to_tile_26_12_3),
		.out_wire_2_0(horizontal_tile_26_12_to_tile_26_11_0),
		.out_wire_2_1(horizontal_tile_26_12_to_tile_26_11_1),
		.out_wire_2_2(horizontal_tile_26_12_to_tile_26_11_2),
		.out_wire_2_3(horizontal_tile_26_12_to_tile_26_11_3),
		.in_wire_2_0(horizontal_tile_26_11_to_tile_26_12_0),
		.in_wire_2_1(horizontal_tile_26_11_to_tile_26_12_1),
		.in_wire_2_2(horizontal_tile_26_11_to_tile_26_12_2),
		.in_wire_2_3(horizontal_tile_26_11_to_tile_26_12_3),
		.out_wire_0_0(horizontal_tile_26_12_to_tile_26_13_0),
		.out_wire_0_1(horizontal_tile_26_12_to_tile_26_13_1),
		.out_wire_0_2(horizontal_tile_26_12_to_tile_26_13_2),
		.out_wire_0_3(horizontal_tile_26_12_to_tile_26_13_3),
		.in_wire_0_0(horizontal_tile_26_13_to_tile_26_12_0),
		.in_wire_0_1(horizontal_tile_26_13_to_tile_26_12_1),
		.in_wire_0_2(horizontal_tile_26_13_to_tile_26_12_2),
		.in_wire_0_3(horizontal_tile_26_13_to_tile_26_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(845)
	);

	pe_tile pe_tile_26_13(
		.out_wire_3_0(vertical_tile_26_13_to_tile_25_13_0),
		.out_wire_3_1(vertical_tile_26_13_to_tile_25_13_1),
		.out_wire_3_2(vertical_tile_26_13_to_tile_25_13_2),
		.out_wire_3_3(vertical_tile_26_13_to_tile_25_13_3),
		.in_wire_3_0(vertical_tile_25_13_to_tile_26_13_0),
		.in_wire_3_1(vertical_tile_25_13_to_tile_26_13_1),
		.in_wire_3_2(vertical_tile_25_13_to_tile_26_13_2),
		.in_wire_3_3(vertical_tile_25_13_to_tile_26_13_3),
		.out_wire_1_0(vertical_tile_26_13_to_tile_27_13_0),
		.out_wire_1_1(vertical_tile_26_13_to_tile_27_13_1),
		.out_wire_1_2(vertical_tile_26_13_to_tile_27_13_2),
		.out_wire_1_3(vertical_tile_26_13_to_tile_27_13_3),
		.in_wire_1_0(vertical_tile_27_13_to_tile_26_13_0),
		.in_wire_1_1(vertical_tile_27_13_to_tile_26_13_1),
		.in_wire_1_2(vertical_tile_27_13_to_tile_26_13_2),
		.in_wire_1_3(vertical_tile_27_13_to_tile_26_13_3),
		.out_wire_2_0(horizontal_tile_26_13_to_tile_26_12_0),
		.out_wire_2_1(horizontal_tile_26_13_to_tile_26_12_1),
		.out_wire_2_2(horizontal_tile_26_13_to_tile_26_12_2),
		.out_wire_2_3(horizontal_tile_26_13_to_tile_26_12_3),
		.in_wire_2_0(horizontal_tile_26_12_to_tile_26_13_0),
		.in_wire_2_1(horizontal_tile_26_12_to_tile_26_13_1),
		.in_wire_2_2(horizontal_tile_26_12_to_tile_26_13_2),
		.in_wire_2_3(horizontal_tile_26_12_to_tile_26_13_3),
		.out_wire_0_0(horizontal_tile_26_13_to_tile_26_14_0),
		.out_wire_0_1(horizontal_tile_26_13_to_tile_26_14_1),
		.out_wire_0_2(horizontal_tile_26_13_to_tile_26_14_2),
		.out_wire_0_3(horizontal_tile_26_13_to_tile_26_14_3),
		.in_wire_0_0(horizontal_tile_26_14_to_tile_26_13_0),
		.in_wire_0_1(horizontal_tile_26_14_to_tile_26_13_1),
		.in_wire_0_2(horizontal_tile_26_14_to_tile_26_13_2),
		.in_wire_0_3(horizontal_tile_26_14_to_tile_26_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(846)
	);

	pe_tile pe_tile_26_14(
		.out_wire_3_0(vertical_tile_26_14_to_tile_25_14_0),
		.out_wire_3_1(vertical_tile_26_14_to_tile_25_14_1),
		.out_wire_3_2(vertical_tile_26_14_to_tile_25_14_2),
		.out_wire_3_3(vertical_tile_26_14_to_tile_25_14_3),
		.in_wire_3_0(vertical_tile_25_14_to_tile_26_14_0),
		.in_wire_3_1(vertical_tile_25_14_to_tile_26_14_1),
		.in_wire_3_2(vertical_tile_25_14_to_tile_26_14_2),
		.in_wire_3_3(vertical_tile_25_14_to_tile_26_14_3),
		.out_wire_1_0(vertical_tile_26_14_to_tile_27_14_0),
		.out_wire_1_1(vertical_tile_26_14_to_tile_27_14_1),
		.out_wire_1_2(vertical_tile_26_14_to_tile_27_14_2),
		.out_wire_1_3(vertical_tile_26_14_to_tile_27_14_3),
		.in_wire_1_0(vertical_tile_27_14_to_tile_26_14_0),
		.in_wire_1_1(vertical_tile_27_14_to_tile_26_14_1),
		.in_wire_1_2(vertical_tile_27_14_to_tile_26_14_2),
		.in_wire_1_3(vertical_tile_27_14_to_tile_26_14_3),
		.out_wire_2_0(horizontal_tile_26_14_to_tile_26_13_0),
		.out_wire_2_1(horizontal_tile_26_14_to_tile_26_13_1),
		.out_wire_2_2(horizontal_tile_26_14_to_tile_26_13_2),
		.out_wire_2_3(horizontal_tile_26_14_to_tile_26_13_3),
		.in_wire_2_0(horizontal_tile_26_13_to_tile_26_14_0),
		.in_wire_2_1(horizontal_tile_26_13_to_tile_26_14_1),
		.in_wire_2_2(horizontal_tile_26_13_to_tile_26_14_2),
		.in_wire_2_3(horizontal_tile_26_13_to_tile_26_14_3),
		.out_wire_0_0(horizontal_tile_26_14_to_tile_26_15_0),
		.out_wire_0_1(horizontal_tile_26_14_to_tile_26_15_1),
		.out_wire_0_2(horizontal_tile_26_14_to_tile_26_15_2),
		.out_wire_0_3(horizontal_tile_26_14_to_tile_26_15_3),
		.in_wire_0_0(horizontal_tile_26_15_to_tile_26_14_0),
		.in_wire_0_1(horizontal_tile_26_15_to_tile_26_14_1),
		.in_wire_0_2(horizontal_tile_26_15_to_tile_26_14_2),
		.in_wire_0_3(horizontal_tile_26_15_to_tile_26_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(847)
	);

	pe_tile pe_tile_26_15(
		.out_wire_3_0(vertical_tile_26_15_to_tile_25_15_0),
		.out_wire_3_1(vertical_tile_26_15_to_tile_25_15_1),
		.out_wire_3_2(vertical_tile_26_15_to_tile_25_15_2),
		.out_wire_3_3(vertical_tile_26_15_to_tile_25_15_3),
		.in_wire_3_0(vertical_tile_25_15_to_tile_26_15_0),
		.in_wire_3_1(vertical_tile_25_15_to_tile_26_15_1),
		.in_wire_3_2(vertical_tile_25_15_to_tile_26_15_2),
		.in_wire_3_3(vertical_tile_25_15_to_tile_26_15_3),
		.out_wire_1_0(vertical_tile_26_15_to_tile_27_15_0),
		.out_wire_1_1(vertical_tile_26_15_to_tile_27_15_1),
		.out_wire_1_2(vertical_tile_26_15_to_tile_27_15_2),
		.out_wire_1_3(vertical_tile_26_15_to_tile_27_15_3),
		.in_wire_1_0(vertical_tile_27_15_to_tile_26_15_0),
		.in_wire_1_1(vertical_tile_27_15_to_tile_26_15_1),
		.in_wire_1_2(vertical_tile_27_15_to_tile_26_15_2),
		.in_wire_1_3(vertical_tile_27_15_to_tile_26_15_3),
		.out_wire_2_0(horizontal_tile_26_15_to_tile_26_14_0),
		.out_wire_2_1(horizontal_tile_26_15_to_tile_26_14_1),
		.out_wire_2_2(horizontal_tile_26_15_to_tile_26_14_2),
		.out_wire_2_3(horizontal_tile_26_15_to_tile_26_14_3),
		.in_wire_2_0(horizontal_tile_26_14_to_tile_26_15_0),
		.in_wire_2_1(horizontal_tile_26_14_to_tile_26_15_1),
		.in_wire_2_2(horizontal_tile_26_14_to_tile_26_15_2),
		.in_wire_2_3(horizontal_tile_26_14_to_tile_26_15_3),
		.out_wire_0_0(horizontal_tile_26_15_to_tile_26_16_0),
		.out_wire_0_1(horizontal_tile_26_15_to_tile_26_16_1),
		.out_wire_0_2(horizontal_tile_26_15_to_tile_26_16_2),
		.out_wire_0_3(horizontal_tile_26_15_to_tile_26_16_3),
		.in_wire_0_0(horizontal_tile_26_16_to_tile_26_15_0),
		.in_wire_0_1(horizontal_tile_26_16_to_tile_26_15_1),
		.in_wire_0_2(horizontal_tile_26_16_to_tile_26_15_2),
		.in_wire_0_3(horizontal_tile_26_16_to_tile_26_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(848)
	);

	pe_tile pe_tile_26_16(
		.out_wire_3_0(vertical_tile_26_16_to_tile_25_16_0),
		.out_wire_3_1(vertical_tile_26_16_to_tile_25_16_1),
		.out_wire_3_2(vertical_tile_26_16_to_tile_25_16_2),
		.out_wire_3_3(vertical_tile_26_16_to_tile_25_16_3),
		.in_wire_3_0(vertical_tile_25_16_to_tile_26_16_0),
		.in_wire_3_1(vertical_tile_25_16_to_tile_26_16_1),
		.in_wire_3_2(vertical_tile_25_16_to_tile_26_16_2),
		.in_wire_3_3(vertical_tile_25_16_to_tile_26_16_3),
		.out_wire_1_0(vertical_tile_26_16_to_tile_27_16_0),
		.out_wire_1_1(vertical_tile_26_16_to_tile_27_16_1),
		.out_wire_1_2(vertical_tile_26_16_to_tile_27_16_2),
		.out_wire_1_3(vertical_tile_26_16_to_tile_27_16_3),
		.in_wire_1_0(vertical_tile_27_16_to_tile_26_16_0),
		.in_wire_1_1(vertical_tile_27_16_to_tile_26_16_1),
		.in_wire_1_2(vertical_tile_27_16_to_tile_26_16_2),
		.in_wire_1_3(vertical_tile_27_16_to_tile_26_16_3),
		.out_wire_2_0(horizontal_tile_26_16_to_tile_26_15_0),
		.out_wire_2_1(horizontal_tile_26_16_to_tile_26_15_1),
		.out_wire_2_2(horizontal_tile_26_16_to_tile_26_15_2),
		.out_wire_2_3(horizontal_tile_26_16_to_tile_26_15_3),
		.in_wire_2_0(horizontal_tile_26_15_to_tile_26_16_0),
		.in_wire_2_1(horizontal_tile_26_15_to_tile_26_16_1),
		.in_wire_2_2(horizontal_tile_26_15_to_tile_26_16_2),
		.in_wire_2_3(horizontal_tile_26_15_to_tile_26_16_3),
		.out_wire_0_0(horizontal_tile_26_16_to_tile_26_17_0),
		.out_wire_0_1(horizontal_tile_26_16_to_tile_26_17_1),
		.out_wire_0_2(horizontal_tile_26_16_to_tile_26_17_2),
		.out_wire_0_3(horizontal_tile_26_16_to_tile_26_17_3),
		.in_wire_0_0(horizontal_tile_26_17_to_tile_26_16_0),
		.in_wire_0_1(horizontal_tile_26_17_to_tile_26_16_1),
		.in_wire_0_2(horizontal_tile_26_17_to_tile_26_16_2),
		.in_wire_0_3(horizontal_tile_26_17_to_tile_26_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(849)
	);

	pe_tile pe_tile_26_17(
		.out_wire_3_0(vertical_tile_26_17_to_tile_25_17_0),
		.out_wire_3_1(vertical_tile_26_17_to_tile_25_17_1),
		.out_wire_3_2(vertical_tile_26_17_to_tile_25_17_2),
		.out_wire_3_3(vertical_tile_26_17_to_tile_25_17_3),
		.in_wire_3_0(vertical_tile_25_17_to_tile_26_17_0),
		.in_wire_3_1(vertical_tile_25_17_to_tile_26_17_1),
		.in_wire_3_2(vertical_tile_25_17_to_tile_26_17_2),
		.in_wire_3_3(vertical_tile_25_17_to_tile_26_17_3),
		.out_wire_1_0(vertical_tile_26_17_to_tile_27_17_0),
		.out_wire_1_1(vertical_tile_26_17_to_tile_27_17_1),
		.out_wire_1_2(vertical_tile_26_17_to_tile_27_17_2),
		.out_wire_1_3(vertical_tile_26_17_to_tile_27_17_3),
		.in_wire_1_0(vertical_tile_27_17_to_tile_26_17_0),
		.in_wire_1_1(vertical_tile_27_17_to_tile_26_17_1),
		.in_wire_1_2(vertical_tile_27_17_to_tile_26_17_2),
		.in_wire_1_3(vertical_tile_27_17_to_tile_26_17_3),
		.out_wire_2_0(horizontal_tile_26_17_to_tile_26_16_0),
		.out_wire_2_1(horizontal_tile_26_17_to_tile_26_16_1),
		.out_wire_2_2(horizontal_tile_26_17_to_tile_26_16_2),
		.out_wire_2_3(horizontal_tile_26_17_to_tile_26_16_3),
		.in_wire_2_0(horizontal_tile_26_16_to_tile_26_17_0),
		.in_wire_2_1(horizontal_tile_26_16_to_tile_26_17_1),
		.in_wire_2_2(horizontal_tile_26_16_to_tile_26_17_2),
		.in_wire_2_3(horizontal_tile_26_16_to_tile_26_17_3),
		.out_wire_0_0(horizontal_tile_26_17_to_tile_26_18_0),
		.out_wire_0_1(horizontal_tile_26_17_to_tile_26_18_1),
		.out_wire_0_2(horizontal_tile_26_17_to_tile_26_18_2),
		.out_wire_0_3(horizontal_tile_26_17_to_tile_26_18_3),
		.in_wire_0_0(horizontal_tile_26_18_to_tile_26_17_0),
		.in_wire_0_1(horizontal_tile_26_18_to_tile_26_17_1),
		.in_wire_0_2(horizontal_tile_26_18_to_tile_26_17_2),
		.in_wire_0_3(horizontal_tile_26_18_to_tile_26_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(850)
	);

	pe_tile pe_tile_26_18(
		.out_wire_3_0(vertical_tile_26_18_to_tile_25_18_0),
		.out_wire_3_1(vertical_tile_26_18_to_tile_25_18_1),
		.out_wire_3_2(vertical_tile_26_18_to_tile_25_18_2),
		.out_wire_3_3(vertical_tile_26_18_to_tile_25_18_3),
		.in_wire_3_0(vertical_tile_25_18_to_tile_26_18_0),
		.in_wire_3_1(vertical_tile_25_18_to_tile_26_18_1),
		.in_wire_3_2(vertical_tile_25_18_to_tile_26_18_2),
		.in_wire_3_3(vertical_tile_25_18_to_tile_26_18_3),
		.out_wire_1_0(vertical_tile_26_18_to_tile_27_18_0),
		.out_wire_1_1(vertical_tile_26_18_to_tile_27_18_1),
		.out_wire_1_2(vertical_tile_26_18_to_tile_27_18_2),
		.out_wire_1_3(vertical_tile_26_18_to_tile_27_18_3),
		.in_wire_1_0(vertical_tile_27_18_to_tile_26_18_0),
		.in_wire_1_1(vertical_tile_27_18_to_tile_26_18_1),
		.in_wire_1_2(vertical_tile_27_18_to_tile_26_18_2),
		.in_wire_1_3(vertical_tile_27_18_to_tile_26_18_3),
		.out_wire_2_0(horizontal_tile_26_18_to_tile_26_17_0),
		.out_wire_2_1(horizontal_tile_26_18_to_tile_26_17_1),
		.out_wire_2_2(horizontal_tile_26_18_to_tile_26_17_2),
		.out_wire_2_3(horizontal_tile_26_18_to_tile_26_17_3),
		.in_wire_2_0(horizontal_tile_26_17_to_tile_26_18_0),
		.in_wire_2_1(horizontal_tile_26_17_to_tile_26_18_1),
		.in_wire_2_2(horizontal_tile_26_17_to_tile_26_18_2),
		.in_wire_2_3(horizontal_tile_26_17_to_tile_26_18_3),
		.out_wire_0_0(horizontal_tile_26_18_to_tile_26_19_0),
		.out_wire_0_1(horizontal_tile_26_18_to_tile_26_19_1),
		.out_wire_0_2(horizontal_tile_26_18_to_tile_26_19_2),
		.out_wire_0_3(horizontal_tile_26_18_to_tile_26_19_3),
		.in_wire_0_0(horizontal_tile_26_19_to_tile_26_18_0),
		.in_wire_0_1(horizontal_tile_26_19_to_tile_26_18_1),
		.in_wire_0_2(horizontal_tile_26_19_to_tile_26_18_2),
		.in_wire_0_3(horizontal_tile_26_19_to_tile_26_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(851)
	);

	pe_tile pe_tile_26_19(
		.out_wire_3_0(vertical_tile_26_19_to_tile_25_19_0),
		.out_wire_3_1(vertical_tile_26_19_to_tile_25_19_1),
		.out_wire_3_2(vertical_tile_26_19_to_tile_25_19_2),
		.out_wire_3_3(vertical_tile_26_19_to_tile_25_19_3),
		.in_wire_3_0(vertical_tile_25_19_to_tile_26_19_0),
		.in_wire_3_1(vertical_tile_25_19_to_tile_26_19_1),
		.in_wire_3_2(vertical_tile_25_19_to_tile_26_19_2),
		.in_wire_3_3(vertical_tile_25_19_to_tile_26_19_3),
		.out_wire_1_0(vertical_tile_26_19_to_tile_27_19_0),
		.out_wire_1_1(vertical_tile_26_19_to_tile_27_19_1),
		.out_wire_1_2(vertical_tile_26_19_to_tile_27_19_2),
		.out_wire_1_3(vertical_tile_26_19_to_tile_27_19_3),
		.in_wire_1_0(vertical_tile_27_19_to_tile_26_19_0),
		.in_wire_1_1(vertical_tile_27_19_to_tile_26_19_1),
		.in_wire_1_2(vertical_tile_27_19_to_tile_26_19_2),
		.in_wire_1_3(vertical_tile_27_19_to_tile_26_19_3),
		.out_wire_2_0(horizontal_tile_26_19_to_tile_26_18_0),
		.out_wire_2_1(horizontal_tile_26_19_to_tile_26_18_1),
		.out_wire_2_2(horizontal_tile_26_19_to_tile_26_18_2),
		.out_wire_2_3(horizontal_tile_26_19_to_tile_26_18_3),
		.in_wire_2_0(horizontal_tile_26_18_to_tile_26_19_0),
		.in_wire_2_1(horizontal_tile_26_18_to_tile_26_19_1),
		.in_wire_2_2(horizontal_tile_26_18_to_tile_26_19_2),
		.in_wire_2_3(horizontal_tile_26_18_to_tile_26_19_3),
		.out_wire_0_0(horizontal_tile_26_19_to_tile_26_20_0),
		.out_wire_0_1(horizontal_tile_26_19_to_tile_26_20_1),
		.out_wire_0_2(horizontal_tile_26_19_to_tile_26_20_2),
		.out_wire_0_3(horizontal_tile_26_19_to_tile_26_20_3),
		.in_wire_0_0(horizontal_tile_26_20_to_tile_26_19_0),
		.in_wire_0_1(horizontal_tile_26_20_to_tile_26_19_1),
		.in_wire_0_2(horizontal_tile_26_20_to_tile_26_19_2),
		.in_wire_0_3(horizontal_tile_26_20_to_tile_26_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(852)
	);

	pe_tile pe_tile_26_20(
		.out_wire_3_0(vertical_tile_26_20_to_tile_25_20_0),
		.out_wire_3_1(vertical_tile_26_20_to_tile_25_20_1),
		.out_wire_3_2(vertical_tile_26_20_to_tile_25_20_2),
		.out_wire_3_3(vertical_tile_26_20_to_tile_25_20_3),
		.in_wire_3_0(vertical_tile_25_20_to_tile_26_20_0),
		.in_wire_3_1(vertical_tile_25_20_to_tile_26_20_1),
		.in_wire_3_2(vertical_tile_25_20_to_tile_26_20_2),
		.in_wire_3_3(vertical_tile_25_20_to_tile_26_20_3),
		.out_wire_1_0(vertical_tile_26_20_to_tile_27_20_0),
		.out_wire_1_1(vertical_tile_26_20_to_tile_27_20_1),
		.out_wire_1_2(vertical_tile_26_20_to_tile_27_20_2),
		.out_wire_1_3(vertical_tile_26_20_to_tile_27_20_3),
		.in_wire_1_0(vertical_tile_27_20_to_tile_26_20_0),
		.in_wire_1_1(vertical_tile_27_20_to_tile_26_20_1),
		.in_wire_1_2(vertical_tile_27_20_to_tile_26_20_2),
		.in_wire_1_3(vertical_tile_27_20_to_tile_26_20_3),
		.out_wire_2_0(horizontal_tile_26_20_to_tile_26_19_0),
		.out_wire_2_1(horizontal_tile_26_20_to_tile_26_19_1),
		.out_wire_2_2(horizontal_tile_26_20_to_tile_26_19_2),
		.out_wire_2_3(horizontal_tile_26_20_to_tile_26_19_3),
		.in_wire_2_0(horizontal_tile_26_19_to_tile_26_20_0),
		.in_wire_2_1(horizontal_tile_26_19_to_tile_26_20_1),
		.in_wire_2_2(horizontal_tile_26_19_to_tile_26_20_2),
		.in_wire_2_3(horizontal_tile_26_19_to_tile_26_20_3),
		.out_wire_0_0(horizontal_tile_26_20_to_tile_26_21_0),
		.out_wire_0_1(horizontal_tile_26_20_to_tile_26_21_1),
		.out_wire_0_2(horizontal_tile_26_20_to_tile_26_21_2),
		.out_wire_0_3(horizontal_tile_26_20_to_tile_26_21_3),
		.in_wire_0_0(horizontal_tile_26_21_to_tile_26_20_0),
		.in_wire_0_1(horizontal_tile_26_21_to_tile_26_20_1),
		.in_wire_0_2(horizontal_tile_26_21_to_tile_26_20_2),
		.in_wire_0_3(horizontal_tile_26_21_to_tile_26_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(853)
	);

	pe_tile pe_tile_26_21(
		.out_wire_3_0(vertical_tile_26_21_to_tile_25_21_0),
		.out_wire_3_1(vertical_tile_26_21_to_tile_25_21_1),
		.out_wire_3_2(vertical_tile_26_21_to_tile_25_21_2),
		.out_wire_3_3(vertical_tile_26_21_to_tile_25_21_3),
		.in_wire_3_0(vertical_tile_25_21_to_tile_26_21_0),
		.in_wire_3_1(vertical_tile_25_21_to_tile_26_21_1),
		.in_wire_3_2(vertical_tile_25_21_to_tile_26_21_2),
		.in_wire_3_3(vertical_tile_25_21_to_tile_26_21_3),
		.out_wire_1_0(vertical_tile_26_21_to_tile_27_21_0),
		.out_wire_1_1(vertical_tile_26_21_to_tile_27_21_1),
		.out_wire_1_2(vertical_tile_26_21_to_tile_27_21_2),
		.out_wire_1_3(vertical_tile_26_21_to_tile_27_21_3),
		.in_wire_1_0(vertical_tile_27_21_to_tile_26_21_0),
		.in_wire_1_1(vertical_tile_27_21_to_tile_26_21_1),
		.in_wire_1_2(vertical_tile_27_21_to_tile_26_21_2),
		.in_wire_1_3(vertical_tile_27_21_to_tile_26_21_3),
		.out_wire_2_0(horizontal_tile_26_21_to_tile_26_20_0),
		.out_wire_2_1(horizontal_tile_26_21_to_tile_26_20_1),
		.out_wire_2_2(horizontal_tile_26_21_to_tile_26_20_2),
		.out_wire_2_3(horizontal_tile_26_21_to_tile_26_20_3),
		.in_wire_2_0(horizontal_tile_26_20_to_tile_26_21_0),
		.in_wire_2_1(horizontal_tile_26_20_to_tile_26_21_1),
		.in_wire_2_2(horizontal_tile_26_20_to_tile_26_21_2),
		.in_wire_2_3(horizontal_tile_26_20_to_tile_26_21_3),
		.out_wire_0_0(horizontal_tile_26_21_to_tile_26_22_0),
		.out_wire_0_1(horizontal_tile_26_21_to_tile_26_22_1),
		.out_wire_0_2(horizontal_tile_26_21_to_tile_26_22_2),
		.out_wire_0_3(horizontal_tile_26_21_to_tile_26_22_3),
		.in_wire_0_0(horizontal_tile_26_22_to_tile_26_21_0),
		.in_wire_0_1(horizontal_tile_26_22_to_tile_26_21_1),
		.in_wire_0_2(horizontal_tile_26_22_to_tile_26_21_2),
		.in_wire_0_3(horizontal_tile_26_22_to_tile_26_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(854)
	);

	pe_tile pe_tile_26_22(
		.out_wire_3_0(vertical_tile_26_22_to_tile_25_22_0),
		.out_wire_3_1(vertical_tile_26_22_to_tile_25_22_1),
		.out_wire_3_2(vertical_tile_26_22_to_tile_25_22_2),
		.out_wire_3_3(vertical_tile_26_22_to_tile_25_22_3),
		.in_wire_3_0(vertical_tile_25_22_to_tile_26_22_0),
		.in_wire_3_1(vertical_tile_25_22_to_tile_26_22_1),
		.in_wire_3_2(vertical_tile_25_22_to_tile_26_22_2),
		.in_wire_3_3(vertical_tile_25_22_to_tile_26_22_3),
		.out_wire_1_0(vertical_tile_26_22_to_tile_27_22_0),
		.out_wire_1_1(vertical_tile_26_22_to_tile_27_22_1),
		.out_wire_1_2(vertical_tile_26_22_to_tile_27_22_2),
		.out_wire_1_3(vertical_tile_26_22_to_tile_27_22_3),
		.in_wire_1_0(vertical_tile_27_22_to_tile_26_22_0),
		.in_wire_1_1(vertical_tile_27_22_to_tile_26_22_1),
		.in_wire_1_2(vertical_tile_27_22_to_tile_26_22_2),
		.in_wire_1_3(vertical_tile_27_22_to_tile_26_22_3),
		.out_wire_2_0(horizontal_tile_26_22_to_tile_26_21_0),
		.out_wire_2_1(horizontal_tile_26_22_to_tile_26_21_1),
		.out_wire_2_2(horizontal_tile_26_22_to_tile_26_21_2),
		.out_wire_2_3(horizontal_tile_26_22_to_tile_26_21_3),
		.in_wire_2_0(horizontal_tile_26_21_to_tile_26_22_0),
		.in_wire_2_1(horizontal_tile_26_21_to_tile_26_22_1),
		.in_wire_2_2(horizontal_tile_26_21_to_tile_26_22_2),
		.in_wire_2_3(horizontal_tile_26_21_to_tile_26_22_3),
		.out_wire_0_0(horizontal_tile_26_22_to_tile_26_23_0),
		.out_wire_0_1(horizontal_tile_26_22_to_tile_26_23_1),
		.out_wire_0_2(horizontal_tile_26_22_to_tile_26_23_2),
		.out_wire_0_3(horizontal_tile_26_22_to_tile_26_23_3),
		.in_wire_0_0(horizontal_tile_26_23_to_tile_26_22_0),
		.in_wire_0_1(horizontal_tile_26_23_to_tile_26_22_1),
		.in_wire_0_2(horizontal_tile_26_23_to_tile_26_22_2),
		.in_wire_0_3(horizontal_tile_26_23_to_tile_26_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(855)
	);

	pe_tile pe_tile_26_23(
		.out_wire_3_0(vertical_tile_26_23_to_tile_25_23_0),
		.out_wire_3_1(vertical_tile_26_23_to_tile_25_23_1),
		.out_wire_3_2(vertical_tile_26_23_to_tile_25_23_2),
		.out_wire_3_3(vertical_tile_26_23_to_tile_25_23_3),
		.in_wire_3_0(vertical_tile_25_23_to_tile_26_23_0),
		.in_wire_3_1(vertical_tile_25_23_to_tile_26_23_1),
		.in_wire_3_2(vertical_tile_25_23_to_tile_26_23_2),
		.in_wire_3_3(vertical_tile_25_23_to_tile_26_23_3),
		.out_wire_1_0(vertical_tile_26_23_to_tile_27_23_0),
		.out_wire_1_1(vertical_tile_26_23_to_tile_27_23_1),
		.out_wire_1_2(vertical_tile_26_23_to_tile_27_23_2),
		.out_wire_1_3(vertical_tile_26_23_to_tile_27_23_3),
		.in_wire_1_0(vertical_tile_27_23_to_tile_26_23_0),
		.in_wire_1_1(vertical_tile_27_23_to_tile_26_23_1),
		.in_wire_1_2(vertical_tile_27_23_to_tile_26_23_2),
		.in_wire_1_3(vertical_tile_27_23_to_tile_26_23_3),
		.out_wire_2_0(horizontal_tile_26_23_to_tile_26_22_0),
		.out_wire_2_1(horizontal_tile_26_23_to_tile_26_22_1),
		.out_wire_2_2(horizontal_tile_26_23_to_tile_26_22_2),
		.out_wire_2_3(horizontal_tile_26_23_to_tile_26_22_3),
		.in_wire_2_0(horizontal_tile_26_22_to_tile_26_23_0),
		.in_wire_2_1(horizontal_tile_26_22_to_tile_26_23_1),
		.in_wire_2_2(horizontal_tile_26_22_to_tile_26_23_2),
		.in_wire_2_3(horizontal_tile_26_22_to_tile_26_23_3),
		.out_wire_0_0(horizontal_tile_26_23_to_tile_26_24_0),
		.out_wire_0_1(horizontal_tile_26_23_to_tile_26_24_1),
		.out_wire_0_2(horizontal_tile_26_23_to_tile_26_24_2),
		.out_wire_0_3(horizontal_tile_26_23_to_tile_26_24_3),
		.in_wire_0_0(horizontal_tile_26_24_to_tile_26_23_0),
		.in_wire_0_1(horizontal_tile_26_24_to_tile_26_23_1),
		.in_wire_0_2(horizontal_tile_26_24_to_tile_26_23_2),
		.in_wire_0_3(horizontal_tile_26_24_to_tile_26_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(856)
	);

	pe_tile pe_tile_26_24(
		.out_wire_3_0(vertical_tile_26_24_to_tile_25_24_0),
		.out_wire_3_1(vertical_tile_26_24_to_tile_25_24_1),
		.out_wire_3_2(vertical_tile_26_24_to_tile_25_24_2),
		.out_wire_3_3(vertical_tile_26_24_to_tile_25_24_3),
		.in_wire_3_0(vertical_tile_25_24_to_tile_26_24_0),
		.in_wire_3_1(vertical_tile_25_24_to_tile_26_24_1),
		.in_wire_3_2(vertical_tile_25_24_to_tile_26_24_2),
		.in_wire_3_3(vertical_tile_25_24_to_tile_26_24_3),
		.out_wire_1_0(vertical_tile_26_24_to_tile_27_24_0),
		.out_wire_1_1(vertical_tile_26_24_to_tile_27_24_1),
		.out_wire_1_2(vertical_tile_26_24_to_tile_27_24_2),
		.out_wire_1_3(vertical_tile_26_24_to_tile_27_24_3),
		.in_wire_1_0(vertical_tile_27_24_to_tile_26_24_0),
		.in_wire_1_1(vertical_tile_27_24_to_tile_26_24_1),
		.in_wire_1_2(vertical_tile_27_24_to_tile_26_24_2),
		.in_wire_1_3(vertical_tile_27_24_to_tile_26_24_3),
		.out_wire_2_0(horizontal_tile_26_24_to_tile_26_23_0),
		.out_wire_2_1(horizontal_tile_26_24_to_tile_26_23_1),
		.out_wire_2_2(horizontal_tile_26_24_to_tile_26_23_2),
		.out_wire_2_3(horizontal_tile_26_24_to_tile_26_23_3),
		.in_wire_2_0(horizontal_tile_26_23_to_tile_26_24_0),
		.in_wire_2_1(horizontal_tile_26_23_to_tile_26_24_1),
		.in_wire_2_2(horizontal_tile_26_23_to_tile_26_24_2),
		.in_wire_2_3(horizontal_tile_26_23_to_tile_26_24_3),
		.out_wire_0_0(horizontal_tile_26_24_to_tile_26_25_0),
		.out_wire_0_1(horizontal_tile_26_24_to_tile_26_25_1),
		.out_wire_0_2(horizontal_tile_26_24_to_tile_26_25_2),
		.out_wire_0_3(horizontal_tile_26_24_to_tile_26_25_3),
		.in_wire_0_0(horizontal_tile_26_25_to_tile_26_24_0),
		.in_wire_0_1(horizontal_tile_26_25_to_tile_26_24_1),
		.in_wire_0_2(horizontal_tile_26_25_to_tile_26_24_2),
		.in_wire_0_3(horizontal_tile_26_25_to_tile_26_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(857)
	);

	pe_tile pe_tile_26_25(
		.out_wire_3_0(vertical_tile_26_25_to_tile_25_25_0),
		.out_wire_3_1(vertical_tile_26_25_to_tile_25_25_1),
		.out_wire_3_2(vertical_tile_26_25_to_tile_25_25_2),
		.out_wire_3_3(vertical_tile_26_25_to_tile_25_25_3),
		.in_wire_3_0(vertical_tile_25_25_to_tile_26_25_0),
		.in_wire_3_1(vertical_tile_25_25_to_tile_26_25_1),
		.in_wire_3_2(vertical_tile_25_25_to_tile_26_25_2),
		.in_wire_3_3(vertical_tile_25_25_to_tile_26_25_3),
		.out_wire_1_0(vertical_tile_26_25_to_tile_27_25_0),
		.out_wire_1_1(vertical_tile_26_25_to_tile_27_25_1),
		.out_wire_1_2(vertical_tile_26_25_to_tile_27_25_2),
		.out_wire_1_3(vertical_tile_26_25_to_tile_27_25_3),
		.in_wire_1_0(vertical_tile_27_25_to_tile_26_25_0),
		.in_wire_1_1(vertical_tile_27_25_to_tile_26_25_1),
		.in_wire_1_2(vertical_tile_27_25_to_tile_26_25_2),
		.in_wire_1_3(vertical_tile_27_25_to_tile_26_25_3),
		.out_wire_2_0(horizontal_tile_26_25_to_tile_26_24_0),
		.out_wire_2_1(horizontal_tile_26_25_to_tile_26_24_1),
		.out_wire_2_2(horizontal_tile_26_25_to_tile_26_24_2),
		.out_wire_2_3(horizontal_tile_26_25_to_tile_26_24_3),
		.in_wire_2_0(horizontal_tile_26_24_to_tile_26_25_0),
		.in_wire_2_1(horizontal_tile_26_24_to_tile_26_25_1),
		.in_wire_2_2(horizontal_tile_26_24_to_tile_26_25_2),
		.in_wire_2_3(horizontal_tile_26_24_to_tile_26_25_3),
		.out_wire_0_0(horizontal_tile_26_25_to_tile_26_26_0),
		.out_wire_0_1(horizontal_tile_26_25_to_tile_26_26_1),
		.out_wire_0_2(horizontal_tile_26_25_to_tile_26_26_2),
		.out_wire_0_3(horizontal_tile_26_25_to_tile_26_26_3),
		.in_wire_0_0(horizontal_tile_26_26_to_tile_26_25_0),
		.in_wire_0_1(horizontal_tile_26_26_to_tile_26_25_1),
		.in_wire_0_2(horizontal_tile_26_26_to_tile_26_25_2),
		.in_wire_0_3(horizontal_tile_26_26_to_tile_26_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(858)
	);

	pe_tile pe_tile_26_26(
		.out_wire_3_0(vertical_tile_26_26_to_tile_25_26_0),
		.out_wire_3_1(vertical_tile_26_26_to_tile_25_26_1),
		.out_wire_3_2(vertical_tile_26_26_to_tile_25_26_2),
		.out_wire_3_3(vertical_tile_26_26_to_tile_25_26_3),
		.in_wire_3_0(vertical_tile_25_26_to_tile_26_26_0),
		.in_wire_3_1(vertical_tile_25_26_to_tile_26_26_1),
		.in_wire_3_2(vertical_tile_25_26_to_tile_26_26_2),
		.in_wire_3_3(vertical_tile_25_26_to_tile_26_26_3),
		.out_wire_1_0(vertical_tile_26_26_to_tile_27_26_0),
		.out_wire_1_1(vertical_tile_26_26_to_tile_27_26_1),
		.out_wire_1_2(vertical_tile_26_26_to_tile_27_26_2),
		.out_wire_1_3(vertical_tile_26_26_to_tile_27_26_3),
		.in_wire_1_0(vertical_tile_27_26_to_tile_26_26_0),
		.in_wire_1_1(vertical_tile_27_26_to_tile_26_26_1),
		.in_wire_1_2(vertical_tile_27_26_to_tile_26_26_2),
		.in_wire_1_3(vertical_tile_27_26_to_tile_26_26_3),
		.out_wire_2_0(horizontal_tile_26_26_to_tile_26_25_0),
		.out_wire_2_1(horizontal_tile_26_26_to_tile_26_25_1),
		.out_wire_2_2(horizontal_tile_26_26_to_tile_26_25_2),
		.out_wire_2_3(horizontal_tile_26_26_to_tile_26_25_3),
		.in_wire_2_0(horizontal_tile_26_25_to_tile_26_26_0),
		.in_wire_2_1(horizontal_tile_26_25_to_tile_26_26_1),
		.in_wire_2_2(horizontal_tile_26_25_to_tile_26_26_2),
		.in_wire_2_3(horizontal_tile_26_25_to_tile_26_26_3),
		.out_wire_0_0(horizontal_tile_26_26_to_tile_26_27_0),
		.out_wire_0_1(horizontal_tile_26_26_to_tile_26_27_1),
		.out_wire_0_2(horizontal_tile_26_26_to_tile_26_27_2),
		.out_wire_0_3(horizontal_tile_26_26_to_tile_26_27_3),
		.in_wire_0_0(horizontal_tile_26_27_to_tile_26_26_0),
		.in_wire_0_1(horizontal_tile_26_27_to_tile_26_26_1),
		.in_wire_0_2(horizontal_tile_26_27_to_tile_26_26_2),
		.in_wire_0_3(horizontal_tile_26_27_to_tile_26_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(859)
	);

	pe_tile pe_tile_26_27(
		.out_wire_3_0(vertical_tile_26_27_to_tile_25_27_0),
		.out_wire_3_1(vertical_tile_26_27_to_tile_25_27_1),
		.out_wire_3_2(vertical_tile_26_27_to_tile_25_27_2),
		.out_wire_3_3(vertical_tile_26_27_to_tile_25_27_3),
		.in_wire_3_0(vertical_tile_25_27_to_tile_26_27_0),
		.in_wire_3_1(vertical_tile_25_27_to_tile_26_27_1),
		.in_wire_3_2(vertical_tile_25_27_to_tile_26_27_2),
		.in_wire_3_3(vertical_tile_25_27_to_tile_26_27_3),
		.out_wire_1_0(vertical_tile_26_27_to_tile_27_27_0),
		.out_wire_1_1(vertical_tile_26_27_to_tile_27_27_1),
		.out_wire_1_2(vertical_tile_26_27_to_tile_27_27_2),
		.out_wire_1_3(vertical_tile_26_27_to_tile_27_27_3),
		.in_wire_1_0(vertical_tile_27_27_to_tile_26_27_0),
		.in_wire_1_1(vertical_tile_27_27_to_tile_26_27_1),
		.in_wire_1_2(vertical_tile_27_27_to_tile_26_27_2),
		.in_wire_1_3(vertical_tile_27_27_to_tile_26_27_3),
		.out_wire_2_0(horizontal_tile_26_27_to_tile_26_26_0),
		.out_wire_2_1(horizontal_tile_26_27_to_tile_26_26_1),
		.out_wire_2_2(horizontal_tile_26_27_to_tile_26_26_2),
		.out_wire_2_3(horizontal_tile_26_27_to_tile_26_26_3),
		.in_wire_2_0(horizontal_tile_26_26_to_tile_26_27_0),
		.in_wire_2_1(horizontal_tile_26_26_to_tile_26_27_1),
		.in_wire_2_2(horizontal_tile_26_26_to_tile_26_27_2),
		.in_wire_2_3(horizontal_tile_26_26_to_tile_26_27_3),
		.out_wire_0_0(horizontal_tile_26_27_to_tile_26_28_0),
		.out_wire_0_1(horizontal_tile_26_27_to_tile_26_28_1),
		.out_wire_0_2(horizontal_tile_26_27_to_tile_26_28_2),
		.out_wire_0_3(horizontal_tile_26_27_to_tile_26_28_3),
		.in_wire_0_0(horizontal_tile_26_28_to_tile_26_27_0),
		.in_wire_0_1(horizontal_tile_26_28_to_tile_26_27_1),
		.in_wire_0_2(horizontal_tile_26_28_to_tile_26_27_2),
		.in_wire_0_3(horizontal_tile_26_28_to_tile_26_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(860)
	);

	pe_tile pe_tile_26_28(
		.out_wire_3_0(vertical_tile_26_28_to_tile_25_28_0),
		.out_wire_3_1(vertical_tile_26_28_to_tile_25_28_1),
		.out_wire_3_2(vertical_tile_26_28_to_tile_25_28_2),
		.out_wire_3_3(vertical_tile_26_28_to_tile_25_28_3),
		.in_wire_3_0(vertical_tile_25_28_to_tile_26_28_0),
		.in_wire_3_1(vertical_tile_25_28_to_tile_26_28_1),
		.in_wire_3_2(vertical_tile_25_28_to_tile_26_28_2),
		.in_wire_3_3(vertical_tile_25_28_to_tile_26_28_3),
		.out_wire_1_0(vertical_tile_26_28_to_tile_27_28_0),
		.out_wire_1_1(vertical_tile_26_28_to_tile_27_28_1),
		.out_wire_1_2(vertical_tile_26_28_to_tile_27_28_2),
		.out_wire_1_3(vertical_tile_26_28_to_tile_27_28_3),
		.in_wire_1_0(vertical_tile_27_28_to_tile_26_28_0),
		.in_wire_1_1(vertical_tile_27_28_to_tile_26_28_1),
		.in_wire_1_2(vertical_tile_27_28_to_tile_26_28_2),
		.in_wire_1_3(vertical_tile_27_28_to_tile_26_28_3),
		.out_wire_2_0(horizontal_tile_26_28_to_tile_26_27_0),
		.out_wire_2_1(horizontal_tile_26_28_to_tile_26_27_1),
		.out_wire_2_2(horizontal_tile_26_28_to_tile_26_27_2),
		.out_wire_2_3(horizontal_tile_26_28_to_tile_26_27_3),
		.in_wire_2_0(horizontal_tile_26_27_to_tile_26_28_0),
		.in_wire_2_1(horizontal_tile_26_27_to_tile_26_28_1),
		.in_wire_2_2(horizontal_tile_26_27_to_tile_26_28_2),
		.in_wire_2_3(horizontal_tile_26_27_to_tile_26_28_3),
		.out_wire_0_0(horizontal_tile_26_28_to_tile_26_29_0),
		.out_wire_0_1(horizontal_tile_26_28_to_tile_26_29_1),
		.out_wire_0_2(horizontal_tile_26_28_to_tile_26_29_2),
		.out_wire_0_3(horizontal_tile_26_28_to_tile_26_29_3),
		.in_wire_0_0(horizontal_tile_26_29_to_tile_26_28_0),
		.in_wire_0_1(horizontal_tile_26_29_to_tile_26_28_1),
		.in_wire_0_2(horizontal_tile_26_29_to_tile_26_28_2),
		.in_wire_0_3(horizontal_tile_26_29_to_tile_26_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(861)
	);

	pe_tile pe_tile_26_29(
		.out_wire_3_0(vertical_tile_26_29_to_tile_25_29_0),
		.out_wire_3_1(vertical_tile_26_29_to_tile_25_29_1),
		.out_wire_3_2(vertical_tile_26_29_to_tile_25_29_2),
		.out_wire_3_3(vertical_tile_26_29_to_tile_25_29_3),
		.in_wire_3_0(vertical_tile_25_29_to_tile_26_29_0),
		.in_wire_3_1(vertical_tile_25_29_to_tile_26_29_1),
		.in_wire_3_2(vertical_tile_25_29_to_tile_26_29_2),
		.in_wire_3_3(vertical_tile_25_29_to_tile_26_29_3),
		.out_wire_1_0(vertical_tile_26_29_to_tile_27_29_0),
		.out_wire_1_1(vertical_tile_26_29_to_tile_27_29_1),
		.out_wire_1_2(vertical_tile_26_29_to_tile_27_29_2),
		.out_wire_1_3(vertical_tile_26_29_to_tile_27_29_3),
		.in_wire_1_0(vertical_tile_27_29_to_tile_26_29_0),
		.in_wire_1_1(vertical_tile_27_29_to_tile_26_29_1),
		.in_wire_1_2(vertical_tile_27_29_to_tile_26_29_2),
		.in_wire_1_3(vertical_tile_27_29_to_tile_26_29_3),
		.out_wire_2_0(horizontal_tile_26_29_to_tile_26_28_0),
		.out_wire_2_1(horizontal_tile_26_29_to_tile_26_28_1),
		.out_wire_2_2(horizontal_tile_26_29_to_tile_26_28_2),
		.out_wire_2_3(horizontal_tile_26_29_to_tile_26_28_3),
		.in_wire_2_0(horizontal_tile_26_28_to_tile_26_29_0),
		.in_wire_2_1(horizontal_tile_26_28_to_tile_26_29_1),
		.in_wire_2_2(horizontal_tile_26_28_to_tile_26_29_2),
		.in_wire_2_3(horizontal_tile_26_28_to_tile_26_29_3),
		.out_wire_0_0(horizontal_tile_26_29_to_tile_26_30_0),
		.out_wire_0_1(horizontal_tile_26_29_to_tile_26_30_1),
		.out_wire_0_2(horizontal_tile_26_29_to_tile_26_30_2),
		.out_wire_0_3(horizontal_tile_26_29_to_tile_26_30_3),
		.in_wire_0_0(horizontal_tile_26_30_to_tile_26_29_0),
		.in_wire_0_1(horizontal_tile_26_30_to_tile_26_29_1),
		.in_wire_0_2(horizontal_tile_26_30_to_tile_26_29_2),
		.in_wire_0_3(horizontal_tile_26_30_to_tile_26_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(862)
	);

	pe_tile pe_tile_26_30(
		.out_wire_3_0(vertical_tile_26_30_to_tile_25_30_0),
		.out_wire_3_1(vertical_tile_26_30_to_tile_25_30_1),
		.out_wire_3_2(vertical_tile_26_30_to_tile_25_30_2),
		.out_wire_3_3(vertical_tile_26_30_to_tile_25_30_3),
		.in_wire_3_0(vertical_tile_25_30_to_tile_26_30_0),
		.in_wire_3_1(vertical_tile_25_30_to_tile_26_30_1),
		.in_wire_3_2(vertical_tile_25_30_to_tile_26_30_2),
		.in_wire_3_3(vertical_tile_25_30_to_tile_26_30_3),
		.out_wire_1_0(vertical_tile_26_30_to_tile_27_30_0),
		.out_wire_1_1(vertical_tile_26_30_to_tile_27_30_1),
		.out_wire_1_2(vertical_tile_26_30_to_tile_27_30_2),
		.out_wire_1_3(vertical_tile_26_30_to_tile_27_30_3),
		.in_wire_1_0(vertical_tile_27_30_to_tile_26_30_0),
		.in_wire_1_1(vertical_tile_27_30_to_tile_26_30_1),
		.in_wire_1_2(vertical_tile_27_30_to_tile_26_30_2),
		.in_wire_1_3(vertical_tile_27_30_to_tile_26_30_3),
		.out_wire_2_0(horizontal_tile_26_30_to_tile_26_29_0),
		.out_wire_2_1(horizontal_tile_26_30_to_tile_26_29_1),
		.out_wire_2_2(horizontal_tile_26_30_to_tile_26_29_2),
		.out_wire_2_3(horizontal_tile_26_30_to_tile_26_29_3),
		.in_wire_2_0(horizontal_tile_26_29_to_tile_26_30_0),
		.in_wire_2_1(horizontal_tile_26_29_to_tile_26_30_1),
		.in_wire_2_2(horizontal_tile_26_29_to_tile_26_30_2),
		.in_wire_2_3(horizontal_tile_26_29_to_tile_26_30_3),
		.out_wire_0_0(horizontal_tile_26_30_to_tile_26_31_0),
		.out_wire_0_1(horizontal_tile_26_30_to_tile_26_31_1),
		.out_wire_0_2(horizontal_tile_26_30_to_tile_26_31_2),
		.out_wire_0_3(horizontal_tile_26_30_to_tile_26_31_3),
		.in_wire_0_0(horizontal_tile_26_31_to_tile_26_30_0),
		.in_wire_0_1(horizontal_tile_26_31_to_tile_26_30_1),
		.in_wire_0_2(horizontal_tile_26_31_to_tile_26_30_2),
		.in_wire_0_3(horizontal_tile_26_31_to_tile_26_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(863)
	);

	pe_tile_right pe_tile_26_31(
		.out_wire_3_0(vertical_tile_26_31_to_tile_25_31_0),
		.out_wire_3_1(vertical_tile_26_31_to_tile_25_31_1),
		.out_wire_3_2(vertical_tile_26_31_to_tile_25_31_2),
		.out_wire_3_3(vertical_tile_26_31_to_tile_25_31_3),
		.in_wire_3_0(vertical_tile_25_31_to_tile_26_31_0),
		.in_wire_3_1(vertical_tile_25_31_to_tile_26_31_1),
		.in_wire_3_2(vertical_tile_25_31_to_tile_26_31_2),
		.in_wire_3_3(vertical_tile_25_31_to_tile_26_31_3),
		.out_wire_1_0(vertical_tile_26_31_to_tile_27_31_0),
		.out_wire_1_1(vertical_tile_26_31_to_tile_27_31_1),
		.out_wire_1_2(vertical_tile_26_31_to_tile_27_31_2),
		.out_wire_1_3(vertical_tile_26_31_to_tile_27_31_3),
		.in_wire_1_0(vertical_tile_27_31_to_tile_26_31_0),
		.in_wire_1_1(vertical_tile_27_31_to_tile_26_31_1),
		.in_wire_1_2(vertical_tile_27_31_to_tile_26_31_2),
		.in_wire_1_3(vertical_tile_27_31_to_tile_26_31_3),
		.out_wire_2_0(horizontal_tile_26_31_to_tile_26_30_0),
		.out_wire_2_1(horizontal_tile_26_31_to_tile_26_30_1),
		.out_wire_2_2(horizontal_tile_26_31_to_tile_26_30_2),
		.out_wire_2_3(horizontal_tile_26_31_to_tile_26_30_3),
		.in_wire_2_0(horizontal_tile_26_30_to_tile_26_31_0),
		.in_wire_2_1(horizontal_tile_26_30_to_tile_26_31_1),
		.in_wire_2_2(horizontal_tile_26_30_to_tile_26_31_2),
		.in_wire_2_3(horizontal_tile_26_30_to_tile_26_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(864)
	);

	pe_tile_left pe_tile_27_0(
		.out_wire_3_0(vertical_tile_27_0_to_tile_26_0_0),
		.out_wire_3_1(vertical_tile_27_0_to_tile_26_0_1),
		.out_wire_3_2(vertical_tile_27_0_to_tile_26_0_2),
		.out_wire_3_3(vertical_tile_27_0_to_tile_26_0_3),
		.in_wire_3_0(vertical_tile_26_0_to_tile_27_0_0),
		.in_wire_3_1(vertical_tile_26_0_to_tile_27_0_1),
		.in_wire_3_2(vertical_tile_26_0_to_tile_27_0_2),
		.in_wire_3_3(vertical_tile_26_0_to_tile_27_0_3),
		.out_wire_1_0(vertical_tile_27_0_to_tile_28_0_0),
		.out_wire_1_1(vertical_tile_27_0_to_tile_28_0_1),
		.out_wire_1_2(vertical_tile_27_0_to_tile_28_0_2),
		.out_wire_1_3(vertical_tile_27_0_to_tile_28_0_3),
		.in_wire_1_0(vertical_tile_28_0_to_tile_27_0_0),
		.in_wire_1_1(vertical_tile_28_0_to_tile_27_0_1),
		.in_wire_1_2(vertical_tile_28_0_to_tile_27_0_2),
		.in_wire_1_3(vertical_tile_28_0_to_tile_27_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_27_0_to_tile_27_1_0),
		.out_wire_0_1(horizontal_tile_27_0_to_tile_27_1_1),
		.out_wire_0_2(horizontal_tile_27_0_to_tile_27_1_2),
		.out_wire_0_3(horizontal_tile_27_0_to_tile_27_1_3),
		.in_wire_0_0(horizontal_tile_27_1_to_tile_27_0_0),
		.in_wire_0_1(horizontal_tile_27_1_to_tile_27_0_1),
		.in_wire_0_2(horizontal_tile_27_1_to_tile_27_0_2),
		.in_wire_0_3(horizontal_tile_27_1_to_tile_27_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(865)
	);

	pe_tile pe_tile_27_1(
		.out_wire_3_0(vertical_tile_27_1_to_tile_26_1_0),
		.out_wire_3_1(vertical_tile_27_1_to_tile_26_1_1),
		.out_wire_3_2(vertical_tile_27_1_to_tile_26_1_2),
		.out_wire_3_3(vertical_tile_27_1_to_tile_26_1_3),
		.in_wire_3_0(vertical_tile_26_1_to_tile_27_1_0),
		.in_wire_3_1(vertical_tile_26_1_to_tile_27_1_1),
		.in_wire_3_2(vertical_tile_26_1_to_tile_27_1_2),
		.in_wire_3_3(vertical_tile_26_1_to_tile_27_1_3),
		.out_wire_1_0(vertical_tile_27_1_to_tile_28_1_0),
		.out_wire_1_1(vertical_tile_27_1_to_tile_28_1_1),
		.out_wire_1_2(vertical_tile_27_1_to_tile_28_1_2),
		.out_wire_1_3(vertical_tile_27_1_to_tile_28_1_3),
		.in_wire_1_0(vertical_tile_28_1_to_tile_27_1_0),
		.in_wire_1_1(vertical_tile_28_1_to_tile_27_1_1),
		.in_wire_1_2(vertical_tile_28_1_to_tile_27_1_2),
		.in_wire_1_3(vertical_tile_28_1_to_tile_27_1_3),
		.out_wire_2_0(horizontal_tile_27_1_to_tile_27_0_0),
		.out_wire_2_1(horizontal_tile_27_1_to_tile_27_0_1),
		.out_wire_2_2(horizontal_tile_27_1_to_tile_27_0_2),
		.out_wire_2_3(horizontal_tile_27_1_to_tile_27_0_3),
		.in_wire_2_0(horizontal_tile_27_0_to_tile_27_1_0),
		.in_wire_2_1(horizontal_tile_27_0_to_tile_27_1_1),
		.in_wire_2_2(horizontal_tile_27_0_to_tile_27_1_2),
		.in_wire_2_3(horizontal_tile_27_0_to_tile_27_1_3),
		.out_wire_0_0(horizontal_tile_27_1_to_tile_27_2_0),
		.out_wire_0_1(horizontal_tile_27_1_to_tile_27_2_1),
		.out_wire_0_2(horizontal_tile_27_1_to_tile_27_2_2),
		.out_wire_0_3(horizontal_tile_27_1_to_tile_27_2_3),
		.in_wire_0_0(horizontal_tile_27_2_to_tile_27_1_0),
		.in_wire_0_1(horizontal_tile_27_2_to_tile_27_1_1),
		.in_wire_0_2(horizontal_tile_27_2_to_tile_27_1_2),
		.in_wire_0_3(horizontal_tile_27_2_to_tile_27_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(866)
	);

	pe_tile pe_tile_27_2(
		.out_wire_3_0(vertical_tile_27_2_to_tile_26_2_0),
		.out_wire_3_1(vertical_tile_27_2_to_tile_26_2_1),
		.out_wire_3_2(vertical_tile_27_2_to_tile_26_2_2),
		.out_wire_3_3(vertical_tile_27_2_to_tile_26_2_3),
		.in_wire_3_0(vertical_tile_26_2_to_tile_27_2_0),
		.in_wire_3_1(vertical_tile_26_2_to_tile_27_2_1),
		.in_wire_3_2(vertical_tile_26_2_to_tile_27_2_2),
		.in_wire_3_3(vertical_tile_26_2_to_tile_27_2_3),
		.out_wire_1_0(vertical_tile_27_2_to_tile_28_2_0),
		.out_wire_1_1(vertical_tile_27_2_to_tile_28_2_1),
		.out_wire_1_2(vertical_tile_27_2_to_tile_28_2_2),
		.out_wire_1_3(vertical_tile_27_2_to_tile_28_2_3),
		.in_wire_1_0(vertical_tile_28_2_to_tile_27_2_0),
		.in_wire_1_1(vertical_tile_28_2_to_tile_27_2_1),
		.in_wire_1_2(vertical_tile_28_2_to_tile_27_2_2),
		.in_wire_1_3(vertical_tile_28_2_to_tile_27_2_3),
		.out_wire_2_0(horizontal_tile_27_2_to_tile_27_1_0),
		.out_wire_2_1(horizontal_tile_27_2_to_tile_27_1_1),
		.out_wire_2_2(horizontal_tile_27_2_to_tile_27_1_2),
		.out_wire_2_3(horizontal_tile_27_2_to_tile_27_1_3),
		.in_wire_2_0(horizontal_tile_27_1_to_tile_27_2_0),
		.in_wire_2_1(horizontal_tile_27_1_to_tile_27_2_1),
		.in_wire_2_2(horizontal_tile_27_1_to_tile_27_2_2),
		.in_wire_2_3(horizontal_tile_27_1_to_tile_27_2_3),
		.out_wire_0_0(horizontal_tile_27_2_to_tile_27_3_0),
		.out_wire_0_1(horizontal_tile_27_2_to_tile_27_3_1),
		.out_wire_0_2(horizontal_tile_27_2_to_tile_27_3_2),
		.out_wire_0_3(horizontal_tile_27_2_to_tile_27_3_3),
		.in_wire_0_0(horizontal_tile_27_3_to_tile_27_2_0),
		.in_wire_0_1(horizontal_tile_27_3_to_tile_27_2_1),
		.in_wire_0_2(horizontal_tile_27_3_to_tile_27_2_2),
		.in_wire_0_3(horizontal_tile_27_3_to_tile_27_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(867)
	);

	pe_tile pe_tile_27_3(
		.out_wire_3_0(vertical_tile_27_3_to_tile_26_3_0),
		.out_wire_3_1(vertical_tile_27_3_to_tile_26_3_1),
		.out_wire_3_2(vertical_tile_27_3_to_tile_26_3_2),
		.out_wire_3_3(vertical_tile_27_3_to_tile_26_3_3),
		.in_wire_3_0(vertical_tile_26_3_to_tile_27_3_0),
		.in_wire_3_1(vertical_tile_26_3_to_tile_27_3_1),
		.in_wire_3_2(vertical_tile_26_3_to_tile_27_3_2),
		.in_wire_3_3(vertical_tile_26_3_to_tile_27_3_3),
		.out_wire_1_0(vertical_tile_27_3_to_tile_28_3_0),
		.out_wire_1_1(vertical_tile_27_3_to_tile_28_3_1),
		.out_wire_1_2(vertical_tile_27_3_to_tile_28_3_2),
		.out_wire_1_3(vertical_tile_27_3_to_tile_28_3_3),
		.in_wire_1_0(vertical_tile_28_3_to_tile_27_3_0),
		.in_wire_1_1(vertical_tile_28_3_to_tile_27_3_1),
		.in_wire_1_2(vertical_tile_28_3_to_tile_27_3_2),
		.in_wire_1_3(vertical_tile_28_3_to_tile_27_3_3),
		.out_wire_2_0(horizontal_tile_27_3_to_tile_27_2_0),
		.out_wire_2_1(horizontal_tile_27_3_to_tile_27_2_1),
		.out_wire_2_2(horizontal_tile_27_3_to_tile_27_2_2),
		.out_wire_2_3(horizontal_tile_27_3_to_tile_27_2_3),
		.in_wire_2_0(horizontal_tile_27_2_to_tile_27_3_0),
		.in_wire_2_1(horizontal_tile_27_2_to_tile_27_3_1),
		.in_wire_2_2(horizontal_tile_27_2_to_tile_27_3_2),
		.in_wire_2_3(horizontal_tile_27_2_to_tile_27_3_3),
		.out_wire_0_0(horizontal_tile_27_3_to_tile_27_4_0),
		.out_wire_0_1(horizontal_tile_27_3_to_tile_27_4_1),
		.out_wire_0_2(horizontal_tile_27_3_to_tile_27_4_2),
		.out_wire_0_3(horizontal_tile_27_3_to_tile_27_4_3),
		.in_wire_0_0(horizontal_tile_27_4_to_tile_27_3_0),
		.in_wire_0_1(horizontal_tile_27_4_to_tile_27_3_1),
		.in_wire_0_2(horizontal_tile_27_4_to_tile_27_3_2),
		.in_wire_0_3(horizontal_tile_27_4_to_tile_27_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(868)
	);

	pe_tile pe_tile_27_4(
		.out_wire_3_0(vertical_tile_27_4_to_tile_26_4_0),
		.out_wire_3_1(vertical_tile_27_4_to_tile_26_4_1),
		.out_wire_3_2(vertical_tile_27_4_to_tile_26_4_2),
		.out_wire_3_3(vertical_tile_27_4_to_tile_26_4_3),
		.in_wire_3_0(vertical_tile_26_4_to_tile_27_4_0),
		.in_wire_3_1(vertical_tile_26_4_to_tile_27_4_1),
		.in_wire_3_2(vertical_tile_26_4_to_tile_27_4_2),
		.in_wire_3_3(vertical_tile_26_4_to_tile_27_4_3),
		.out_wire_1_0(vertical_tile_27_4_to_tile_28_4_0),
		.out_wire_1_1(vertical_tile_27_4_to_tile_28_4_1),
		.out_wire_1_2(vertical_tile_27_4_to_tile_28_4_2),
		.out_wire_1_3(vertical_tile_27_4_to_tile_28_4_3),
		.in_wire_1_0(vertical_tile_28_4_to_tile_27_4_0),
		.in_wire_1_1(vertical_tile_28_4_to_tile_27_4_1),
		.in_wire_1_2(vertical_tile_28_4_to_tile_27_4_2),
		.in_wire_1_3(vertical_tile_28_4_to_tile_27_4_3),
		.out_wire_2_0(horizontal_tile_27_4_to_tile_27_3_0),
		.out_wire_2_1(horizontal_tile_27_4_to_tile_27_3_1),
		.out_wire_2_2(horizontal_tile_27_4_to_tile_27_3_2),
		.out_wire_2_3(horizontal_tile_27_4_to_tile_27_3_3),
		.in_wire_2_0(horizontal_tile_27_3_to_tile_27_4_0),
		.in_wire_2_1(horizontal_tile_27_3_to_tile_27_4_1),
		.in_wire_2_2(horizontal_tile_27_3_to_tile_27_4_2),
		.in_wire_2_3(horizontal_tile_27_3_to_tile_27_4_3),
		.out_wire_0_0(horizontal_tile_27_4_to_tile_27_5_0),
		.out_wire_0_1(horizontal_tile_27_4_to_tile_27_5_1),
		.out_wire_0_2(horizontal_tile_27_4_to_tile_27_5_2),
		.out_wire_0_3(horizontal_tile_27_4_to_tile_27_5_3),
		.in_wire_0_0(horizontal_tile_27_5_to_tile_27_4_0),
		.in_wire_0_1(horizontal_tile_27_5_to_tile_27_4_1),
		.in_wire_0_2(horizontal_tile_27_5_to_tile_27_4_2),
		.in_wire_0_3(horizontal_tile_27_5_to_tile_27_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(869)
	);

	pe_tile pe_tile_27_5(
		.out_wire_3_0(vertical_tile_27_5_to_tile_26_5_0),
		.out_wire_3_1(vertical_tile_27_5_to_tile_26_5_1),
		.out_wire_3_2(vertical_tile_27_5_to_tile_26_5_2),
		.out_wire_3_3(vertical_tile_27_5_to_tile_26_5_3),
		.in_wire_3_0(vertical_tile_26_5_to_tile_27_5_0),
		.in_wire_3_1(vertical_tile_26_5_to_tile_27_5_1),
		.in_wire_3_2(vertical_tile_26_5_to_tile_27_5_2),
		.in_wire_3_3(vertical_tile_26_5_to_tile_27_5_3),
		.out_wire_1_0(vertical_tile_27_5_to_tile_28_5_0),
		.out_wire_1_1(vertical_tile_27_5_to_tile_28_5_1),
		.out_wire_1_2(vertical_tile_27_5_to_tile_28_5_2),
		.out_wire_1_3(vertical_tile_27_5_to_tile_28_5_3),
		.in_wire_1_0(vertical_tile_28_5_to_tile_27_5_0),
		.in_wire_1_1(vertical_tile_28_5_to_tile_27_5_1),
		.in_wire_1_2(vertical_tile_28_5_to_tile_27_5_2),
		.in_wire_1_3(vertical_tile_28_5_to_tile_27_5_3),
		.out_wire_2_0(horizontal_tile_27_5_to_tile_27_4_0),
		.out_wire_2_1(horizontal_tile_27_5_to_tile_27_4_1),
		.out_wire_2_2(horizontal_tile_27_5_to_tile_27_4_2),
		.out_wire_2_3(horizontal_tile_27_5_to_tile_27_4_3),
		.in_wire_2_0(horizontal_tile_27_4_to_tile_27_5_0),
		.in_wire_2_1(horizontal_tile_27_4_to_tile_27_5_1),
		.in_wire_2_2(horizontal_tile_27_4_to_tile_27_5_2),
		.in_wire_2_3(horizontal_tile_27_4_to_tile_27_5_3),
		.out_wire_0_0(horizontal_tile_27_5_to_tile_27_6_0),
		.out_wire_0_1(horizontal_tile_27_5_to_tile_27_6_1),
		.out_wire_0_2(horizontal_tile_27_5_to_tile_27_6_2),
		.out_wire_0_3(horizontal_tile_27_5_to_tile_27_6_3),
		.in_wire_0_0(horizontal_tile_27_6_to_tile_27_5_0),
		.in_wire_0_1(horizontal_tile_27_6_to_tile_27_5_1),
		.in_wire_0_2(horizontal_tile_27_6_to_tile_27_5_2),
		.in_wire_0_3(horizontal_tile_27_6_to_tile_27_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(870)
	);

	pe_tile pe_tile_27_6(
		.out_wire_3_0(vertical_tile_27_6_to_tile_26_6_0),
		.out_wire_3_1(vertical_tile_27_6_to_tile_26_6_1),
		.out_wire_3_2(vertical_tile_27_6_to_tile_26_6_2),
		.out_wire_3_3(vertical_tile_27_6_to_tile_26_6_3),
		.in_wire_3_0(vertical_tile_26_6_to_tile_27_6_0),
		.in_wire_3_1(vertical_tile_26_6_to_tile_27_6_1),
		.in_wire_3_2(vertical_tile_26_6_to_tile_27_6_2),
		.in_wire_3_3(vertical_tile_26_6_to_tile_27_6_3),
		.out_wire_1_0(vertical_tile_27_6_to_tile_28_6_0),
		.out_wire_1_1(vertical_tile_27_6_to_tile_28_6_1),
		.out_wire_1_2(vertical_tile_27_6_to_tile_28_6_2),
		.out_wire_1_3(vertical_tile_27_6_to_tile_28_6_3),
		.in_wire_1_0(vertical_tile_28_6_to_tile_27_6_0),
		.in_wire_1_1(vertical_tile_28_6_to_tile_27_6_1),
		.in_wire_1_2(vertical_tile_28_6_to_tile_27_6_2),
		.in_wire_1_3(vertical_tile_28_6_to_tile_27_6_3),
		.out_wire_2_0(horizontal_tile_27_6_to_tile_27_5_0),
		.out_wire_2_1(horizontal_tile_27_6_to_tile_27_5_1),
		.out_wire_2_2(horizontal_tile_27_6_to_tile_27_5_2),
		.out_wire_2_3(horizontal_tile_27_6_to_tile_27_5_3),
		.in_wire_2_0(horizontal_tile_27_5_to_tile_27_6_0),
		.in_wire_2_1(horizontal_tile_27_5_to_tile_27_6_1),
		.in_wire_2_2(horizontal_tile_27_5_to_tile_27_6_2),
		.in_wire_2_3(horizontal_tile_27_5_to_tile_27_6_3),
		.out_wire_0_0(horizontal_tile_27_6_to_tile_27_7_0),
		.out_wire_0_1(horizontal_tile_27_6_to_tile_27_7_1),
		.out_wire_0_2(horizontal_tile_27_6_to_tile_27_7_2),
		.out_wire_0_3(horizontal_tile_27_6_to_tile_27_7_3),
		.in_wire_0_0(horizontal_tile_27_7_to_tile_27_6_0),
		.in_wire_0_1(horizontal_tile_27_7_to_tile_27_6_1),
		.in_wire_0_2(horizontal_tile_27_7_to_tile_27_6_2),
		.in_wire_0_3(horizontal_tile_27_7_to_tile_27_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(871)
	);

	pe_tile pe_tile_27_7(
		.out_wire_3_0(vertical_tile_27_7_to_tile_26_7_0),
		.out_wire_3_1(vertical_tile_27_7_to_tile_26_7_1),
		.out_wire_3_2(vertical_tile_27_7_to_tile_26_7_2),
		.out_wire_3_3(vertical_tile_27_7_to_tile_26_7_3),
		.in_wire_3_0(vertical_tile_26_7_to_tile_27_7_0),
		.in_wire_3_1(vertical_tile_26_7_to_tile_27_7_1),
		.in_wire_3_2(vertical_tile_26_7_to_tile_27_7_2),
		.in_wire_3_3(vertical_tile_26_7_to_tile_27_7_3),
		.out_wire_1_0(vertical_tile_27_7_to_tile_28_7_0),
		.out_wire_1_1(vertical_tile_27_7_to_tile_28_7_1),
		.out_wire_1_2(vertical_tile_27_7_to_tile_28_7_2),
		.out_wire_1_3(vertical_tile_27_7_to_tile_28_7_3),
		.in_wire_1_0(vertical_tile_28_7_to_tile_27_7_0),
		.in_wire_1_1(vertical_tile_28_7_to_tile_27_7_1),
		.in_wire_1_2(vertical_tile_28_7_to_tile_27_7_2),
		.in_wire_1_3(vertical_tile_28_7_to_tile_27_7_3),
		.out_wire_2_0(horizontal_tile_27_7_to_tile_27_6_0),
		.out_wire_2_1(horizontal_tile_27_7_to_tile_27_6_1),
		.out_wire_2_2(horizontal_tile_27_7_to_tile_27_6_2),
		.out_wire_2_3(horizontal_tile_27_7_to_tile_27_6_3),
		.in_wire_2_0(horizontal_tile_27_6_to_tile_27_7_0),
		.in_wire_2_1(horizontal_tile_27_6_to_tile_27_7_1),
		.in_wire_2_2(horizontal_tile_27_6_to_tile_27_7_2),
		.in_wire_2_3(horizontal_tile_27_6_to_tile_27_7_3),
		.out_wire_0_0(horizontal_tile_27_7_to_tile_27_8_0),
		.out_wire_0_1(horizontal_tile_27_7_to_tile_27_8_1),
		.out_wire_0_2(horizontal_tile_27_7_to_tile_27_8_2),
		.out_wire_0_3(horizontal_tile_27_7_to_tile_27_8_3),
		.in_wire_0_0(horizontal_tile_27_8_to_tile_27_7_0),
		.in_wire_0_1(horizontal_tile_27_8_to_tile_27_7_1),
		.in_wire_0_2(horizontal_tile_27_8_to_tile_27_7_2),
		.in_wire_0_3(horizontal_tile_27_8_to_tile_27_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(872)
	);

	pe_tile pe_tile_27_8(
		.out_wire_3_0(vertical_tile_27_8_to_tile_26_8_0),
		.out_wire_3_1(vertical_tile_27_8_to_tile_26_8_1),
		.out_wire_3_2(vertical_tile_27_8_to_tile_26_8_2),
		.out_wire_3_3(vertical_tile_27_8_to_tile_26_8_3),
		.in_wire_3_0(vertical_tile_26_8_to_tile_27_8_0),
		.in_wire_3_1(vertical_tile_26_8_to_tile_27_8_1),
		.in_wire_3_2(vertical_tile_26_8_to_tile_27_8_2),
		.in_wire_3_3(vertical_tile_26_8_to_tile_27_8_3),
		.out_wire_1_0(vertical_tile_27_8_to_tile_28_8_0),
		.out_wire_1_1(vertical_tile_27_8_to_tile_28_8_1),
		.out_wire_1_2(vertical_tile_27_8_to_tile_28_8_2),
		.out_wire_1_3(vertical_tile_27_8_to_tile_28_8_3),
		.in_wire_1_0(vertical_tile_28_8_to_tile_27_8_0),
		.in_wire_1_1(vertical_tile_28_8_to_tile_27_8_1),
		.in_wire_1_2(vertical_tile_28_8_to_tile_27_8_2),
		.in_wire_1_3(vertical_tile_28_8_to_tile_27_8_3),
		.out_wire_2_0(horizontal_tile_27_8_to_tile_27_7_0),
		.out_wire_2_1(horizontal_tile_27_8_to_tile_27_7_1),
		.out_wire_2_2(horizontal_tile_27_8_to_tile_27_7_2),
		.out_wire_2_3(horizontal_tile_27_8_to_tile_27_7_3),
		.in_wire_2_0(horizontal_tile_27_7_to_tile_27_8_0),
		.in_wire_2_1(horizontal_tile_27_7_to_tile_27_8_1),
		.in_wire_2_2(horizontal_tile_27_7_to_tile_27_8_2),
		.in_wire_2_3(horizontal_tile_27_7_to_tile_27_8_3),
		.out_wire_0_0(horizontal_tile_27_8_to_tile_27_9_0),
		.out_wire_0_1(horizontal_tile_27_8_to_tile_27_9_1),
		.out_wire_0_2(horizontal_tile_27_8_to_tile_27_9_2),
		.out_wire_0_3(horizontal_tile_27_8_to_tile_27_9_3),
		.in_wire_0_0(horizontal_tile_27_9_to_tile_27_8_0),
		.in_wire_0_1(horizontal_tile_27_9_to_tile_27_8_1),
		.in_wire_0_2(horizontal_tile_27_9_to_tile_27_8_2),
		.in_wire_0_3(horizontal_tile_27_9_to_tile_27_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(873)
	);

	pe_tile pe_tile_27_9(
		.out_wire_3_0(vertical_tile_27_9_to_tile_26_9_0),
		.out_wire_3_1(vertical_tile_27_9_to_tile_26_9_1),
		.out_wire_3_2(vertical_tile_27_9_to_tile_26_9_2),
		.out_wire_3_3(vertical_tile_27_9_to_tile_26_9_3),
		.in_wire_3_0(vertical_tile_26_9_to_tile_27_9_0),
		.in_wire_3_1(vertical_tile_26_9_to_tile_27_9_1),
		.in_wire_3_2(vertical_tile_26_9_to_tile_27_9_2),
		.in_wire_3_3(vertical_tile_26_9_to_tile_27_9_3),
		.out_wire_1_0(vertical_tile_27_9_to_tile_28_9_0),
		.out_wire_1_1(vertical_tile_27_9_to_tile_28_9_1),
		.out_wire_1_2(vertical_tile_27_9_to_tile_28_9_2),
		.out_wire_1_3(vertical_tile_27_9_to_tile_28_9_3),
		.in_wire_1_0(vertical_tile_28_9_to_tile_27_9_0),
		.in_wire_1_1(vertical_tile_28_9_to_tile_27_9_1),
		.in_wire_1_2(vertical_tile_28_9_to_tile_27_9_2),
		.in_wire_1_3(vertical_tile_28_9_to_tile_27_9_3),
		.out_wire_2_0(horizontal_tile_27_9_to_tile_27_8_0),
		.out_wire_2_1(horizontal_tile_27_9_to_tile_27_8_1),
		.out_wire_2_2(horizontal_tile_27_9_to_tile_27_8_2),
		.out_wire_2_3(horizontal_tile_27_9_to_tile_27_8_3),
		.in_wire_2_0(horizontal_tile_27_8_to_tile_27_9_0),
		.in_wire_2_1(horizontal_tile_27_8_to_tile_27_9_1),
		.in_wire_2_2(horizontal_tile_27_8_to_tile_27_9_2),
		.in_wire_2_3(horizontal_tile_27_8_to_tile_27_9_3),
		.out_wire_0_0(horizontal_tile_27_9_to_tile_27_10_0),
		.out_wire_0_1(horizontal_tile_27_9_to_tile_27_10_1),
		.out_wire_0_2(horizontal_tile_27_9_to_tile_27_10_2),
		.out_wire_0_3(horizontal_tile_27_9_to_tile_27_10_3),
		.in_wire_0_0(horizontal_tile_27_10_to_tile_27_9_0),
		.in_wire_0_1(horizontal_tile_27_10_to_tile_27_9_1),
		.in_wire_0_2(horizontal_tile_27_10_to_tile_27_9_2),
		.in_wire_0_3(horizontal_tile_27_10_to_tile_27_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(874)
	);

	pe_tile pe_tile_27_10(
		.out_wire_3_0(vertical_tile_27_10_to_tile_26_10_0),
		.out_wire_3_1(vertical_tile_27_10_to_tile_26_10_1),
		.out_wire_3_2(vertical_tile_27_10_to_tile_26_10_2),
		.out_wire_3_3(vertical_tile_27_10_to_tile_26_10_3),
		.in_wire_3_0(vertical_tile_26_10_to_tile_27_10_0),
		.in_wire_3_1(vertical_tile_26_10_to_tile_27_10_1),
		.in_wire_3_2(vertical_tile_26_10_to_tile_27_10_2),
		.in_wire_3_3(vertical_tile_26_10_to_tile_27_10_3),
		.out_wire_1_0(vertical_tile_27_10_to_tile_28_10_0),
		.out_wire_1_1(vertical_tile_27_10_to_tile_28_10_1),
		.out_wire_1_2(vertical_tile_27_10_to_tile_28_10_2),
		.out_wire_1_3(vertical_tile_27_10_to_tile_28_10_3),
		.in_wire_1_0(vertical_tile_28_10_to_tile_27_10_0),
		.in_wire_1_1(vertical_tile_28_10_to_tile_27_10_1),
		.in_wire_1_2(vertical_tile_28_10_to_tile_27_10_2),
		.in_wire_1_3(vertical_tile_28_10_to_tile_27_10_3),
		.out_wire_2_0(horizontal_tile_27_10_to_tile_27_9_0),
		.out_wire_2_1(horizontal_tile_27_10_to_tile_27_9_1),
		.out_wire_2_2(horizontal_tile_27_10_to_tile_27_9_2),
		.out_wire_2_3(horizontal_tile_27_10_to_tile_27_9_3),
		.in_wire_2_0(horizontal_tile_27_9_to_tile_27_10_0),
		.in_wire_2_1(horizontal_tile_27_9_to_tile_27_10_1),
		.in_wire_2_2(horizontal_tile_27_9_to_tile_27_10_2),
		.in_wire_2_3(horizontal_tile_27_9_to_tile_27_10_3),
		.out_wire_0_0(horizontal_tile_27_10_to_tile_27_11_0),
		.out_wire_0_1(horizontal_tile_27_10_to_tile_27_11_1),
		.out_wire_0_2(horizontal_tile_27_10_to_tile_27_11_2),
		.out_wire_0_3(horizontal_tile_27_10_to_tile_27_11_3),
		.in_wire_0_0(horizontal_tile_27_11_to_tile_27_10_0),
		.in_wire_0_1(horizontal_tile_27_11_to_tile_27_10_1),
		.in_wire_0_2(horizontal_tile_27_11_to_tile_27_10_2),
		.in_wire_0_3(horizontal_tile_27_11_to_tile_27_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(875)
	);

	pe_tile pe_tile_27_11(
		.out_wire_3_0(vertical_tile_27_11_to_tile_26_11_0),
		.out_wire_3_1(vertical_tile_27_11_to_tile_26_11_1),
		.out_wire_3_2(vertical_tile_27_11_to_tile_26_11_2),
		.out_wire_3_3(vertical_tile_27_11_to_tile_26_11_3),
		.in_wire_3_0(vertical_tile_26_11_to_tile_27_11_0),
		.in_wire_3_1(vertical_tile_26_11_to_tile_27_11_1),
		.in_wire_3_2(vertical_tile_26_11_to_tile_27_11_2),
		.in_wire_3_3(vertical_tile_26_11_to_tile_27_11_3),
		.out_wire_1_0(vertical_tile_27_11_to_tile_28_11_0),
		.out_wire_1_1(vertical_tile_27_11_to_tile_28_11_1),
		.out_wire_1_2(vertical_tile_27_11_to_tile_28_11_2),
		.out_wire_1_3(vertical_tile_27_11_to_tile_28_11_3),
		.in_wire_1_0(vertical_tile_28_11_to_tile_27_11_0),
		.in_wire_1_1(vertical_tile_28_11_to_tile_27_11_1),
		.in_wire_1_2(vertical_tile_28_11_to_tile_27_11_2),
		.in_wire_1_3(vertical_tile_28_11_to_tile_27_11_3),
		.out_wire_2_0(horizontal_tile_27_11_to_tile_27_10_0),
		.out_wire_2_1(horizontal_tile_27_11_to_tile_27_10_1),
		.out_wire_2_2(horizontal_tile_27_11_to_tile_27_10_2),
		.out_wire_2_3(horizontal_tile_27_11_to_tile_27_10_3),
		.in_wire_2_0(horizontal_tile_27_10_to_tile_27_11_0),
		.in_wire_2_1(horizontal_tile_27_10_to_tile_27_11_1),
		.in_wire_2_2(horizontal_tile_27_10_to_tile_27_11_2),
		.in_wire_2_3(horizontal_tile_27_10_to_tile_27_11_3),
		.out_wire_0_0(horizontal_tile_27_11_to_tile_27_12_0),
		.out_wire_0_1(horizontal_tile_27_11_to_tile_27_12_1),
		.out_wire_0_2(horizontal_tile_27_11_to_tile_27_12_2),
		.out_wire_0_3(horizontal_tile_27_11_to_tile_27_12_3),
		.in_wire_0_0(horizontal_tile_27_12_to_tile_27_11_0),
		.in_wire_0_1(horizontal_tile_27_12_to_tile_27_11_1),
		.in_wire_0_2(horizontal_tile_27_12_to_tile_27_11_2),
		.in_wire_0_3(horizontal_tile_27_12_to_tile_27_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(876)
	);

	pe_tile pe_tile_27_12(
		.out_wire_3_0(vertical_tile_27_12_to_tile_26_12_0),
		.out_wire_3_1(vertical_tile_27_12_to_tile_26_12_1),
		.out_wire_3_2(vertical_tile_27_12_to_tile_26_12_2),
		.out_wire_3_3(vertical_tile_27_12_to_tile_26_12_3),
		.in_wire_3_0(vertical_tile_26_12_to_tile_27_12_0),
		.in_wire_3_1(vertical_tile_26_12_to_tile_27_12_1),
		.in_wire_3_2(vertical_tile_26_12_to_tile_27_12_2),
		.in_wire_3_3(vertical_tile_26_12_to_tile_27_12_3),
		.out_wire_1_0(vertical_tile_27_12_to_tile_28_12_0),
		.out_wire_1_1(vertical_tile_27_12_to_tile_28_12_1),
		.out_wire_1_2(vertical_tile_27_12_to_tile_28_12_2),
		.out_wire_1_3(vertical_tile_27_12_to_tile_28_12_3),
		.in_wire_1_0(vertical_tile_28_12_to_tile_27_12_0),
		.in_wire_1_1(vertical_tile_28_12_to_tile_27_12_1),
		.in_wire_1_2(vertical_tile_28_12_to_tile_27_12_2),
		.in_wire_1_3(vertical_tile_28_12_to_tile_27_12_3),
		.out_wire_2_0(horizontal_tile_27_12_to_tile_27_11_0),
		.out_wire_2_1(horizontal_tile_27_12_to_tile_27_11_1),
		.out_wire_2_2(horizontal_tile_27_12_to_tile_27_11_2),
		.out_wire_2_3(horizontal_tile_27_12_to_tile_27_11_3),
		.in_wire_2_0(horizontal_tile_27_11_to_tile_27_12_0),
		.in_wire_2_1(horizontal_tile_27_11_to_tile_27_12_1),
		.in_wire_2_2(horizontal_tile_27_11_to_tile_27_12_2),
		.in_wire_2_3(horizontal_tile_27_11_to_tile_27_12_3),
		.out_wire_0_0(horizontal_tile_27_12_to_tile_27_13_0),
		.out_wire_0_1(horizontal_tile_27_12_to_tile_27_13_1),
		.out_wire_0_2(horizontal_tile_27_12_to_tile_27_13_2),
		.out_wire_0_3(horizontal_tile_27_12_to_tile_27_13_3),
		.in_wire_0_0(horizontal_tile_27_13_to_tile_27_12_0),
		.in_wire_0_1(horizontal_tile_27_13_to_tile_27_12_1),
		.in_wire_0_2(horizontal_tile_27_13_to_tile_27_12_2),
		.in_wire_0_3(horizontal_tile_27_13_to_tile_27_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(877)
	);

	pe_tile pe_tile_27_13(
		.out_wire_3_0(vertical_tile_27_13_to_tile_26_13_0),
		.out_wire_3_1(vertical_tile_27_13_to_tile_26_13_1),
		.out_wire_3_2(vertical_tile_27_13_to_tile_26_13_2),
		.out_wire_3_3(vertical_tile_27_13_to_tile_26_13_3),
		.in_wire_3_0(vertical_tile_26_13_to_tile_27_13_0),
		.in_wire_3_1(vertical_tile_26_13_to_tile_27_13_1),
		.in_wire_3_2(vertical_tile_26_13_to_tile_27_13_2),
		.in_wire_3_3(vertical_tile_26_13_to_tile_27_13_3),
		.out_wire_1_0(vertical_tile_27_13_to_tile_28_13_0),
		.out_wire_1_1(vertical_tile_27_13_to_tile_28_13_1),
		.out_wire_1_2(vertical_tile_27_13_to_tile_28_13_2),
		.out_wire_1_3(vertical_tile_27_13_to_tile_28_13_3),
		.in_wire_1_0(vertical_tile_28_13_to_tile_27_13_0),
		.in_wire_1_1(vertical_tile_28_13_to_tile_27_13_1),
		.in_wire_1_2(vertical_tile_28_13_to_tile_27_13_2),
		.in_wire_1_3(vertical_tile_28_13_to_tile_27_13_3),
		.out_wire_2_0(horizontal_tile_27_13_to_tile_27_12_0),
		.out_wire_2_1(horizontal_tile_27_13_to_tile_27_12_1),
		.out_wire_2_2(horizontal_tile_27_13_to_tile_27_12_2),
		.out_wire_2_3(horizontal_tile_27_13_to_tile_27_12_3),
		.in_wire_2_0(horizontal_tile_27_12_to_tile_27_13_0),
		.in_wire_2_1(horizontal_tile_27_12_to_tile_27_13_1),
		.in_wire_2_2(horizontal_tile_27_12_to_tile_27_13_2),
		.in_wire_2_3(horizontal_tile_27_12_to_tile_27_13_3),
		.out_wire_0_0(horizontal_tile_27_13_to_tile_27_14_0),
		.out_wire_0_1(horizontal_tile_27_13_to_tile_27_14_1),
		.out_wire_0_2(horizontal_tile_27_13_to_tile_27_14_2),
		.out_wire_0_3(horizontal_tile_27_13_to_tile_27_14_3),
		.in_wire_0_0(horizontal_tile_27_14_to_tile_27_13_0),
		.in_wire_0_1(horizontal_tile_27_14_to_tile_27_13_1),
		.in_wire_0_2(horizontal_tile_27_14_to_tile_27_13_2),
		.in_wire_0_3(horizontal_tile_27_14_to_tile_27_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(878)
	);

	pe_tile pe_tile_27_14(
		.out_wire_3_0(vertical_tile_27_14_to_tile_26_14_0),
		.out_wire_3_1(vertical_tile_27_14_to_tile_26_14_1),
		.out_wire_3_2(vertical_tile_27_14_to_tile_26_14_2),
		.out_wire_3_3(vertical_tile_27_14_to_tile_26_14_3),
		.in_wire_3_0(vertical_tile_26_14_to_tile_27_14_0),
		.in_wire_3_1(vertical_tile_26_14_to_tile_27_14_1),
		.in_wire_3_2(vertical_tile_26_14_to_tile_27_14_2),
		.in_wire_3_3(vertical_tile_26_14_to_tile_27_14_3),
		.out_wire_1_0(vertical_tile_27_14_to_tile_28_14_0),
		.out_wire_1_1(vertical_tile_27_14_to_tile_28_14_1),
		.out_wire_1_2(vertical_tile_27_14_to_tile_28_14_2),
		.out_wire_1_3(vertical_tile_27_14_to_tile_28_14_3),
		.in_wire_1_0(vertical_tile_28_14_to_tile_27_14_0),
		.in_wire_1_1(vertical_tile_28_14_to_tile_27_14_1),
		.in_wire_1_2(vertical_tile_28_14_to_tile_27_14_2),
		.in_wire_1_3(vertical_tile_28_14_to_tile_27_14_3),
		.out_wire_2_0(horizontal_tile_27_14_to_tile_27_13_0),
		.out_wire_2_1(horizontal_tile_27_14_to_tile_27_13_1),
		.out_wire_2_2(horizontal_tile_27_14_to_tile_27_13_2),
		.out_wire_2_3(horizontal_tile_27_14_to_tile_27_13_3),
		.in_wire_2_0(horizontal_tile_27_13_to_tile_27_14_0),
		.in_wire_2_1(horizontal_tile_27_13_to_tile_27_14_1),
		.in_wire_2_2(horizontal_tile_27_13_to_tile_27_14_2),
		.in_wire_2_3(horizontal_tile_27_13_to_tile_27_14_3),
		.out_wire_0_0(horizontal_tile_27_14_to_tile_27_15_0),
		.out_wire_0_1(horizontal_tile_27_14_to_tile_27_15_1),
		.out_wire_0_2(horizontal_tile_27_14_to_tile_27_15_2),
		.out_wire_0_3(horizontal_tile_27_14_to_tile_27_15_3),
		.in_wire_0_0(horizontal_tile_27_15_to_tile_27_14_0),
		.in_wire_0_1(horizontal_tile_27_15_to_tile_27_14_1),
		.in_wire_0_2(horizontal_tile_27_15_to_tile_27_14_2),
		.in_wire_0_3(horizontal_tile_27_15_to_tile_27_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(879)
	);

	pe_tile pe_tile_27_15(
		.out_wire_3_0(vertical_tile_27_15_to_tile_26_15_0),
		.out_wire_3_1(vertical_tile_27_15_to_tile_26_15_1),
		.out_wire_3_2(vertical_tile_27_15_to_tile_26_15_2),
		.out_wire_3_3(vertical_tile_27_15_to_tile_26_15_3),
		.in_wire_3_0(vertical_tile_26_15_to_tile_27_15_0),
		.in_wire_3_1(vertical_tile_26_15_to_tile_27_15_1),
		.in_wire_3_2(vertical_tile_26_15_to_tile_27_15_2),
		.in_wire_3_3(vertical_tile_26_15_to_tile_27_15_3),
		.out_wire_1_0(vertical_tile_27_15_to_tile_28_15_0),
		.out_wire_1_1(vertical_tile_27_15_to_tile_28_15_1),
		.out_wire_1_2(vertical_tile_27_15_to_tile_28_15_2),
		.out_wire_1_3(vertical_tile_27_15_to_tile_28_15_3),
		.in_wire_1_0(vertical_tile_28_15_to_tile_27_15_0),
		.in_wire_1_1(vertical_tile_28_15_to_tile_27_15_1),
		.in_wire_1_2(vertical_tile_28_15_to_tile_27_15_2),
		.in_wire_1_3(vertical_tile_28_15_to_tile_27_15_3),
		.out_wire_2_0(horizontal_tile_27_15_to_tile_27_14_0),
		.out_wire_2_1(horizontal_tile_27_15_to_tile_27_14_1),
		.out_wire_2_2(horizontal_tile_27_15_to_tile_27_14_2),
		.out_wire_2_3(horizontal_tile_27_15_to_tile_27_14_3),
		.in_wire_2_0(horizontal_tile_27_14_to_tile_27_15_0),
		.in_wire_2_1(horizontal_tile_27_14_to_tile_27_15_1),
		.in_wire_2_2(horizontal_tile_27_14_to_tile_27_15_2),
		.in_wire_2_3(horizontal_tile_27_14_to_tile_27_15_3),
		.out_wire_0_0(horizontal_tile_27_15_to_tile_27_16_0),
		.out_wire_0_1(horizontal_tile_27_15_to_tile_27_16_1),
		.out_wire_0_2(horizontal_tile_27_15_to_tile_27_16_2),
		.out_wire_0_3(horizontal_tile_27_15_to_tile_27_16_3),
		.in_wire_0_0(horizontal_tile_27_16_to_tile_27_15_0),
		.in_wire_0_1(horizontal_tile_27_16_to_tile_27_15_1),
		.in_wire_0_2(horizontal_tile_27_16_to_tile_27_15_2),
		.in_wire_0_3(horizontal_tile_27_16_to_tile_27_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(880)
	);

	pe_tile pe_tile_27_16(
		.out_wire_3_0(vertical_tile_27_16_to_tile_26_16_0),
		.out_wire_3_1(vertical_tile_27_16_to_tile_26_16_1),
		.out_wire_3_2(vertical_tile_27_16_to_tile_26_16_2),
		.out_wire_3_3(vertical_tile_27_16_to_tile_26_16_3),
		.in_wire_3_0(vertical_tile_26_16_to_tile_27_16_0),
		.in_wire_3_1(vertical_tile_26_16_to_tile_27_16_1),
		.in_wire_3_2(vertical_tile_26_16_to_tile_27_16_2),
		.in_wire_3_3(vertical_tile_26_16_to_tile_27_16_3),
		.out_wire_1_0(vertical_tile_27_16_to_tile_28_16_0),
		.out_wire_1_1(vertical_tile_27_16_to_tile_28_16_1),
		.out_wire_1_2(vertical_tile_27_16_to_tile_28_16_2),
		.out_wire_1_3(vertical_tile_27_16_to_tile_28_16_3),
		.in_wire_1_0(vertical_tile_28_16_to_tile_27_16_0),
		.in_wire_1_1(vertical_tile_28_16_to_tile_27_16_1),
		.in_wire_1_2(vertical_tile_28_16_to_tile_27_16_2),
		.in_wire_1_3(vertical_tile_28_16_to_tile_27_16_3),
		.out_wire_2_0(horizontal_tile_27_16_to_tile_27_15_0),
		.out_wire_2_1(horizontal_tile_27_16_to_tile_27_15_1),
		.out_wire_2_2(horizontal_tile_27_16_to_tile_27_15_2),
		.out_wire_2_3(horizontal_tile_27_16_to_tile_27_15_3),
		.in_wire_2_0(horizontal_tile_27_15_to_tile_27_16_0),
		.in_wire_2_1(horizontal_tile_27_15_to_tile_27_16_1),
		.in_wire_2_2(horizontal_tile_27_15_to_tile_27_16_2),
		.in_wire_2_3(horizontal_tile_27_15_to_tile_27_16_3),
		.out_wire_0_0(horizontal_tile_27_16_to_tile_27_17_0),
		.out_wire_0_1(horizontal_tile_27_16_to_tile_27_17_1),
		.out_wire_0_2(horizontal_tile_27_16_to_tile_27_17_2),
		.out_wire_0_3(horizontal_tile_27_16_to_tile_27_17_3),
		.in_wire_0_0(horizontal_tile_27_17_to_tile_27_16_0),
		.in_wire_0_1(horizontal_tile_27_17_to_tile_27_16_1),
		.in_wire_0_2(horizontal_tile_27_17_to_tile_27_16_2),
		.in_wire_0_3(horizontal_tile_27_17_to_tile_27_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(881)
	);

	pe_tile pe_tile_27_17(
		.out_wire_3_0(vertical_tile_27_17_to_tile_26_17_0),
		.out_wire_3_1(vertical_tile_27_17_to_tile_26_17_1),
		.out_wire_3_2(vertical_tile_27_17_to_tile_26_17_2),
		.out_wire_3_3(vertical_tile_27_17_to_tile_26_17_3),
		.in_wire_3_0(vertical_tile_26_17_to_tile_27_17_0),
		.in_wire_3_1(vertical_tile_26_17_to_tile_27_17_1),
		.in_wire_3_2(vertical_tile_26_17_to_tile_27_17_2),
		.in_wire_3_3(vertical_tile_26_17_to_tile_27_17_3),
		.out_wire_1_0(vertical_tile_27_17_to_tile_28_17_0),
		.out_wire_1_1(vertical_tile_27_17_to_tile_28_17_1),
		.out_wire_1_2(vertical_tile_27_17_to_tile_28_17_2),
		.out_wire_1_3(vertical_tile_27_17_to_tile_28_17_3),
		.in_wire_1_0(vertical_tile_28_17_to_tile_27_17_0),
		.in_wire_1_1(vertical_tile_28_17_to_tile_27_17_1),
		.in_wire_1_2(vertical_tile_28_17_to_tile_27_17_2),
		.in_wire_1_3(vertical_tile_28_17_to_tile_27_17_3),
		.out_wire_2_0(horizontal_tile_27_17_to_tile_27_16_0),
		.out_wire_2_1(horizontal_tile_27_17_to_tile_27_16_1),
		.out_wire_2_2(horizontal_tile_27_17_to_tile_27_16_2),
		.out_wire_2_3(horizontal_tile_27_17_to_tile_27_16_3),
		.in_wire_2_0(horizontal_tile_27_16_to_tile_27_17_0),
		.in_wire_2_1(horizontal_tile_27_16_to_tile_27_17_1),
		.in_wire_2_2(horizontal_tile_27_16_to_tile_27_17_2),
		.in_wire_2_3(horizontal_tile_27_16_to_tile_27_17_3),
		.out_wire_0_0(horizontal_tile_27_17_to_tile_27_18_0),
		.out_wire_0_1(horizontal_tile_27_17_to_tile_27_18_1),
		.out_wire_0_2(horizontal_tile_27_17_to_tile_27_18_2),
		.out_wire_0_3(horizontal_tile_27_17_to_tile_27_18_3),
		.in_wire_0_0(horizontal_tile_27_18_to_tile_27_17_0),
		.in_wire_0_1(horizontal_tile_27_18_to_tile_27_17_1),
		.in_wire_0_2(horizontal_tile_27_18_to_tile_27_17_2),
		.in_wire_0_3(horizontal_tile_27_18_to_tile_27_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(882)
	);

	pe_tile pe_tile_27_18(
		.out_wire_3_0(vertical_tile_27_18_to_tile_26_18_0),
		.out_wire_3_1(vertical_tile_27_18_to_tile_26_18_1),
		.out_wire_3_2(vertical_tile_27_18_to_tile_26_18_2),
		.out_wire_3_3(vertical_tile_27_18_to_tile_26_18_3),
		.in_wire_3_0(vertical_tile_26_18_to_tile_27_18_0),
		.in_wire_3_1(vertical_tile_26_18_to_tile_27_18_1),
		.in_wire_3_2(vertical_tile_26_18_to_tile_27_18_2),
		.in_wire_3_3(vertical_tile_26_18_to_tile_27_18_3),
		.out_wire_1_0(vertical_tile_27_18_to_tile_28_18_0),
		.out_wire_1_1(vertical_tile_27_18_to_tile_28_18_1),
		.out_wire_1_2(vertical_tile_27_18_to_tile_28_18_2),
		.out_wire_1_3(vertical_tile_27_18_to_tile_28_18_3),
		.in_wire_1_0(vertical_tile_28_18_to_tile_27_18_0),
		.in_wire_1_1(vertical_tile_28_18_to_tile_27_18_1),
		.in_wire_1_2(vertical_tile_28_18_to_tile_27_18_2),
		.in_wire_1_3(vertical_tile_28_18_to_tile_27_18_3),
		.out_wire_2_0(horizontal_tile_27_18_to_tile_27_17_0),
		.out_wire_2_1(horizontal_tile_27_18_to_tile_27_17_1),
		.out_wire_2_2(horizontal_tile_27_18_to_tile_27_17_2),
		.out_wire_2_3(horizontal_tile_27_18_to_tile_27_17_3),
		.in_wire_2_0(horizontal_tile_27_17_to_tile_27_18_0),
		.in_wire_2_1(horizontal_tile_27_17_to_tile_27_18_1),
		.in_wire_2_2(horizontal_tile_27_17_to_tile_27_18_2),
		.in_wire_2_3(horizontal_tile_27_17_to_tile_27_18_3),
		.out_wire_0_0(horizontal_tile_27_18_to_tile_27_19_0),
		.out_wire_0_1(horizontal_tile_27_18_to_tile_27_19_1),
		.out_wire_0_2(horizontal_tile_27_18_to_tile_27_19_2),
		.out_wire_0_3(horizontal_tile_27_18_to_tile_27_19_3),
		.in_wire_0_0(horizontal_tile_27_19_to_tile_27_18_0),
		.in_wire_0_1(horizontal_tile_27_19_to_tile_27_18_1),
		.in_wire_0_2(horizontal_tile_27_19_to_tile_27_18_2),
		.in_wire_0_3(horizontal_tile_27_19_to_tile_27_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(883)
	);

	pe_tile pe_tile_27_19(
		.out_wire_3_0(vertical_tile_27_19_to_tile_26_19_0),
		.out_wire_3_1(vertical_tile_27_19_to_tile_26_19_1),
		.out_wire_3_2(vertical_tile_27_19_to_tile_26_19_2),
		.out_wire_3_3(vertical_tile_27_19_to_tile_26_19_3),
		.in_wire_3_0(vertical_tile_26_19_to_tile_27_19_0),
		.in_wire_3_1(vertical_tile_26_19_to_tile_27_19_1),
		.in_wire_3_2(vertical_tile_26_19_to_tile_27_19_2),
		.in_wire_3_3(vertical_tile_26_19_to_tile_27_19_3),
		.out_wire_1_0(vertical_tile_27_19_to_tile_28_19_0),
		.out_wire_1_1(vertical_tile_27_19_to_tile_28_19_1),
		.out_wire_1_2(vertical_tile_27_19_to_tile_28_19_2),
		.out_wire_1_3(vertical_tile_27_19_to_tile_28_19_3),
		.in_wire_1_0(vertical_tile_28_19_to_tile_27_19_0),
		.in_wire_1_1(vertical_tile_28_19_to_tile_27_19_1),
		.in_wire_1_2(vertical_tile_28_19_to_tile_27_19_2),
		.in_wire_1_3(vertical_tile_28_19_to_tile_27_19_3),
		.out_wire_2_0(horizontal_tile_27_19_to_tile_27_18_0),
		.out_wire_2_1(horizontal_tile_27_19_to_tile_27_18_1),
		.out_wire_2_2(horizontal_tile_27_19_to_tile_27_18_2),
		.out_wire_2_3(horizontal_tile_27_19_to_tile_27_18_3),
		.in_wire_2_0(horizontal_tile_27_18_to_tile_27_19_0),
		.in_wire_2_1(horizontal_tile_27_18_to_tile_27_19_1),
		.in_wire_2_2(horizontal_tile_27_18_to_tile_27_19_2),
		.in_wire_2_3(horizontal_tile_27_18_to_tile_27_19_3),
		.out_wire_0_0(horizontal_tile_27_19_to_tile_27_20_0),
		.out_wire_0_1(horizontal_tile_27_19_to_tile_27_20_1),
		.out_wire_0_2(horizontal_tile_27_19_to_tile_27_20_2),
		.out_wire_0_3(horizontal_tile_27_19_to_tile_27_20_3),
		.in_wire_0_0(horizontal_tile_27_20_to_tile_27_19_0),
		.in_wire_0_1(horizontal_tile_27_20_to_tile_27_19_1),
		.in_wire_0_2(horizontal_tile_27_20_to_tile_27_19_2),
		.in_wire_0_3(horizontal_tile_27_20_to_tile_27_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(884)
	);

	pe_tile pe_tile_27_20(
		.out_wire_3_0(vertical_tile_27_20_to_tile_26_20_0),
		.out_wire_3_1(vertical_tile_27_20_to_tile_26_20_1),
		.out_wire_3_2(vertical_tile_27_20_to_tile_26_20_2),
		.out_wire_3_3(vertical_tile_27_20_to_tile_26_20_3),
		.in_wire_3_0(vertical_tile_26_20_to_tile_27_20_0),
		.in_wire_3_1(vertical_tile_26_20_to_tile_27_20_1),
		.in_wire_3_2(vertical_tile_26_20_to_tile_27_20_2),
		.in_wire_3_3(vertical_tile_26_20_to_tile_27_20_3),
		.out_wire_1_0(vertical_tile_27_20_to_tile_28_20_0),
		.out_wire_1_1(vertical_tile_27_20_to_tile_28_20_1),
		.out_wire_1_2(vertical_tile_27_20_to_tile_28_20_2),
		.out_wire_1_3(vertical_tile_27_20_to_tile_28_20_3),
		.in_wire_1_0(vertical_tile_28_20_to_tile_27_20_0),
		.in_wire_1_1(vertical_tile_28_20_to_tile_27_20_1),
		.in_wire_1_2(vertical_tile_28_20_to_tile_27_20_2),
		.in_wire_1_3(vertical_tile_28_20_to_tile_27_20_3),
		.out_wire_2_0(horizontal_tile_27_20_to_tile_27_19_0),
		.out_wire_2_1(horizontal_tile_27_20_to_tile_27_19_1),
		.out_wire_2_2(horizontal_tile_27_20_to_tile_27_19_2),
		.out_wire_2_3(horizontal_tile_27_20_to_tile_27_19_3),
		.in_wire_2_0(horizontal_tile_27_19_to_tile_27_20_0),
		.in_wire_2_1(horizontal_tile_27_19_to_tile_27_20_1),
		.in_wire_2_2(horizontal_tile_27_19_to_tile_27_20_2),
		.in_wire_2_3(horizontal_tile_27_19_to_tile_27_20_3),
		.out_wire_0_0(horizontal_tile_27_20_to_tile_27_21_0),
		.out_wire_0_1(horizontal_tile_27_20_to_tile_27_21_1),
		.out_wire_0_2(horizontal_tile_27_20_to_tile_27_21_2),
		.out_wire_0_3(horizontal_tile_27_20_to_tile_27_21_3),
		.in_wire_0_0(horizontal_tile_27_21_to_tile_27_20_0),
		.in_wire_0_1(horizontal_tile_27_21_to_tile_27_20_1),
		.in_wire_0_2(horizontal_tile_27_21_to_tile_27_20_2),
		.in_wire_0_3(horizontal_tile_27_21_to_tile_27_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(885)
	);

	pe_tile pe_tile_27_21(
		.out_wire_3_0(vertical_tile_27_21_to_tile_26_21_0),
		.out_wire_3_1(vertical_tile_27_21_to_tile_26_21_1),
		.out_wire_3_2(vertical_tile_27_21_to_tile_26_21_2),
		.out_wire_3_3(vertical_tile_27_21_to_tile_26_21_3),
		.in_wire_3_0(vertical_tile_26_21_to_tile_27_21_0),
		.in_wire_3_1(vertical_tile_26_21_to_tile_27_21_1),
		.in_wire_3_2(vertical_tile_26_21_to_tile_27_21_2),
		.in_wire_3_3(vertical_tile_26_21_to_tile_27_21_3),
		.out_wire_1_0(vertical_tile_27_21_to_tile_28_21_0),
		.out_wire_1_1(vertical_tile_27_21_to_tile_28_21_1),
		.out_wire_1_2(vertical_tile_27_21_to_tile_28_21_2),
		.out_wire_1_3(vertical_tile_27_21_to_tile_28_21_3),
		.in_wire_1_0(vertical_tile_28_21_to_tile_27_21_0),
		.in_wire_1_1(vertical_tile_28_21_to_tile_27_21_1),
		.in_wire_1_2(vertical_tile_28_21_to_tile_27_21_2),
		.in_wire_1_3(vertical_tile_28_21_to_tile_27_21_3),
		.out_wire_2_0(horizontal_tile_27_21_to_tile_27_20_0),
		.out_wire_2_1(horizontal_tile_27_21_to_tile_27_20_1),
		.out_wire_2_2(horizontal_tile_27_21_to_tile_27_20_2),
		.out_wire_2_3(horizontal_tile_27_21_to_tile_27_20_3),
		.in_wire_2_0(horizontal_tile_27_20_to_tile_27_21_0),
		.in_wire_2_1(horizontal_tile_27_20_to_tile_27_21_1),
		.in_wire_2_2(horizontal_tile_27_20_to_tile_27_21_2),
		.in_wire_2_3(horizontal_tile_27_20_to_tile_27_21_3),
		.out_wire_0_0(horizontal_tile_27_21_to_tile_27_22_0),
		.out_wire_0_1(horizontal_tile_27_21_to_tile_27_22_1),
		.out_wire_0_2(horizontal_tile_27_21_to_tile_27_22_2),
		.out_wire_0_3(horizontal_tile_27_21_to_tile_27_22_3),
		.in_wire_0_0(horizontal_tile_27_22_to_tile_27_21_0),
		.in_wire_0_1(horizontal_tile_27_22_to_tile_27_21_1),
		.in_wire_0_2(horizontal_tile_27_22_to_tile_27_21_2),
		.in_wire_0_3(horizontal_tile_27_22_to_tile_27_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(886)
	);

	pe_tile pe_tile_27_22(
		.out_wire_3_0(vertical_tile_27_22_to_tile_26_22_0),
		.out_wire_3_1(vertical_tile_27_22_to_tile_26_22_1),
		.out_wire_3_2(vertical_tile_27_22_to_tile_26_22_2),
		.out_wire_3_3(vertical_tile_27_22_to_tile_26_22_3),
		.in_wire_3_0(vertical_tile_26_22_to_tile_27_22_0),
		.in_wire_3_1(vertical_tile_26_22_to_tile_27_22_1),
		.in_wire_3_2(vertical_tile_26_22_to_tile_27_22_2),
		.in_wire_3_3(vertical_tile_26_22_to_tile_27_22_3),
		.out_wire_1_0(vertical_tile_27_22_to_tile_28_22_0),
		.out_wire_1_1(vertical_tile_27_22_to_tile_28_22_1),
		.out_wire_1_2(vertical_tile_27_22_to_tile_28_22_2),
		.out_wire_1_3(vertical_tile_27_22_to_tile_28_22_3),
		.in_wire_1_0(vertical_tile_28_22_to_tile_27_22_0),
		.in_wire_1_1(vertical_tile_28_22_to_tile_27_22_1),
		.in_wire_1_2(vertical_tile_28_22_to_tile_27_22_2),
		.in_wire_1_3(vertical_tile_28_22_to_tile_27_22_3),
		.out_wire_2_0(horizontal_tile_27_22_to_tile_27_21_0),
		.out_wire_2_1(horizontal_tile_27_22_to_tile_27_21_1),
		.out_wire_2_2(horizontal_tile_27_22_to_tile_27_21_2),
		.out_wire_2_3(horizontal_tile_27_22_to_tile_27_21_3),
		.in_wire_2_0(horizontal_tile_27_21_to_tile_27_22_0),
		.in_wire_2_1(horizontal_tile_27_21_to_tile_27_22_1),
		.in_wire_2_2(horizontal_tile_27_21_to_tile_27_22_2),
		.in_wire_2_3(horizontal_tile_27_21_to_tile_27_22_3),
		.out_wire_0_0(horizontal_tile_27_22_to_tile_27_23_0),
		.out_wire_0_1(horizontal_tile_27_22_to_tile_27_23_1),
		.out_wire_0_2(horizontal_tile_27_22_to_tile_27_23_2),
		.out_wire_0_3(horizontal_tile_27_22_to_tile_27_23_3),
		.in_wire_0_0(horizontal_tile_27_23_to_tile_27_22_0),
		.in_wire_0_1(horizontal_tile_27_23_to_tile_27_22_1),
		.in_wire_0_2(horizontal_tile_27_23_to_tile_27_22_2),
		.in_wire_0_3(horizontal_tile_27_23_to_tile_27_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(887)
	);

	pe_tile pe_tile_27_23(
		.out_wire_3_0(vertical_tile_27_23_to_tile_26_23_0),
		.out_wire_3_1(vertical_tile_27_23_to_tile_26_23_1),
		.out_wire_3_2(vertical_tile_27_23_to_tile_26_23_2),
		.out_wire_3_3(vertical_tile_27_23_to_tile_26_23_3),
		.in_wire_3_0(vertical_tile_26_23_to_tile_27_23_0),
		.in_wire_3_1(vertical_tile_26_23_to_tile_27_23_1),
		.in_wire_3_2(vertical_tile_26_23_to_tile_27_23_2),
		.in_wire_3_3(vertical_tile_26_23_to_tile_27_23_3),
		.out_wire_1_0(vertical_tile_27_23_to_tile_28_23_0),
		.out_wire_1_1(vertical_tile_27_23_to_tile_28_23_1),
		.out_wire_1_2(vertical_tile_27_23_to_tile_28_23_2),
		.out_wire_1_3(vertical_tile_27_23_to_tile_28_23_3),
		.in_wire_1_0(vertical_tile_28_23_to_tile_27_23_0),
		.in_wire_1_1(vertical_tile_28_23_to_tile_27_23_1),
		.in_wire_1_2(vertical_tile_28_23_to_tile_27_23_2),
		.in_wire_1_3(vertical_tile_28_23_to_tile_27_23_3),
		.out_wire_2_0(horizontal_tile_27_23_to_tile_27_22_0),
		.out_wire_2_1(horizontal_tile_27_23_to_tile_27_22_1),
		.out_wire_2_2(horizontal_tile_27_23_to_tile_27_22_2),
		.out_wire_2_3(horizontal_tile_27_23_to_tile_27_22_3),
		.in_wire_2_0(horizontal_tile_27_22_to_tile_27_23_0),
		.in_wire_2_1(horizontal_tile_27_22_to_tile_27_23_1),
		.in_wire_2_2(horizontal_tile_27_22_to_tile_27_23_2),
		.in_wire_2_3(horizontal_tile_27_22_to_tile_27_23_3),
		.out_wire_0_0(horizontal_tile_27_23_to_tile_27_24_0),
		.out_wire_0_1(horizontal_tile_27_23_to_tile_27_24_1),
		.out_wire_0_2(horizontal_tile_27_23_to_tile_27_24_2),
		.out_wire_0_3(horizontal_tile_27_23_to_tile_27_24_3),
		.in_wire_0_0(horizontal_tile_27_24_to_tile_27_23_0),
		.in_wire_0_1(horizontal_tile_27_24_to_tile_27_23_1),
		.in_wire_0_2(horizontal_tile_27_24_to_tile_27_23_2),
		.in_wire_0_3(horizontal_tile_27_24_to_tile_27_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(888)
	);

	pe_tile pe_tile_27_24(
		.out_wire_3_0(vertical_tile_27_24_to_tile_26_24_0),
		.out_wire_3_1(vertical_tile_27_24_to_tile_26_24_1),
		.out_wire_3_2(vertical_tile_27_24_to_tile_26_24_2),
		.out_wire_3_3(vertical_tile_27_24_to_tile_26_24_3),
		.in_wire_3_0(vertical_tile_26_24_to_tile_27_24_0),
		.in_wire_3_1(vertical_tile_26_24_to_tile_27_24_1),
		.in_wire_3_2(vertical_tile_26_24_to_tile_27_24_2),
		.in_wire_3_3(vertical_tile_26_24_to_tile_27_24_3),
		.out_wire_1_0(vertical_tile_27_24_to_tile_28_24_0),
		.out_wire_1_1(vertical_tile_27_24_to_tile_28_24_1),
		.out_wire_1_2(vertical_tile_27_24_to_tile_28_24_2),
		.out_wire_1_3(vertical_tile_27_24_to_tile_28_24_3),
		.in_wire_1_0(vertical_tile_28_24_to_tile_27_24_0),
		.in_wire_1_1(vertical_tile_28_24_to_tile_27_24_1),
		.in_wire_1_2(vertical_tile_28_24_to_tile_27_24_2),
		.in_wire_1_3(vertical_tile_28_24_to_tile_27_24_3),
		.out_wire_2_0(horizontal_tile_27_24_to_tile_27_23_0),
		.out_wire_2_1(horizontal_tile_27_24_to_tile_27_23_1),
		.out_wire_2_2(horizontal_tile_27_24_to_tile_27_23_2),
		.out_wire_2_3(horizontal_tile_27_24_to_tile_27_23_3),
		.in_wire_2_0(horizontal_tile_27_23_to_tile_27_24_0),
		.in_wire_2_1(horizontal_tile_27_23_to_tile_27_24_1),
		.in_wire_2_2(horizontal_tile_27_23_to_tile_27_24_2),
		.in_wire_2_3(horizontal_tile_27_23_to_tile_27_24_3),
		.out_wire_0_0(horizontal_tile_27_24_to_tile_27_25_0),
		.out_wire_0_1(horizontal_tile_27_24_to_tile_27_25_1),
		.out_wire_0_2(horizontal_tile_27_24_to_tile_27_25_2),
		.out_wire_0_3(horizontal_tile_27_24_to_tile_27_25_3),
		.in_wire_0_0(horizontal_tile_27_25_to_tile_27_24_0),
		.in_wire_0_1(horizontal_tile_27_25_to_tile_27_24_1),
		.in_wire_0_2(horizontal_tile_27_25_to_tile_27_24_2),
		.in_wire_0_3(horizontal_tile_27_25_to_tile_27_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(889)
	);

	pe_tile pe_tile_27_25(
		.out_wire_3_0(vertical_tile_27_25_to_tile_26_25_0),
		.out_wire_3_1(vertical_tile_27_25_to_tile_26_25_1),
		.out_wire_3_2(vertical_tile_27_25_to_tile_26_25_2),
		.out_wire_3_3(vertical_tile_27_25_to_tile_26_25_3),
		.in_wire_3_0(vertical_tile_26_25_to_tile_27_25_0),
		.in_wire_3_1(vertical_tile_26_25_to_tile_27_25_1),
		.in_wire_3_2(vertical_tile_26_25_to_tile_27_25_2),
		.in_wire_3_3(vertical_tile_26_25_to_tile_27_25_3),
		.out_wire_1_0(vertical_tile_27_25_to_tile_28_25_0),
		.out_wire_1_1(vertical_tile_27_25_to_tile_28_25_1),
		.out_wire_1_2(vertical_tile_27_25_to_tile_28_25_2),
		.out_wire_1_3(vertical_tile_27_25_to_tile_28_25_3),
		.in_wire_1_0(vertical_tile_28_25_to_tile_27_25_0),
		.in_wire_1_1(vertical_tile_28_25_to_tile_27_25_1),
		.in_wire_1_2(vertical_tile_28_25_to_tile_27_25_2),
		.in_wire_1_3(vertical_tile_28_25_to_tile_27_25_3),
		.out_wire_2_0(horizontal_tile_27_25_to_tile_27_24_0),
		.out_wire_2_1(horizontal_tile_27_25_to_tile_27_24_1),
		.out_wire_2_2(horizontal_tile_27_25_to_tile_27_24_2),
		.out_wire_2_3(horizontal_tile_27_25_to_tile_27_24_3),
		.in_wire_2_0(horizontal_tile_27_24_to_tile_27_25_0),
		.in_wire_2_1(horizontal_tile_27_24_to_tile_27_25_1),
		.in_wire_2_2(horizontal_tile_27_24_to_tile_27_25_2),
		.in_wire_2_3(horizontal_tile_27_24_to_tile_27_25_3),
		.out_wire_0_0(horizontal_tile_27_25_to_tile_27_26_0),
		.out_wire_0_1(horizontal_tile_27_25_to_tile_27_26_1),
		.out_wire_0_2(horizontal_tile_27_25_to_tile_27_26_2),
		.out_wire_0_3(horizontal_tile_27_25_to_tile_27_26_3),
		.in_wire_0_0(horizontal_tile_27_26_to_tile_27_25_0),
		.in_wire_0_1(horizontal_tile_27_26_to_tile_27_25_1),
		.in_wire_0_2(horizontal_tile_27_26_to_tile_27_25_2),
		.in_wire_0_3(horizontal_tile_27_26_to_tile_27_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(890)
	);

	pe_tile pe_tile_27_26(
		.out_wire_3_0(vertical_tile_27_26_to_tile_26_26_0),
		.out_wire_3_1(vertical_tile_27_26_to_tile_26_26_1),
		.out_wire_3_2(vertical_tile_27_26_to_tile_26_26_2),
		.out_wire_3_3(vertical_tile_27_26_to_tile_26_26_3),
		.in_wire_3_0(vertical_tile_26_26_to_tile_27_26_0),
		.in_wire_3_1(vertical_tile_26_26_to_tile_27_26_1),
		.in_wire_3_2(vertical_tile_26_26_to_tile_27_26_2),
		.in_wire_3_3(vertical_tile_26_26_to_tile_27_26_3),
		.out_wire_1_0(vertical_tile_27_26_to_tile_28_26_0),
		.out_wire_1_1(vertical_tile_27_26_to_tile_28_26_1),
		.out_wire_1_2(vertical_tile_27_26_to_tile_28_26_2),
		.out_wire_1_3(vertical_tile_27_26_to_tile_28_26_3),
		.in_wire_1_0(vertical_tile_28_26_to_tile_27_26_0),
		.in_wire_1_1(vertical_tile_28_26_to_tile_27_26_1),
		.in_wire_1_2(vertical_tile_28_26_to_tile_27_26_2),
		.in_wire_1_3(vertical_tile_28_26_to_tile_27_26_3),
		.out_wire_2_0(horizontal_tile_27_26_to_tile_27_25_0),
		.out_wire_2_1(horizontal_tile_27_26_to_tile_27_25_1),
		.out_wire_2_2(horizontal_tile_27_26_to_tile_27_25_2),
		.out_wire_2_3(horizontal_tile_27_26_to_tile_27_25_3),
		.in_wire_2_0(horizontal_tile_27_25_to_tile_27_26_0),
		.in_wire_2_1(horizontal_tile_27_25_to_tile_27_26_1),
		.in_wire_2_2(horizontal_tile_27_25_to_tile_27_26_2),
		.in_wire_2_3(horizontal_tile_27_25_to_tile_27_26_3),
		.out_wire_0_0(horizontal_tile_27_26_to_tile_27_27_0),
		.out_wire_0_1(horizontal_tile_27_26_to_tile_27_27_1),
		.out_wire_0_2(horizontal_tile_27_26_to_tile_27_27_2),
		.out_wire_0_3(horizontal_tile_27_26_to_tile_27_27_3),
		.in_wire_0_0(horizontal_tile_27_27_to_tile_27_26_0),
		.in_wire_0_1(horizontal_tile_27_27_to_tile_27_26_1),
		.in_wire_0_2(horizontal_tile_27_27_to_tile_27_26_2),
		.in_wire_0_3(horizontal_tile_27_27_to_tile_27_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(891)
	);

	pe_tile pe_tile_27_27(
		.out_wire_3_0(vertical_tile_27_27_to_tile_26_27_0),
		.out_wire_3_1(vertical_tile_27_27_to_tile_26_27_1),
		.out_wire_3_2(vertical_tile_27_27_to_tile_26_27_2),
		.out_wire_3_3(vertical_tile_27_27_to_tile_26_27_3),
		.in_wire_3_0(vertical_tile_26_27_to_tile_27_27_0),
		.in_wire_3_1(vertical_tile_26_27_to_tile_27_27_1),
		.in_wire_3_2(vertical_tile_26_27_to_tile_27_27_2),
		.in_wire_3_3(vertical_tile_26_27_to_tile_27_27_3),
		.out_wire_1_0(vertical_tile_27_27_to_tile_28_27_0),
		.out_wire_1_1(vertical_tile_27_27_to_tile_28_27_1),
		.out_wire_1_2(vertical_tile_27_27_to_tile_28_27_2),
		.out_wire_1_3(vertical_tile_27_27_to_tile_28_27_3),
		.in_wire_1_0(vertical_tile_28_27_to_tile_27_27_0),
		.in_wire_1_1(vertical_tile_28_27_to_tile_27_27_1),
		.in_wire_1_2(vertical_tile_28_27_to_tile_27_27_2),
		.in_wire_1_3(vertical_tile_28_27_to_tile_27_27_3),
		.out_wire_2_0(horizontal_tile_27_27_to_tile_27_26_0),
		.out_wire_2_1(horizontal_tile_27_27_to_tile_27_26_1),
		.out_wire_2_2(horizontal_tile_27_27_to_tile_27_26_2),
		.out_wire_2_3(horizontal_tile_27_27_to_tile_27_26_3),
		.in_wire_2_0(horizontal_tile_27_26_to_tile_27_27_0),
		.in_wire_2_1(horizontal_tile_27_26_to_tile_27_27_1),
		.in_wire_2_2(horizontal_tile_27_26_to_tile_27_27_2),
		.in_wire_2_3(horizontal_tile_27_26_to_tile_27_27_3),
		.out_wire_0_0(horizontal_tile_27_27_to_tile_27_28_0),
		.out_wire_0_1(horizontal_tile_27_27_to_tile_27_28_1),
		.out_wire_0_2(horizontal_tile_27_27_to_tile_27_28_2),
		.out_wire_0_3(horizontal_tile_27_27_to_tile_27_28_3),
		.in_wire_0_0(horizontal_tile_27_28_to_tile_27_27_0),
		.in_wire_0_1(horizontal_tile_27_28_to_tile_27_27_1),
		.in_wire_0_2(horizontal_tile_27_28_to_tile_27_27_2),
		.in_wire_0_3(horizontal_tile_27_28_to_tile_27_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(892)
	);

	pe_tile pe_tile_27_28(
		.out_wire_3_0(vertical_tile_27_28_to_tile_26_28_0),
		.out_wire_3_1(vertical_tile_27_28_to_tile_26_28_1),
		.out_wire_3_2(vertical_tile_27_28_to_tile_26_28_2),
		.out_wire_3_3(vertical_tile_27_28_to_tile_26_28_3),
		.in_wire_3_0(vertical_tile_26_28_to_tile_27_28_0),
		.in_wire_3_1(vertical_tile_26_28_to_tile_27_28_1),
		.in_wire_3_2(vertical_tile_26_28_to_tile_27_28_2),
		.in_wire_3_3(vertical_tile_26_28_to_tile_27_28_3),
		.out_wire_1_0(vertical_tile_27_28_to_tile_28_28_0),
		.out_wire_1_1(vertical_tile_27_28_to_tile_28_28_1),
		.out_wire_1_2(vertical_tile_27_28_to_tile_28_28_2),
		.out_wire_1_3(vertical_tile_27_28_to_tile_28_28_3),
		.in_wire_1_0(vertical_tile_28_28_to_tile_27_28_0),
		.in_wire_1_1(vertical_tile_28_28_to_tile_27_28_1),
		.in_wire_1_2(vertical_tile_28_28_to_tile_27_28_2),
		.in_wire_1_3(vertical_tile_28_28_to_tile_27_28_3),
		.out_wire_2_0(horizontal_tile_27_28_to_tile_27_27_0),
		.out_wire_2_1(horizontal_tile_27_28_to_tile_27_27_1),
		.out_wire_2_2(horizontal_tile_27_28_to_tile_27_27_2),
		.out_wire_2_3(horizontal_tile_27_28_to_tile_27_27_3),
		.in_wire_2_0(horizontal_tile_27_27_to_tile_27_28_0),
		.in_wire_2_1(horizontal_tile_27_27_to_tile_27_28_1),
		.in_wire_2_2(horizontal_tile_27_27_to_tile_27_28_2),
		.in_wire_2_3(horizontal_tile_27_27_to_tile_27_28_3),
		.out_wire_0_0(horizontal_tile_27_28_to_tile_27_29_0),
		.out_wire_0_1(horizontal_tile_27_28_to_tile_27_29_1),
		.out_wire_0_2(horizontal_tile_27_28_to_tile_27_29_2),
		.out_wire_0_3(horizontal_tile_27_28_to_tile_27_29_3),
		.in_wire_0_0(horizontal_tile_27_29_to_tile_27_28_0),
		.in_wire_0_1(horizontal_tile_27_29_to_tile_27_28_1),
		.in_wire_0_2(horizontal_tile_27_29_to_tile_27_28_2),
		.in_wire_0_3(horizontal_tile_27_29_to_tile_27_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(893)
	);

	pe_tile pe_tile_27_29(
		.out_wire_3_0(vertical_tile_27_29_to_tile_26_29_0),
		.out_wire_3_1(vertical_tile_27_29_to_tile_26_29_1),
		.out_wire_3_2(vertical_tile_27_29_to_tile_26_29_2),
		.out_wire_3_3(vertical_tile_27_29_to_tile_26_29_3),
		.in_wire_3_0(vertical_tile_26_29_to_tile_27_29_0),
		.in_wire_3_1(vertical_tile_26_29_to_tile_27_29_1),
		.in_wire_3_2(vertical_tile_26_29_to_tile_27_29_2),
		.in_wire_3_3(vertical_tile_26_29_to_tile_27_29_3),
		.out_wire_1_0(vertical_tile_27_29_to_tile_28_29_0),
		.out_wire_1_1(vertical_tile_27_29_to_tile_28_29_1),
		.out_wire_1_2(vertical_tile_27_29_to_tile_28_29_2),
		.out_wire_1_3(vertical_tile_27_29_to_tile_28_29_3),
		.in_wire_1_0(vertical_tile_28_29_to_tile_27_29_0),
		.in_wire_1_1(vertical_tile_28_29_to_tile_27_29_1),
		.in_wire_1_2(vertical_tile_28_29_to_tile_27_29_2),
		.in_wire_1_3(vertical_tile_28_29_to_tile_27_29_3),
		.out_wire_2_0(horizontal_tile_27_29_to_tile_27_28_0),
		.out_wire_2_1(horizontal_tile_27_29_to_tile_27_28_1),
		.out_wire_2_2(horizontal_tile_27_29_to_tile_27_28_2),
		.out_wire_2_3(horizontal_tile_27_29_to_tile_27_28_3),
		.in_wire_2_0(horizontal_tile_27_28_to_tile_27_29_0),
		.in_wire_2_1(horizontal_tile_27_28_to_tile_27_29_1),
		.in_wire_2_2(horizontal_tile_27_28_to_tile_27_29_2),
		.in_wire_2_3(horizontal_tile_27_28_to_tile_27_29_3),
		.out_wire_0_0(horizontal_tile_27_29_to_tile_27_30_0),
		.out_wire_0_1(horizontal_tile_27_29_to_tile_27_30_1),
		.out_wire_0_2(horizontal_tile_27_29_to_tile_27_30_2),
		.out_wire_0_3(horizontal_tile_27_29_to_tile_27_30_3),
		.in_wire_0_0(horizontal_tile_27_30_to_tile_27_29_0),
		.in_wire_0_1(horizontal_tile_27_30_to_tile_27_29_1),
		.in_wire_0_2(horizontal_tile_27_30_to_tile_27_29_2),
		.in_wire_0_3(horizontal_tile_27_30_to_tile_27_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(894)
	);

	pe_tile pe_tile_27_30(
		.out_wire_3_0(vertical_tile_27_30_to_tile_26_30_0),
		.out_wire_3_1(vertical_tile_27_30_to_tile_26_30_1),
		.out_wire_3_2(vertical_tile_27_30_to_tile_26_30_2),
		.out_wire_3_3(vertical_tile_27_30_to_tile_26_30_3),
		.in_wire_3_0(vertical_tile_26_30_to_tile_27_30_0),
		.in_wire_3_1(vertical_tile_26_30_to_tile_27_30_1),
		.in_wire_3_2(vertical_tile_26_30_to_tile_27_30_2),
		.in_wire_3_3(vertical_tile_26_30_to_tile_27_30_3),
		.out_wire_1_0(vertical_tile_27_30_to_tile_28_30_0),
		.out_wire_1_1(vertical_tile_27_30_to_tile_28_30_1),
		.out_wire_1_2(vertical_tile_27_30_to_tile_28_30_2),
		.out_wire_1_3(vertical_tile_27_30_to_tile_28_30_3),
		.in_wire_1_0(vertical_tile_28_30_to_tile_27_30_0),
		.in_wire_1_1(vertical_tile_28_30_to_tile_27_30_1),
		.in_wire_1_2(vertical_tile_28_30_to_tile_27_30_2),
		.in_wire_1_3(vertical_tile_28_30_to_tile_27_30_3),
		.out_wire_2_0(horizontal_tile_27_30_to_tile_27_29_0),
		.out_wire_2_1(horizontal_tile_27_30_to_tile_27_29_1),
		.out_wire_2_2(horizontal_tile_27_30_to_tile_27_29_2),
		.out_wire_2_3(horizontal_tile_27_30_to_tile_27_29_3),
		.in_wire_2_0(horizontal_tile_27_29_to_tile_27_30_0),
		.in_wire_2_1(horizontal_tile_27_29_to_tile_27_30_1),
		.in_wire_2_2(horizontal_tile_27_29_to_tile_27_30_2),
		.in_wire_2_3(horizontal_tile_27_29_to_tile_27_30_3),
		.out_wire_0_0(horizontal_tile_27_30_to_tile_27_31_0),
		.out_wire_0_1(horizontal_tile_27_30_to_tile_27_31_1),
		.out_wire_0_2(horizontal_tile_27_30_to_tile_27_31_2),
		.out_wire_0_3(horizontal_tile_27_30_to_tile_27_31_3),
		.in_wire_0_0(horizontal_tile_27_31_to_tile_27_30_0),
		.in_wire_0_1(horizontal_tile_27_31_to_tile_27_30_1),
		.in_wire_0_2(horizontal_tile_27_31_to_tile_27_30_2),
		.in_wire_0_3(horizontal_tile_27_31_to_tile_27_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(895)
	);

	pe_tile_right pe_tile_27_31(
		.out_wire_3_0(vertical_tile_27_31_to_tile_26_31_0),
		.out_wire_3_1(vertical_tile_27_31_to_tile_26_31_1),
		.out_wire_3_2(vertical_tile_27_31_to_tile_26_31_2),
		.out_wire_3_3(vertical_tile_27_31_to_tile_26_31_3),
		.in_wire_3_0(vertical_tile_26_31_to_tile_27_31_0),
		.in_wire_3_1(vertical_tile_26_31_to_tile_27_31_1),
		.in_wire_3_2(vertical_tile_26_31_to_tile_27_31_2),
		.in_wire_3_3(vertical_tile_26_31_to_tile_27_31_3),
		.out_wire_1_0(vertical_tile_27_31_to_tile_28_31_0),
		.out_wire_1_1(vertical_tile_27_31_to_tile_28_31_1),
		.out_wire_1_2(vertical_tile_27_31_to_tile_28_31_2),
		.out_wire_1_3(vertical_tile_27_31_to_tile_28_31_3),
		.in_wire_1_0(vertical_tile_28_31_to_tile_27_31_0),
		.in_wire_1_1(vertical_tile_28_31_to_tile_27_31_1),
		.in_wire_1_2(vertical_tile_28_31_to_tile_27_31_2),
		.in_wire_1_3(vertical_tile_28_31_to_tile_27_31_3),
		.out_wire_2_0(horizontal_tile_27_31_to_tile_27_30_0),
		.out_wire_2_1(horizontal_tile_27_31_to_tile_27_30_1),
		.out_wire_2_2(horizontal_tile_27_31_to_tile_27_30_2),
		.out_wire_2_3(horizontal_tile_27_31_to_tile_27_30_3),
		.in_wire_2_0(horizontal_tile_27_30_to_tile_27_31_0),
		.in_wire_2_1(horizontal_tile_27_30_to_tile_27_31_1),
		.in_wire_2_2(horizontal_tile_27_30_to_tile_27_31_2),
		.in_wire_2_3(horizontal_tile_27_30_to_tile_27_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(896)
	);

	pe_tile_left pe_tile_28_0(
		.out_wire_3_0(vertical_tile_28_0_to_tile_27_0_0),
		.out_wire_3_1(vertical_tile_28_0_to_tile_27_0_1),
		.out_wire_3_2(vertical_tile_28_0_to_tile_27_0_2),
		.out_wire_3_3(vertical_tile_28_0_to_tile_27_0_3),
		.in_wire_3_0(vertical_tile_27_0_to_tile_28_0_0),
		.in_wire_3_1(vertical_tile_27_0_to_tile_28_0_1),
		.in_wire_3_2(vertical_tile_27_0_to_tile_28_0_2),
		.in_wire_3_3(vertical_tile_27_0_to_tile_28_0_3),
		.out_wire_1_0(vertical_tile_28_0_to_tile_29_0_0),
		.out_wire_1_1(vertical_tile_28_0_to_tile_29_0_1),
		.out_wire_1_2(vertical_tile_28_0_to_tile_29_0_2),
		.out_wire_1_3(vertical_tile_28_0_to_tile_29_0_3),
		.in_wire_1_0(vertical_tile_29_0_to_tile_28_0_0),
		.in_wire_1_1(vertical_tile_29_0_to_tile_28_0_1),
		.in_wire_1_2(vertical_tile_29_0_to_tile_28_0_2),
		.in_wire_1_3(vertical_tile_29_0_to_tile_28_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_28_0_to_tile_28_1_0),
		.out_wire_0_1(horizontal_tile_28_0_to_tile_28_1_1),
		.out_wire_0_2(horizontal_tile_28_0_to_tile_28_1_2),
		.out_wire_0_3(horizontal_tile_28_0_to_tile_28_1_3),
		.in_wire_0_0(horizontal_tile_28_1_to_tile_28_0_0),
		.in_wire_0_1(horizontal_tile_28_1_to_tile_28_0_1),
		.in_wire_0_2(horizontal_tile_28_1_to_tile_28_0_2),
		.in_wire_0_3(horizontal_tile_28_1_to_tile_28_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(897)
	);

	pe_tile pe_tile_28_1(
		.out_wire_3_0(vertical_tile_28_1_to_tile_27_1_0),
		.out_wire_3_1(vertical_tile_28_1_to_tile_27_1_1),
		.out_wire_3_2(vertical_tile_28_1_to_tile_27_1_2),
		.out_wire_3_3(vertical_tile_28_1_to_tile_27_1_3),
		.in_wire_3_0(vertical_tile_27_1_to_tile_28_1_0),
		.in_wire_3_1(vertical_tile_27_1_to_tile_28_1_1),
		.in_wire_3_2(vertical_tile_27_1_to_tile_28_1_2),
		.in_wire_3_3(vertical_tile_27_1_to_tile_28_1_3),
		.out_wire_1_0(vertical_tile_28_1_to_tile_29_1_0),
		.out_wire_1_1(vertical_tile_28_1_to_tile_29_1_1),
		.out_wire_1_2(vertical_tile_28_1_to_tile_29_1_2),
		.out_wire_1_3(vertical_tile_28_1_to_tile_29_1_3),
		.in_wire_1_0(vertical_tile_29_1_to_tile_28_1_0),
		.in_wire_1_1(vertical_tile_29_1_to_tile_28_1_1),
		.in_wire_1_2(vertical_tile_29_1_to_tile_28_1_2),
		.in_wire_1_3(vertical_tile_29_1_to_tile_28_1_3),
		.out_wire_2_0(horizontal_tile_28_1_to_tile_28_0_0),
		.out_wire_2_1(horizontal_tile_28_1_to_tile_28_0_1),
		.out_wire_2_2(horizontal_tile_28_1_to_tile_28_0_2),
		.out_wire_2_3(horizontal_tile_28_1_to_tile_28_0_3),
		.in_wire_2_0(horizontal_tile_28_0_to_tile_28_1_0),
		.in_wire_2_1(horizontal_tile_28_0_to_tile_28_1_1),
		.in_wire_2_2(horizontal_tile_28_0_to_tile_28_1_2),
		.in_wire_2_3(horizontal_tile_28_0_to_tile_28_1_3),
		.out_wire_0_0(horizontal_tile_28_1_to_tile_28_2_0),
		.out_wire_0_1(horizontal_tile_28_1_to_tile_28_2_1),
		.out_wire_0_2(horizontal_tile_28_1_to_tile_28_2_2),
		.out_wire_0_3(horizontal_tile_28_1_to_tile_28_2_3),
		.in_wire_0_0(horizontal_tile_28_2_to_tile_28_1_0),
		.in_wire_0_1(horizontal_tile_28_2_to_tile_28_1_1),
		.in_wire_0_2(horizontal_tile_28_2_to_tile_28_1_2),
		.in_wire_0_3(horizontal_tile_28_2_to_tile_28_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(898)
	);

	pe_tile pe_tile_28_2(
		.out_wire_3_0(vertical_tile_28_2_to_tile_27_2_0),
		.out_wire_3_1(vertical_tile_28_2_to_tile_27_2_1),
		.out_wire_3_2(vertical_tile_28_2_to_tile_27_2_2),
		.out_wire_3_3(vertical_tile_28_2_to_tile_27_2_3),
		.in_wire_3_0(vertical_tile_27_2_to_tile_28_2_0),
		.in_wire_3_1(vertical_tile_27_2_to_tile_28_2_1),
		.in_wire_3_2(vertical_tile_27_2_to_tile_28_2_2),
		.in_wire_3_3(vertical_tile_27_2_to_tile_28_2_3),
		.out_wire_1_0(vertical_tile_28_2_to_tile_29_2_0),
		.out_wire_1_1(vertical_tile_28_2_to_tile_29_2_1),
		.out_wire_1_2(vertical_tile_28_2_to_tile_29_2_2),
		.out_wire_1_3(vertical_tile_28_2_to_tile_29_2_3),
		.in_wire_1_0(vertical_tile_29_2_to_tile_28_2_0),
		.in_wire_1_1(vertical_tile_29_2_to_tile_28_2_1),
		.in_wire_1_2(vertical_tile_29_2_to_tile_28_2_2),
		.in_wire_1_3(vertical_tile_29_2_to_tile_28_2_3),
		.out_wire_2_0(horizontal_tile_28_2_to_tile_28_1_0),
		.out_wire_2_1(horizontal_tile_28_2_to_tile_28_1_1),
		.out_wire_2_2(horizontal_tile_28_2_to_tile_28_1_2),
		.out_wire_2_3(horizontal_tile_28_2_to_tile_28_1_3),
		.in_wire_2_0(horizontal_tile_28_1_to_tile_28_2_0),
		.in_wire_2_1(horizontal_tile_28_1_to_tile_28_2_1),
		.in_wire_2_2(horizontal_tile_28_1_to_tile_28_2_2),
		.in_wire_2_3(horizontal_tile_28_1_to_tile_28_2_3),
		.out_wire_0_0(horizontal_tile_28_2_to_tile_28_3_0),
		.out_wire_0_1(horizontal_tile_28_2_to_tile_28_3_1),
		.out_wire_0_2(horizontal_tile_28_2_to_tile_28_3_2),
		.out_wire_0_3(horizontal_tile_28_2_to_tile_28_3_3),
		.in_wire_0_0(horizontal_tile_28_3_to_tile_28_2_0),
		.in_wire_0_1(horizontal_tile_28_3_to_tile_28_2_1),
		.in_wire_0_2(horizontal_tile_28_3_to_tile_28_2_2),
		.in_wire_0_3(horizontal_tile_28_3_to_tile_28_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(899)
	);

	pe_tile pe_tile_28_3(
		.out_wire_3_0(vertical_tile_28_3_to_tile_27_3_0),
		.out_wire_3_1(vertical_tile_28_3_to_tile_27_3_1),
		.out_wire_3_2(vertical_tile_28_3_to_tile_27_3_2),
		.out_wire_3_3(vertical_tile_28_3_to_tile_27_3_3),
		.in_wire_3_0(vertical_tile_27_3_to_tile_28_3_0),
		.in_wire_3_1(vertical_tile_27_3_to_tile_28_3_1),
		.in_wire_3_2(vertical_tile_27_3_to_tile_28_3_2),
		.in_wire_3_3(vertical_tile_27_3_to_tile_28_3_3),
		.out_wire_1_0(vertical_tile_28_3_to_tile_29_3_0),
		.out_wire_1_1(vertical_tile_28_3_to_tile_29_3_1),
		.out_wire_1_2(vertical_tile_28_3_to_tile_29_3_2),
		.out_wire_1_3(vertical_tile_28_3_to_tile_29_3_3),
		.in_wire_1_0(vertical_tile_29_3_to_tile_28_3_0),
		.in_wire_1_1(vertical_tile_29_3_to_tile_28_3_1),
		.in_wire_1_2(vertical_tile_29_3_to_tile_28_3_2),
		.in_wire_1_3(vertical_tile_29_3_to_tile_28_3_3),
		.out_wire_2_0(horizontal_tile_28_3_to_tile_28_2_0),
		.out_wire_2_1(horizontal_tile_28_3_to_tile_28_2_1),
		.out_wire_2_2(horizontal_tile_28_3_to_tile_28_2_2),
		.out_wire_2_3(horizontal_tile_28_3_to_tile_28_2_3),
		.in_wire_2_0(horizontal_tile_28_2_to_tile_28_3_0),
		.in_wire_2_1(horizontal_tile_28_2_to_tile_28_3_1),
		.in_wire_2_2(horizontal_tile_28_2_to_tile_28_3_2),
		.in_wire_2_3(horizontal_tile_28_2_to_tile_28_3_3),
		.out_wire_0_0(horizontal_tile_28_3_to_tile_28_4_0),
		.out_wire_0_1(horizontal_tile_28_3_to_tile_28_4_1),
		.out_wire_0_2(horizontal_tile_28_3_to_tile_28_4_2),
		.out_wire_0_3(horizontal_tile_28_3_to_tile_28_4_3),
		.in_wire_0_0(horizontal_tile_28_4_to_tile_28_3_0),
		.in_wire_0_1(horizontal_tile_28_4_to_tile_28_3_1),
		.in_wire_0_2(horizontal_tile_28_4_to_tile_28_3_2),
		.in_wire_0_3(horizontal_tile_28_4_to_tile_28_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(900)
	);

	pe_tile pe_tile_28_4(
		.out_wire_3_0(vertical_tile_28_4_to_tile_27_4_0),
		.out_wire_3_1(vertical_tile_28_4_to_tile_27_4_1),
		.out_wire_3_2(vertical_tile_28_4_to_tile_27_4_2),
		.out_wire_3_3(vertical_tile_28_4_to_tile_27_4_3),
		.in_wire_3_0(vertical_tile_27_4_to_tile_28_4_0),
		.in_wire_3_1(vertical_tile_27_4_to_tile_28_4_1),
		.in_wire_3_2(vertical_tile_27_4_to_tile_28_4_2),
		.in_wire_3_3(vertical_tile_27_4_to_tile_28_4_3),
		.out_wire_1_0(vertical_tile_28_4_to_tile_29_4_0),
		.out_wire_1_1(vertical_tile_28_4_to_tile_29_4_1),
		.out_wire_1_2(vertical_tile_28_4_to_tile_29_4_2),
		.out_wire_1_3(vertical_tile_28_4_to_tile_29_4_3),
		.in_wire_1_0(vertical_tile_29_4_to_tile_28_4_0),
		.in_wire_1_1(vertical_tile_29_4_to_tile_28_4_1),
		.in_wire_1_2(vertical_tile_29_4_to_tile_28_4_2),
		.in_wire_1_3(vertical_tile_29_4_to_tile_28_4_3),
		.out_wire_2_0(horizontal_tile_28_4_to_tile_28_3_0),
		.out_wire_2_1(horizontal_tile_28_4_to_tile_28_3_1),
		.out_wire_2_2(horizontal_tile_28_4_to_tile_28_3_2),
		.out_wire_2_3(horizontal_tile_28_4_to_tile_28_3_3),
		.in_wire_2_0(horizontal_tile_28_3_to_tile_28_4_0),
		.in_wire_2_1(horizontal_tile_28_3_to_tile_28_4_1),
		.in_wire_2_2(horizontal_tile_28_3_to_tile_28_4_2),
		.in_wire_2_3(horizontal_tile_28_3_to_tile_28_4_3),
		.out_wire_0_0(horizontal_tile_28_4_to_tile_28_5_0),
		.out_wire_0_1(horizontal_tile_28_4_to_tile_28_5_1),
		.out_wire_0_2(horizontal_tile_28_4_to_tile_28_5_2),
		.out_wire_0_3(horizontal_tile_28_4_to_tile_28_5_3),
		.in_wire_0_0(horizontal_tile_28_5_to_tile_28_4_0),
		.in_wire_0_1(horizontal_tile_28_5_to_tile_28_4_1),
		.in_wire_0_2(horizontal_tile_28_5_to_tile_28_4_2),
		.in_wire_0_3(horizontal_tile_28_5_to_tile_28_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(901)
	);

	pe_tile pe_tile_28_5(
		.out_wire_3_0(vertical_tile_28_5_to_tile_27_5_0),
		.out_wire_3_1(vertical_tile_28_5_to_tile_27_5_1),
		.out_wire_3_2(vertical_tile_28_5_to_tile_27_5_2),
		.out_wire_3_3(vertical_tile_28_5_to_tile_27_5_3),
		.in_wire_3_0(vertical_tile_27_5_to_tile_28_5_0),
		.in_wire_3_1(vertical_tile_27_5_to_tile_28_5_1),
		.in_wire_3_2(vertical_tile_27_5_to_tile_28_5_2),
		.in_wire_3_3(vertical_tile_27_5_to_tile_28_5_3),
		.out_wire_1_0(vertical_tile_28_5_to_tile_29_5_0),
		.out_wire_1_1(vertical_tile_28_5_to_tile_29_5_1),
		.out_wire_1_2(vertical_tile_28_5_to_tile_29_5_2),
		.out_wire_1_3(vertical_tile_28_5_to_tile_29_5_3),
		.in_wire_1_0(vertical_tile_29_5_to_tile_28_5_0),
		.in_wire_1_1(vertical_tile_29_5_to_tile_28_5_1),
		.in_wire_1_2(vertical_tile_29_5_to_tile_28_5_2),
		.in_wire_1_3(vertical_tile_29_5_to_tile_28_5_3),
		.out_wire_2_0(horizontal_tile_28_5_to_tile_28_4_0),
		.out_wire_2_1(horizontal_tile_28_5_to_tile_28_4_1),
		.out_wire_2_2(horizontal_tile_28_5_to_tile_28_4_2),
		.out_wire_2_3(horizontal_tile_28_5_to_tile_28_4_3),
		.in_wire_2_0(horizontal_tile_28_4_to_tile_28_5_0),
		.in_wire_2_1(horizontal_tile_28_4_to_tile_28_5_1),
		.in_wire_2_2(horizontal_tile_28_4_to_tile_28_5_2),
		.in_wire_2_3(horizontal_tile_28_4_to_tile_28_5_3),
		.out_wire_0_0(horizontal_tile_28_5_to_tile_28_6_0),
		.out_wire_0_1(horizontal_tile_28_5_to_tile_28_6_1),
		.out_wire_0_2(horizontal_tile_28_5_to_tile_28_6_2),
		.out_wire_0_3(horizontal_tile_28_5_to_tile_28_6_3),
		.in_wire_0_0(horizontal_tile_28_6_to_tile_28_5_0),
		.in_wire_0_1(horizontal_tile_28_6_to_tile_28_5_1),
		.in_wire_0_2(horizontal_tile_28_6_to_tile_28_5_2),
		.in_wire_0_3(horizontal_tile_28_6_to_tile_28_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(902)
	);

	pe_tile pe_tile_28_6(
		.out_wire_3_0(vertical_tile_28_6_to_tile_27_6_0),
		.out_wire_3_1(vertical_tile_28_6_to_tile_27_6_1),
		.out_wire_3_2(vertical_tile_28_6_to_tile_27_6_2),
		.out_wire_3_3(vertical_tile_28_6_to_tile_27_6_3),
		.in_wire_3_0(vertical_tile_27_6_to_tile_28_6_0),
		.in_wire_3_1(vertical_tile_27_6_to_tile_28_6_1),
		.in_wire_3_2(vertical_tile_27_6_to_tile_28_6_2),
		.in_wire_3_3(vertical_tile_27_6_to_tile_28_6_3),
		.out_wire_1_0(vertical_tile_28_6_to_tile_29_6_0),
		.out_wire_1_1(vertical_tile_28_6_to_tile_29_6_1),
		.out_wire_1_2(vertical_tile_28_6_to_tile_29_6_2),
		.out_wire_1_3(vertical_tile_28_6_to_tile_29_6_3),
		.in_wire_1_0(vertical_tile_29_6_to_tile_28_6_0),
		.in_wire_1_1(vertical_tile_29_6_to_tile_28_6_1),
		.in_wire_1_2(vertical_tile_29_6_to_tile_28_6_2),
		.in_wire_1_3(vertical_tile_29_6_to_tile_28_6_3),
		.out_wire_2_0(horizontal_tile_28_6_to_tile_28_5_0),
		.out_wire_2_1(horizontal_tile_28_6_to_tile_28_5_1),
		.out_wire_2_2(horizontal_tile_28_6_to_tile_28_5_2),
		.out_wire_2_3(horizontal_tile_28_6_to_tile_28_5_3),
		.in_wire_2_0(horizontal_tile_28_5_to_tile_28_6_0),
		.in_wire_2_1(horizontal_tile_28_5_to_tile_28_6_1),
		.in_wire_2_2(horizontal_tile_28_5_to_tile_28_6_2),
		.in_wire_2_3(horizontal_tile_28_5_to_tile_28_6_3),
		.out_wire_0_0(horizontal_tile_28_6_to_tile_28_7_0),
		.out_wire_0_1(horizontal_tile_28_6_to_tile_28_7_1),
		.out_wire_0_2(horizontal_tile_28_6_to_tile_28_7_2),
		.out_wire_0_3(horizontal_tile_28_6_to_tile_28_7_3),
		.in_wire_0_0(horizontal_tile_28_7_to_tile_28_6_0),
		.in_wire_0_1(horizontal_tile_28_7_to_tile_28_6_1),
		.in_wire_0_2(horizontal_tile_28_7_to_tile_28_6_2),
		.in_wire_0_3(horizontal_tile_28_7_to_tile_28_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(903)
	);

	pe_tile pe_tile_28_7(
		.out_wire_3_0(vertical_tile_28_7_to_tile_27_7_0),
		.out_wire_3_1(vertical_tile_28_7_to_tile_27_7_1),
		.out_wire_3_2(vertical_tile_28_7_to_tile_27_7_2),
		.out_wire_3_3(vertical_tile_28_7_to_tile_27_7_3),
		.in_wire_3_0(vertical_tile_27_7_to_tile_28_7_0),
		.in_wire_3_1(vertical_tile_27_7_to_tile_28_7_1),
		.in_wire_3_2(vertical_tile_27_7_to_tile_28_7_2),
		.in_wire_3_3(vertical_tile_27_7_to_tile_28_7_3),
		.out_wire_1_0(vertical_tile_28_7_to_tile_29_7_0),
		.out_wire_1_1(vertical_tile_28_7_to_tile_29_7_1),
		.out_wire_1_2(vertical_tile_28_7_to_tile_29_7_2),
		.out_wire_1_3(vertical_tile_28_7_to_tile_29_7_3),
		.in_wire_1_0(vertical_tile_29_7_to_tile_28_7_0),
		.in_wire_1_1(vertical_tile_29_7_to_tile_28_7_1),
		.in_wire_1_2(vertical_tile_29_7_to_tile_28_7_2),
		.in_wire_1_3(vertical_tile_29_7_to_tile_28_7_3),
		.out_wire_2_0(horizontal_tile_28_7_to_tile_28_6_0),
		.out_wire_2_1(horizontal_tile_28_7_to_tile_28_6_1),
		.out_wire_2_2(horizontal_tile_28_7_to_tile_28_6_2),
		.out_wire_2_3(horizontal_tile_28_7_to_tile_28_6_3),
		.in_wire_2_0(horizontal_tile_28_6_to_tile_28_7_0),
		.in_wire_2_1(horizontal_tile_28_6_to_tile_28_7_1),
		.in_wire_2_2(horizontal_tile_28_6_to_tile_28_7_2),
		.in_wire_2_3(horizontal_tile_28_6_to_tile_28_7_3),
		.out_wire_0_0(horizontal_tile_28_7_to_tile_28_8_0),
		.out_wire_0_1(horizontal_tile_28_7_to_tile_28_8_1),
		.out_wire_0_2(horizontal_tile_28_7_to_tile_28_8_2),
		.out_wire_0_3(horizontal_tile_28_7_to_tile_28_8_3),
		.in_wire_0_0(horizontal_tile_28_8_to_tile_28_7_0),
		.in_wire_0_1(horizontal_tile_28_8_to_tile_28_7_1),
		.in_wire_0_2(horizontal_tile_28_8_to_tile_28_7_2),
		.in_wire_0_3(horizontal_tile_28_8_to_tile_28_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(904)
	);

	pe_tile pe_tile_28_8(
		.out_wire_3_0(vertical_tile_28_8_to_tile_27_8_0),
		.out_wire_3_1(vertical_tile_28_8_to_tile_27_8_1),
		.out_wire_3_2(vertical_tile_28_8_to_tile_27_8_2),
		.out_wire_3_3(vertical_tile_28_8_to_tile_27_8_3),
		.in_wire_3_0(vertical_tile_27_8_to_tile_28_8_0),
		.in_wire_3_1(vertical_tile_27_8_to_tile_28_8_1),
		.in_wire_3_2(vertical_tile_27_8_to_tile_28_8_2),
		.in_wire_3_3(vertical_tile_27_8_to_tile_28_8_3),
		.out_wire_1_0(vertical_tile_28_8_to_tile_29_8_0),
		.out_wire_1_1(vertical_tile_28_8_to_tile_29_8_1),
		.out_wire_1_2(vertical_tile_28_8_to_tile_29_8_2),
		.out_wire_1_3(vertical_tile_28_8_to_tile_29_8_3),
		.in_wire_1_0(vertical_tile_29_8_to_tile_28_8_0),
		.in_wire_1_1(vertical_tile_29_8_to_tile_28_8_1),
		.in_wire_1_2(vertical_tile_29_8_to_tile_28_8_2),
		.in_wire_1_3(vertical_tile_29_8_to_tile_28_8_3),
		.out_wire_2_0(horizontal_tile_28_8_to_tile_28_7_0),
		.out_wire_2_1(horizontal_tile_28_8_to_tile_28_7_1),
		.out_wire_2_2(horizontal_tile_28_8_to_tile_28_7_2),
		.out_wire_2_3(horizontal_tile_28_8_to_tile_28_7_3),
		.in_wire_2_0(horizontal_tile_28_7_to_tile_28_8_0),
		.in_wire_2_1(horizontal_tile_28_7_to_tile_28_8_1),
		.in_wire_2_2(horizontal_tile_28_7_to_tile_28_8_2),
		.in_wire_2_3(horizontal_tile_28_7_to_tile_28_8_3),
		.out_wire_0_0(horizontal_tile_28_8_to_tile_28_9_0),
		.out_wire_0_1(horizontal_tile_28_8_to_tile_28_9_1),
		.out_wire_0_2(horizontal_tile_28_8_to_tile_28_9_2),
		.out_wire_0_3(horizontal_tile_28_8_to_tile_28_9_3),
		.in_wire_0_0(horizontal_tile_28_9_to_tile_28_8_0),
		.in_wire_0_1(horizontal_tile_28_9_to_tile_28_8_1),
		.in_wire_0_2(horizontal_tile_28_9_to_tile_28_8_2),
		.in_wire_0_3(horizontal_tile_28_9_to_tile_28_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(905)
	);

	pe_tile pe_tile_28_9(
		.out_wire_3_0(vertical_tile_28_9_to_tile_27_9_0),
		.out_wire_3_1(vertical_tile_28_9_to_tile_27_9_1),
		.out_wire_3_2(vertical_tile_28_9_to_tile_27_9_2),
		.out_wire_3_3(vertical_tile_28_9_to_tile_27_9_3),
		.in_wire_3_0(vertical_tile_27_9_to_tile_28_9_0),
		.in_wire_3_1(vertical_tile_27_9_to_tile_28_9_1),
		.in_wire_3_2(vertical_tile_27_9_to_tile_28_9_2),
		.in_wire_3_3(vertical_tile_27_9_to_tile_28_9_3),
		.out_wire_1_0(vertical_tile_28_9_to_tile_29_9_0),
		.out_wire_1_1(vertical_tile_28_9_to_tile_29_9_1),
		.out_wire_1_2(vertical_tile_28_9_to_tile_29_9_2),
		.out_wire_1_3(vertical_tile_28_9_to_tile_29_9_3),
		.in_wire_1_0(vertical_tile_29_9_to_tile_28_9_0),
		.in_wire_1_1(vertical_tile_29_9_to_tile_28_9_1),
		.in_wire_1_2(vertical_tile_29_9_to_tile_28_9_2),
		.in_wire_1_3(vertical_tile_29_9_to_tile_28_9_3),
		.out_wire_2_0(horizontal_tile_28_9_to_tile_28_8_0),
		.out_wire_2_1(horizontal_tile_28_9_to_tile_28_8_1),
		.out_wire_2_2(horizontal_tile_28_9_to_tile_28_8_2),
		.out_wire_2_3(horizontal_tile_28_9_to_tile_28_8_3),
		.in_wire_2_0(horizontal_tile_28_8_to_tile_28_9_0),
		.in_wire_2_1(horizontal_tile_28_8_to_tile_28_9_1),
		.in_wire_2_2(horizontal_tile_28_8_to_tile_28_9_2),
		.in_wire_2_3(horizontal_tile_28_8_to_tile_28_9_3),
		.out_wire_0_0(horizontal_tile_28_9_to_tile_28_10_0),
		.out_wire_0_1(horizontal_tile_28_9_to_tile_28_10_1),
		.out_wire_0_2(horizontal_tile_28_9_to_tile_28_10_2),
		.out_wire_0_3(horizontal_tile_28_9_to_tile_28_10_3),
		.in_wire_0_0(horizontal_tile_28_10_to_tile_28_9_0),
		.in_wire_0_1(horizontal_tile_28_10_to_tile_28_9_1),
		.in_wire_0_2(horizontal_tile_28_10_to_tile_28_9_2),
		.in_wire_0_3(horizontal_tile_28_10_to_tile_28_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(906)
	);

	pe_tile pe_tile_28_10(
		.out_wire_3_0(vertical_tile_28_10_to_tile_27_10_0),
		.out_wire_3_1(vertical_tile_28_10_to_tile_27_10_1),
		.out_wire_3_2(vertical_tile_28_10_to_tile_27_10_2),
		.out_wire_3_3(vertical_tile_28_10_to_tile_27_10_3),
		.in_wire_3_0(vertical_tile_27_10_to_tile_28_10_0),
		.in_wire_3_1(vertical_tile_27_10_to_tile_28_10_1),
		.in_wire_3_2(vertical_tile_27_10_to_tile_28_10_2),
		.in_wire_3_3(vertical_tile_27_10_to_tile_28_10_3),
		.out_wire_1_0(vertical_tile_28_10_to_tile_29_10_0),
		.out_wire_1_1(vertical_tile_28_10_to_tile_29_10_1),
		.out_wire_1_2(vertical_tile_28_10_to_tile_29_10_2),
		.out_wire_1_3(vertical_tile_28_10_to_tile_29_10_3),
		.in_wire_1_0(vertical_tile_29_10_to_tile_28_10_0),
		.in_wire_1_1(vertical_tile_29_10_to_tile_28_10_1),
		.in_wire_1_2(vertical_tile_29_10_to_tile_28_10_2),
		.in_wire_1_3(vertical_tile_29_10_to_tile_28_10_3),
		.out_wire_2_0(horizontal_tile_28_10_to_tile_28_9_0),
		.out_wire_2_1(horizontal_tile_28_10_to_tile_28_9_1),
		.out_wire_2_2(horizontal_tile_28_10_to_tile_28_9_2),
		.out_wire_2_3(horizontal_tile_28_10_to_tile_28_9_3),
		.in_wire_2_0(horizontal_tile_28_9_to_tile_28_10_0),
		.in_wire_2_1(horizontal_tile_28_9_to_tile_28_10_1),
		.in_wire_2_2(horizontal_tile_28_9_to_tile_28_10_2),
		.in_wire_2_3(horizontal_tile_28_9_to_tile_28_10_3),
		.out_wire_0_0(horizontal_tile_28_10_to_tile_28_11_0),
		.out_wire_0_1(horizontal_tile_28_10_to_tile_28_11_1),
		.out_wire_0_2(horizontal_tile_28_10_to_tile_28_11_2),
		.out_wire_0_3(horizontal_tile_28_10_to_tile_28_11_3),
		.in_wire_0_0(horizontal_tile_28_11_to_tile_28_10_0),
		.in_wire_0_1(horizontal_tile_28_11_to_tile_28_10_1),
		.in_wire_0_2(horizontal_tile_28_11_to_tile_28_10_2),
		.in_wire_0_3(horizontal_tile_28_11_to_tile_28_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(907)
	);

	pe_tile pe_tile_28_11(
		.out_wire_3_0(vertical_tile_28_11_to_tile_27_11_0),
		.out_wire_3_1(vertical_tile_28_11_to_tile_27_11_1),
		.out_wire_3_2(vertical_tile_28_11_to_tile_27_11_2),
		.out_wire_3_3(vertical_tile_28_11_to_tile_27_11_3),
		.in_wire_3_0(vertical_tile_27_11_to_tile_28_11_0),
		.in_wire_3_1(vertical_tile_27_11_to_tile_28_11_1),
		.in_wire_3_2(vertical_tile_27_11_to_tile_28_11_2),
		.in_wire_3_3(vertical_tile_27_11_to_tile_28_11_3),
		.out_wire_1_0(vertical_tile_28_11_to_tile_29_11_0),
		.out_wire_1_1(vertical_tile_28_11_to_tile_29_11_1),
		.out_wire_1_2(vertical_tile_28_11_to_tile_29_11_2),
		.out_wire_1_3(vertical_tile_28_11_to_tile_29_11_3),
		.in_wire_1_0(vertical_tile_29_11_to_tile_28_11_0),
		.in_wire_1_1(vertical_tile_29_11_to_tile_28_11_1),
		.in_wire_1_2(vertical_tile_29_11_to_tile_28_11_2),
		.in_wire_1_3(vertical_tile_29_11_to_tile_28_11_3),
		.out_wire_2_0(horizontal_tile_28_11_to_tile_28_10_0),
		.out_wire_2_1(horizontal_tile_28_11_to_tile_28_10_1),
		.out_wire_2_2(horizontal_tile_28_11_to_tile_28_10_2),
		.out_wire_2_3(horizontal_tile_28_11_to_tile_28_10_3),
		.in_wire_2_0(horizontal_tile_28_10_to_tile_28_11_0),
		.in_wire_2_1(horizontal_tile_28_10_to_tile_28_11_1),
		.in_wire_2_2(horizontal_tile_28_10_to_tile_28_11_2),
		.in_wire_2_3(horizontal_tile_28_10_to_tile_28_11_3),
		.out_wire_0_0(horizontal_tile_28_11_to_tile_28_12_0),
		.out_wire_0_1(horizontal_tile_28_11_to_tile_28_12_1),
		.out_wire_0_2(horizontal_tile_28_11_to_tile_28_12_2),
		.out_wire_0_3(horizontal_tile_28_11_to_tile_28_12_3),
		.in_wire_0_0(horizontal_tile_28_12_to_tile_28_11_0),
		.in_wire_0_1(horizontal_tile_28_12_to_tile_28_11_1),
		.in_wire_0_2(horizontal_tile_28_12_to_tile_28_11_2),
		.in_wire_0_3(horizontal_tile_28_12_to_tile_28_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(908)
	);

	pe_tile pe_tile_28_12(
		.out_wire_3_0(vertical_tile_28_12_to_tile_27_12_0),
		.out_wire_3_1(vertical_tile_28_12_to_tile_27_12_1),
		.out_wire_3_2(vertical_tile_28_12_to_tile_27_12_2),
		.out_wire_3_3(vertical_tile_28_12_to_tile_27_12_3),
		.in_wire_3_0(vertical_tile_27_12_to_tile_28_12_0),
		.in_wire_3_1(vertical_tile_27_12_to_tile_28_12_1),
		.in_wire_3_2(vertical_tile_27_12_to_tile_28_12_2),
		.in_wire_3_3(vertical_tile_27_12_to_tile_28_12_3),
		.out_wire_1_0(vertical_tile_28_12_to_tile_29_12_0),
		.out_wire_1_1(vertical_tile_28_12_to_tile_29_12_1),
		.out_wire_1_2(vertical_tile_28_12_to_tile_29_12_2),
		.out_wire_1_3(vertical_tile_28_12_to_tile_29_12_3),
		.in_wire_1_0(vertical_tile_29_12_to_tile_28_12_0),
		.in_wire_1_1(vertical_tile_29_12_to_tile_28_12_1),
		.in_wire_1_2(vertical_tile_29_12_to_tile_28_12_2),
		.in_wire_1_3(vertical_tile_29_12_to_tile_28_12_3),
		.out_wire_2_0(horizontal_tile_28_12_to_tile_28_11_0),
		.out_wire_2_1(horizontal_tile_28_12_to_tile_28_11_1),
		.out_wire_2_2(horizontal_tile_28_12_to_tile_28_11_2),
		.out_wire_2_3(horizontal_tile_28_12_to_tile_28_11_3),
		.in_wire_2_0(horizontal_tile_28_11_to_tile_28_12_0),
		.in_wire_2_1(horizontal_tile_28_11_to_tile_28_12_1),
		.in_wire_2_2(horizontal_tile_28_11_to_tile_28_12_2),
		.in_wire_2_3(horizontal_tile_28_11_to_tile_28_12_3),
		.out_wire_0_0(horizontal_tile_28_12_to_tile_28_13_0),
		.out_wire_0_1(horizontal_tile_28_12_to_tile_28_13_1),
		.out_wire_0_2(horizontal_tile_28_12_to_tile_28_13_2),
		.out_wire_0_3(horizontal_tile_28_12_to_tile_28_13_3),
		.in_wire_0_0(horizontal_tile_28_13_to_tile_28_12_0),
		.in_wire_0_1(horizontal_tile_28_13_to_tile_28_12_1),
		.in_wire_0_2(horizontal_tile_28_13_to_tile_28_12_2),
		.in_wire_0_3(horizontal_tile_28_13_to_tile_28_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(909)
	);

	pe_tile pe_tile_28_13(
		.out_wire_3_0(vertical_tile_28_13_to_tile_27_13_0),
		.out_wire_3_1(vertical_tile_28_13_to_tile_27_13_1),
		.out_wire_3_2(vertical_tile_28_13_to_tile_27_13_2),
		.out_wire_3_3(vertical_tile_28_13_to_tile_27_13_3),
		.in_wire_3_0(vertical_tile_27_13_to_tile_28_13_0),
		.in_wire_3_1(vertical_tile_27_13_to_tile_28_13_1),
		.in_wire_3_2(vertical_tile_27_13_to_tile_28_13_2),
		.in_wire_3_3(vertical_tile_27_13_to_tile_28_13_3),
		.out_wire_1_0(vertical_tile_28_13_to_tile_29_13_0),
		.out_wire_1_1(vertical_tile_28_13_to_tile_29_13_1),
		.out_wire_1_2(vertical_tile_28_13_to_tile_29_13_2),
		.out_wire_1_3(vertical_tile_28_13_to_tile_29_13_3),
		.in_wire_1_0(vertical_tile_29_13_to_tile_28_13_0),
		.in_wire_1_1(vertical_tile_29_13_to_tile_28_13_1),
		.in_wire_1_2(vertical_tile_29_13_to_tile_28_13_2),
		.in_wire_1_3(vertical_tile_29_13_to_tile_28_13_3),
		.out_wire_2_0(horizontal_tile_28_13_to_tile_28_12_0),
		.out_wire_2_1(horizontal_tile_28_13_to_tile_28_12_1),
		.out_wire_2_2(horizontal_tile_28_13_to_tile_28_12_2),
		.out_wire_2_3(horizontal_tile_28_13_to_tile_28_12_3),
		.in_wire_2_0(horizontal_tile_28_12_to_tile_28_13_0),
		.in_wire_2_1(horizontal_tile_28_12_to_tile_28_13_1),
		.in_wire_2_2(horizontal_tile_28_12_to_tile_28_13_2),
		.in_wire_2_3(horizontal_tile_28_12_to_tile_28_13_3),
		.out_wire_0_0(horizontal_tile_28_13_to_tile_28_14_0),
		.out_wire_0_1(horizontal_tile_28_13_to_tile_28_14_1),
		.out_wire_0_2(horizontal_tile_28_13_to_tile_28_14_2),
		.out_wire_0_3(horizontal_tile_28_13_to_tile_28_14_3),
		.in_wire_0_0(horizontal_tile_28_14_to_tile_28_13_0),
		.in_wire_0_1(horizontal_tile_28_14_to_tile_28_13_1),
		.in_wire_0_2(horizontal_tile_28_14_to_tile_28_13_2),
		.in_wire_0_3(horizontal_tile_28_14_to_tile_28_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(910)
	);

	pe_tile pe_tile_28_14(
		.out_wire_3_0(vertical_tile_28_14_to_tile_27_14_0),
		.out_wire_3_1(vertical_tile_28_14_to_tile_27_14_1),
		.out_wire_3_2(vertical_tile_28_14_to_tile_27_14_2),
		.out_wire_3_3(vertical_tile_28_14_to_tile_27_14_3),
		.in_wire_3_0(vertical_tile_27_14_to_tile_28_14_0),
		.in_wire_3_1(vertical_tile_27_14_to_tile_28_14_1),
		.in_wire_3_2(vertical_tile_27_14_to_tile_28_14_2),
		.in_wire_3_3(vertical_tile_27_14_to_tile_28_14_3),
		.out_wire_1_0(vertical_tile_28_14_to_tile_29_14_0),
		.out_wire_1_1(vertical_tile_28_14_to_tile_29_14_1),
		.out_wire_1_2(vertical_tile_28_14_to_tile_29_14_2),
		.out_wire_1_3(vertical_tile_28_14_to_tile_29_14_3),
		.in_wire_1_0(vertical_tile_29_14_to_tile_28_14_0),
		.in_wire_1_1(vertical_tile_29_14_to_tile_28_14_1),
		.in_wire_1_2(vertical_tile_29_14_to_tile_28_14_2),
		.in_wire_1_3(vertical_tile_29_14_to_tile_28_14_3),
		.out_wire_2_0(horizontal_tile_28_14_to_tile_28_13_0),
		.out_wire_2_1(horizontal_tile_28_14_to_tile_28_13_1),
		.out_wire_2_2(horizontal_tile_28_14_to_tile_28_13_2),
		.out_wire_2_3(horizontal_tile_28_14_to_tile_28_13_3),
		.in_wire_2_0(horizontal_tile_28_13_to_tile_28_14_0),
		.in_wire_2_1(horizontal_tile_28_13_to_tile_28_14_1),
		.in_wire_2_2(horizontal_tile_28_13_to_tile_28_14_2),
		.in_wire_2_3(horizontal_tile_28_13_to_tile_28_14_3),
		.out_wire_0_0(horizontal_tile_28_14_to_tile_28_15_0),
		.out_wire_0_1(horizontal_tile_28_14_to_tile_28_15_1),
		.out_wire_0_2(horizontal_tile_28_14_to_tile_28_15_2),
		.out_wire_0_3(horizontal_tile_28_14_to_tile_28_15_3),
		.in_wire_0_0(horizontal_tile_28_15_to_tile_28_14_0),
		.in_wire_0_1(horizontal_tile_28_15_to_tile_28_14_1),
		.in_wire_0_2(horizontal_tile_28_15_to_tile_28_14_2),
		.in_wire_0_3(horizontal_tile_28_15_to_tile_28_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(911)
	);

	pe_tile pe_tile_28_15(
		.out_wire_3_0(vertical_tile_28_15_to_tile_27_15_0),
		.out_wire_3_1(vertical_tile_28_15_to_tile_27_15_1),
		.out_wire_3_2(vertical_tile_28_15_to_tile_27_15_2),
		.out_wire_3_3(vertical_tile_28_15_to_tile_27_15_3),
		.in_wire_3_0(vertical_tile_27_15_to_tile_28_15_0),
		.in_wire_3_1(vertical_tile_27_15_to_tile_28_15_1),
		.in_wire_3_2(vertical_tile_27_15_to_tile_28_15_2),
		.in_wire_3_3(vertical_tile_27_15_to_tile_28_15_3),
		.out_wire_1_0(vertical_tile_28_15_to_tile_29_15_0),
		.out_wire_1_1(vertical_tile_28_15_to_tile_29_15_1),
		.out_wire_1_2(vertical_tile_28_15_to_tile_29_15_2),
		.out_wire_1_3(vertical_tile_28_15_to_tile_29_15_3),
		.in_wire_1_0(vertical_tile_29_15_to_tile_28_15_0),
		.in_wire_1_1(vertical_tile_29_15_to_tile_28_15_1),
		.in_wire_1_2(vertical_tile_29_15_to_tile_28_15_2),
		.in_wire_1_3(vertical_tile_29_15_to_tile_28_15_3),
		.out_wire_2_0(horizontal_tile_28_15_to_tile_28_14_0),
		.out_wire_2_1(horizontal_tile_28_15_to_tile_28_14_1),
		.out_wire_2_2(horizontal_tile_28_15_to_tile_28_14_2),
		.out_wire_2_3(horizontal_tile_28_15_to_tile_28_14_3),
		.in_wire_2_0(horizontal_tile_28_14_to_tile_28_15_0),
		.in_wire_2_1(horizontal_tile_28_14_to_tile_28_15_1),
		.in_wire_2_2(horizontal_tile_28_14_to_tile_28_15_2),
		.in_wire_2_3(horizontal_tile_28_14_to_tile_28_15_3),
		.out_wire_0_0(horizontal_tile_28_15_to_tile_28_16_0),
		.out_wire_0_1(horizontal_tile_28_15_to_tile_28_16_1),
		.out_wire_0_2(horizontal_tile_28_15_to_tile_28_16_2),
		.out_wire_0_3(horizontal_tile_28_15_to_tile_28_16_3),
		.in_wire_0_0(horizontal_tile_28_16_to_tile_28_15_0),
		.in_wire_0_1(horizontal_tile_28_16_to_tile_28_15_1),
		.in_wire_0_2(horizontal_tile_28_16_to_tile_28_15_2),
		.in_wire_0_3(horizontal_tile_28_16_to_tile_28_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(912)
	);

	pe_tile pe_tile_28_16(
		.out_wire_3_0(vertical_tile_28_16_to_tile_27_16_0),
		.out_wire_3_1(vertical_tile_28_16_to_tile_27_16_1),
		.out_wire_3_2(vertical_tile_28_16_to_tile_27_16_2),
		.out_wire_3_3(vertical_tile_28_16_to_tile_27_16_3),
		.in_wire_3_0(vertical_tile_27_16_to_tile_28_16_0),
		.in_wire_3_1(vertical_tile_27_16_to_tile_28_16_1),
		.in_wire_3_2(vertical_tile_27_16_to_tile_28_16_2),
		.in_wire_3_3(vertical_tile_27_16_to_tile_28_16_3),
		.out_wire_1_0(vertical_tile_28_16_to_tile_29_16_0),
		.out_wire_1_1(vertical_tile_28_16_to_tile_29_16_1),
		.out_wire_1_2(vertical_tile_28_16_to_tile_29_16_2),
		.out_wire_1_3(vertical_tile_28_16_to_tile_29_16_3),
		.in_wire_1_0(vertical_tile_29_16_to_tile_28_16_0),
		.in_wire_1_1(vertical_tile_29_16_to_tile_28_16_1),
		.in_wire_1_2(vertical_tile_29_16_to_tile_28_16_2),
		.in_wire_1_3(vertical_tile_29_16_to_tile_28_16_3),
		.out_wire_2_0(horizontal_tile_28_16_to_tile_28_15_0),
		.out_wire_2_1(horizontal_tile_28_16_to_tile_28_15_1),
		.out_wire_2_2(horizontal_tile_28_16_to_tile_28_15_2),
		.out_wire_2_3(horizontal_tile_28_16_to_tile_28_15_3),
		.in_wire_2_0(horizontal_tile_28_15_to_tile_28_16_0),
		.in_wire_2_1(horizontal_tile_28_15_to_tile_28_16_1),
		.in_wire_2_2(horizontal_tile_28_15_to_tile_28_16_2),
		.in_wire_2_3(horizontal_tile_28_15_to_tile_28_16_3),
		.out_wire_0_0(horizontal_tile_28_16_to_tile_28_17_0),
		.out_wire_0_1(horizontal_tile_28_16_to_tile_28_17_1),
		.out_wire_0_2(horizontal_tile_28_16_to_tile_28_17_2),
		.out_wire_0_3(horizontal_tile_28_16_to_tile_28_17_3),
		.in_wire_0_0(horizontal_tile_28_17_to_tile_28_16_0),
		.in_wire_0_1(horizontal_tile_28_17_to_tile_28_16_1),
		.in_wire_0_2(horizontal_tile_28_17_to_tile_28_16_2),
		.in_wire_0_3(horizontal_tile_28_17_to_tile_28_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(913)
	);

	pe_tile pe_tile_28_17(
		.out_wire_3_0(vertical_tile_28_17_to_tile_27_17_0),
		.out_wire_3_1(vertical_tile_28_17_to_tile_27_17_1),
		.out_wire_3_2(vertical_tile_28_17_to_tile_27_17_2),
		.out_wire_3_3(vertical_tile_28_17_to_tile_27_17_3),
		.in_wire_3_0(vertical_tile_27_17_to_tile_28_17_0),
		.in_wire_3_1(vertical_tile_27_17_to_tile_28_17_1),
		.in_wire_3_2(vertical_tile_27_17_to_tile_28_17_2),
		.in_wire_3_3(vertical_tile_27_17_to_tile_28_17_3),
		.out_wire_1_0(vertical_tile_28_17_to_tile_29_17_0),
		.out_wire_1_1(vertical_tile_28_17_to_tile_29_17_1),
		.out_wire_1_2(vertical_tile_28_17_to_tile_29_17_2),
		.out_wire_1_3(vertical_tile_28_17_to_tile_29_17_3),
		.in_wire_1_0(vertical_tile_29_17_to_tile_28_17_0),
		.in_wire_1_1(vertical_tile_29_17_to_tile_28_17_1),
		.in_wire_1_2(vertical_tile_29_17_to_tile_28_17_2),
		.in_wire_1_3(vertical_tile_29_17_to_tile_28_17_3),
		.out_wire_2_0(horizontal_tile_28_17_to_tile_28_16_0),
		.out_wire_2_1(horizontal_tile_28_17_to_tile_28_16_1),
		.out_wire_2_2(horizontal_tile_28_17_to_tile_28_16_2),
		.out_wire_2_3(horizontal_tile_28_17_to_tile_28_16_3),
		.in_wire_2_0(horizontal_tile_28_16_to_tile_28_17_0),
		.in_wire_2_1(horizontal_tile_28_16_to_tile_28_17_1),
		.in_wire_2_2(horizontal_tile_28_16_to_tile_28_17_2),
		.in_wire_2_3(horizontal_tile_28_16_to_tile_28_17_3),
		.out_wire_0_0(horizontal_tile_28_17_to_tile_28_18_0),
		.out_wire_0_1(horizontal_tile_28_17_to_tile_28_18_1),
		.out_wire_0_2(horizontal_tile_28_17_to_tile_28_18_2),
		.out_wire_0_3(horizontal_tile_28_17_to_tile_28_18_3),
		.in_wire_0_0(horizontal_tile_28_18_to_tile_28_17_0),
		.in_wire_0_1(horizontal_tile_28_18_to_tile_28_17_1),
		.in_wire_0_2(horizontal_tile_28_18_to_tile_28_17_2),
		.in_wire_0_3(horizontal_tile_28_18_to_tile_28_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(914)
	);

	pe_tile pe_tile_28_18(
		.out_wire_3_0(vertical_tile_28_18_to_tile_27_18_0),
		.out_wire_3_1(vertical_tile_28_18_to_tile_27_18_1),
		.out_wire_3_2(vertical_tile_28_18_to_tile_27_18_2),
		.out_wire_3_3(vertical_tile_28_18_to_tile_27_18_3),
		.in_wire_3_0(vertical_tile_27_18_to_tile_28_18_0),
		.in_wire_3_1(vertical_tile_27_18_to_tile_28_18_1),
		.in_wire_3_2(vertical_tile_27_18_to_tile_28_18_2),
		.in_wire_3_3(vertical_tile_27_18_to_tile_28_18_3),
		.out_wire_1_0(vertical_tile_28_18_to_tile_29_18_0),
		.out_wire_1_1(vertical_tile_28_18_to_tile_29_18_1),
		.out_wire_1_2(vertical_tile_28_18_to_tile_29_18_2),
		.out_wire_1_3(vertical_tile_28_18_to_tile_29_18_3),
		.in_wire_1_0(vertical_tile_29_18_to_tile_28_18_0),
		.in_wire_1_1(vertical_tile_29_18_to_tile_28_18_1),
		.in_wire_1_2(vertical_tile_29_18_to_tile_28_18_2),
		.in_wire_1_3(vertical_tile_29_18_to_tile_28_18_3),
		.out_wire_2_0(horizontal_tile_28_18_to_tile_28_17_0),
		.out_wire_2_1(horizontal_tile_28_18_to_tile_28_17_1),
		.out_wire_2_2(horizontal_tile_28_18_to_tile_28_17_2),
		.out_wire_2_3(horizontal_tile_28_18_to_tile_28_17_3),
		.in_wire_2_0(horizontal_tile_28_17_to_tile_28_18_0),
		.in_wire_2_1(horizontal_tile_28_17_to_tile_28_18_1),
		.in_wire_2_2(horizontal_tile_28_17_to_tile_28_18_2),
		.in_wire_2_3(horizontal_tile_28_17_to_tile_28_18_3),
		.out_wire_0_0(horizontal_tile_28_18_to_tile_28_19_0),
		.out_wire_0_1(horizontal_tile_28_18_to_tile_28_19_1),
		.out_wire_0_2(horizontal_tile_28_18_to_tile_28_19_2),
		.out_wire_0_3(horizontal_tile_28_18_to_tile_28_19_3),
		.in_wire_0_0(horizontal_tile_28_19_to_tile_28_18_0),
		.in_wire_0_1(horizontal_tile_28_19_to_tile_28_18_1),
		.in_wire_0_2(horizontal_tile_28_19_to_tile_28_18_2),
		.in_wire_0_3(horizontal_tile_28_19_to_tile_28_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(915)
	);

	pe_tile pe_tile_28_19(
		.out_wire_3_0(vertical_tile_28_19_to_tile_27_19_0),
		.out_wire_3_1(vertical_tile_28_19_to_tile_27_19_1),
		.out_wire_3_2(vertical_tile_28_19_to_tile_27_19_2),
		.out_wire_3_3(vertical_tile_28_19_to_tile_27_19_3),
		.in_wire_3_0(vertical_tile_27_19_to_tile_28_19_0),
		.in_wire_3_1(vertical_tile_27_19_to_tile_28_19_1),
		.in_wire_3_2(vertical_tile_27_19_to_tile_28_19_2),
		.in_wire_3_3(vertical_tile_27_19_to_tile_28_19_3),
		.out_wire_1_0(vertical_tile_28_19_to_tile_29_19_0),
		.out_wire_1_1(vertical_tile_28_19_to_tile_29_19_1),
		.out_wire_1_2(vertical_tile_28_19_to_tile_29_19_2),
		.out_wire_1_3(vertical_tile_28_19_to_tile_29_19_3),
		.in_wire_1_0(vertical_tile_29_19_to_tile_28_19_0),
		.in_wire_1_1(vertical_tile_29_19_to_tile_28_19_1),
		.in_wire_1_2(vertical_tile_29_19_to_tile_28_19_2),
		.in_wire_1_3(vertical_tile_29_19_to_tile_28_19_3),
		.out_wire_2_0(horizontal_tile_28_19_to_tile_28_18_0),
		.out_wire_2_1(horizontal_tile_28_19_to_tile_28_18_1),
		.out_wire_2_2(horizontal_tile_28_19_to_tile_28_18_2),
		.out_wire_2_3(horizontal_tile_28_19_to_tile_28_18_3),
		.in_wire_2_0(horizontal_tile_28_18_to_tile_28_19_0),
		.in_wire_2_1(horizontal_tile_28_18_to_tile_28_19_1),
		.in_wire_2_2(horizontal_tile_28_18_to_tile_28_19_2),
		.in_wire_2_3(horizontal_tile_28_18_to_tile_28_19_3),
		.out_wire_0_0(horizontal_tile_28_19_to_tile_28_20_0),
		.out_wire_0_1(horizontal_tile_28_19_to_tile_28_20_1),
		.out_wire_0_2(horizontal_tile_28_19_to_tile_28_20_2),
		.out_wire_0_3(horizontal_tile_28_19_to_tile_28_20_3),
		.in_wire_0_0(horizontal_tile_28_20_to_tile_28_19_0),
		.in_wire_0_1(horizontal_tile_28_20_to_tile_28_19_1),
		.in_wire_0_2(horizontal_tile_28_20_to_tile_28_19_2),
		.in_wire_0_3(horizontal_tile_28_20_to_tile_28_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(916)
	);

	pe_tile pe_tile_28_20(
		.out_wire_3_0(vertical_tile_28_20_to_tile_27_20_0),
		.out_wire_3_1(vertical_tile_28_20_to_tile_27_20_1),
		.out_wire_3_2(vertical_tile_28_20_to_tile_27_20_2),
		.out_wire_3_3(vertical_tile_28_20_to_tile_27_20_3),
		.in_wire_3_0(vertical_tile_27_20_to_tile_28_20_0),
		.in_wire_3_1(vertical_tile_27_20_to_tile_28_20_1),
		.in_wire_3_2(vertical_tile_27_20_to_tile_28_20_2),
		.in_wire_3_3(vertical_tile_27_20_to_tile_28_20_3),
		.out_wire_1_0(vertical_tile_28_20_to_tile_29_20_0),
		.out_wire_1_1(vertical_tile_28_20_to_tile_29_20_1),
		.out_wire_1_2(vertical_tile_28_20_to_tile_29_20_2),
		.out_wire_1_3(vertical_tile_28_20_to_tile_29_20_3),
		.in_wire_1_0(vertical_tile_29_20_to_tile_28_20_0),
		.in_wire_1_1(vertical_tile_29_20_to_tile_28_20_1),
		.in_wire_1_2(vertical_tile_29_20_to_tile_28_20_2),
		.in_wire_1_3(vertical_tile_29_20_to_tile_28_20_3),
		.out_wire_2_0(horizontal_tile_28_20_to_tile_28_19_0),
		.out_wire_2_1(horizontal_tile_28_20_to_tile_28_19_1),
		.out_wire_2_2(horizontal_tile_28_20_to_tile_28_19_2),
		.out_wire_2_3(horizontal_tile_28_20_to_tile_28_19_3),
		.in_wire_2_0(horizontal_tile_28_19_to_tile_28_20_0),
		.in_wire_2_1(horizontal_tile_28_19_to_tile_28_20_1),
		.in_wire_2_2(horizontal_tile_28_19_to_tile_28_20_2),
		.in_wire_2_3(horizontal_tile_28_19_to_tile_28_20_3),
		.out_wire_0_0(horizontal_tile_28_20_to_tile_28_21_0),
		.out_wire_0_1(horizontal_tile_28_20_to_tile_28_21_1),
		.out_wire_0_2(horizontal_tile_28_20_to_tile_28_21_2),
		.out_wire_0_3(horizontal_tile_28_20_to_tile_28_21_3),
		.in_wire_0_0(horizontal_tile_28_21_to_tile_28_20_0),
		.in_wire_0_1(horizontal_tile_28_21_to_tile_28_20_1),
		.in_wire_0_2(horizontal_tile_28_21_to_tile_28_20_2),
		.in_wire_0_3(horizontal_tile_28_21_to_tile_28_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(917)
	);

	pe_tile pe_tile_28_21(
		.out_wire_3_0(vertical_tile_28_21_to_tile_27_21_0),
		.out_wire_3_1(vertical_tile_28_21_to_tile_27_21_1),
		.out_wire_3_2(vertical_tile_28_21_to_tile_27_21_2),
		.out_wire_3_3(vertical_tile_28_21_to_tile_27_21_3),
		.in_wire_3_0(vertical_tile_27_21_to_tile_28_21_0),
		.in_wire_3_1(vertical_tile_27_21_to_tile_28_21_1),
		.in_wire_3_2(vertical_tile_27_21_to_tile_28_21_2),
		.in_wire_3_3(vertical_tile_27_21_to_tile_28_21_3),
		.out_wire_1_0(vertical_tile_28_21_to_tile_29_21_0),
		.out_wire_1_1(vertical_tile_28_21_to_tile_29_21_1),
		.out_wire_1_2(vertical_tile_28_21_to_tile_29_21_2),
		.out_wire_1_3(vertical_tile_28_21_to_tile_29_21_3),
		.in_wire_1_0(vertical_tile_29_21_to_tile_28_21_0),
		.in_wire_1_1(vertical_tile_29_21_to_tile_28_21_1),
		.in_wire_1_2(vertical_tile_29_21_to_tile_28_21_2),
		.in_wire_1_3(vertical_tile_29_21_to_tile_28_21_3),
		.out_wire_2_0(horizontal_tile_28_21_to_tile_28_20_0),
		.out_wire_2_1(horizontal_tile_28_21_to_tile_28_20_1),
		.out_wire_2_2(horizontal_tile_28_21_to_tile_28_20_2),
		.out_wire_2_3(horizontal_tile_28_21_to_tile_28_20_3),
		.in_wire_2_0(horizontal_tile_28_20_to_tile_28_21_0),
		.in_wire_2_1(horizontal_tile_28_20_to_tile_28_21_1),
		.in_wire_2_2(horizontal_tile_28_20_to_tile_28_21_2),
		.in_wire_2_3(horizontal_tile_28_20_to_tile_28_21_3),
		.out_wire_0_0(horizontal_tile_28_21_to_tile_28_22_0),
		.out_wire_0_1(horizontal_tile_28_21_to_tile_28_22_1),
		.out_wire_0_2(horizontal_tile_28_21_to_tile_28_22_2),
		.out_wire_0_3(horizontal_tile_28_21_to_tile_28_22_3),
		.in_wire_0_0(horizontal_tile_28_22_to_tile_28_21_0),
		.in_wire_0_1(horizontal_tile_28_22_to_tile_28_21_1),
		.in_wire_0_2(horizontal_tile_28_22_to_tile_28_21_2),
		.in_wire_0_3(horizontal_tile_28_22_to_tile_28_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(918)
	);

	pe_tile pe_tile_28_22(
		.out_wire_3_0(vertical_tile_28_22_to_tile_27_22_0),
		.out_wire_3_1(vertical_tile_28_22_to_tile_27_22_1),
		.out_wire_3_2(vertical_tile_28_22_to_tile_27_22_2),
		.out_wire_3_3(vertical_tile_28_22_to_tile_27_22_3),
		.in_wire_3_0(vertical_tile_27_22_to_tile_28_22_0),
		.in_wire_3_1(vertical_tile_27_22_to_tile_28_22_1),
		.in_wire_3_2(vertical_tile_27_22_to_tile_28_22_2),
		.in_wire_3_3(vertical_tile_27_22_to_tile_28_22_3),
		.out_wire_1_0(vertical_tile_28_22_to_tile_29_22_0),
		.out_wire_1_1(vertical_tile_28_22_to_tile_29_22_1),
		.out_wire_1_2(vertical_tile_28_22_to_tile_29_22_2),
		.out_wire_1_3(vertical_tile_28_22_to_tile_29_22_3),
		.in_wire_1_0(vertical_tile_29_22_to_tile_28_22_0),
		.in_wire_1_1(vertical_tile_29_22_to_tile_28_22_1),
		.in_wire_1_2(vertical_tile_29_22_to_tile_28_22_2),
		.in_wire_1_3(vertical_tile_29_22_to_tile_28_22_3),
		.out_wire_2_0(horizontal_tile_28_22_to_tile_28_21_0),
		.out_wire_2_1(horizontal_tile_28_22_to_tile_28_21_1),
		.out_wire_2_2(horizontal_tile_28_22_to_tile_28_21_2),
		.out_wire_2_3(horizontal_tile_28_22_to_tile_28_21_3),
		.in_wire_2_0(horizontal_tile_28_21_to_tile_28_22_0),
		.in_wire_2_1(horizontal_tile_28_21_to_tile_28_22_1),
		.in_wire_2_2(horizontal_tile_28_21_to_tile_28_22_2),
		.in_wire_2_3(horizontal_tile_28_21_to_tile_28_22_3),
		.out_wire_0_0(horizontal_tile_28_22_to_tile_28_23_0),
		.out_wire_0_1(horizontal_tile_28_22_to_tile_28_23_1),
		.out_wire_0_2(horizontal_tile_28_22_to_tile_28_23_2),
		.out_wire_0_3(horizontal_tile_28_22_to_tile_28_23_3),
		.in_wire_0_0(horizontal_tile_28_23_to_tile_28_22_0),
		.in_wire_0_1(horizontal_tile_28_23_to_tile_28_22_1),
		.in_wire_0_2(horizontal_tile_28_23_to_tile_28_22_2),
		.in_wire_0_3(horizontal_tile_28_23_to_tile_28_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(919)
	);

	pe_tile pe_tile_28_23(
		.out_wire_3_0(vertical_tile_28_23_to_tile_27_23_0),
		.out_wire_3_1(vertical_tile_28_23_to_tile_27_23_1),
		.out_wire_3_2(vertical_tile_28_23_to_tile_27_23_2),
		.out_wire_3_3(vertical_tile_28_23_to_tile_27_23_3),
		.in_wire_3_0(vertical_tile_27_23_to_tile_28_23_0),
		.in_wire_3_1(vertical_tile_27_23_to_tile_28_23_1),
		.in_wire_3_2(vertical_tile_27_23_to_tile_28_23_2),
		.in_wire_3_3(vertical_tile_27_23_to_tile_28_23_3),
		.out_wire_1_0(vertical_tile_28_23_to_tile_29_23_0),
		.out_wire_1_1(vertical_tile_28_23_to_tile_29_23_1),
		.out_wire_1_2(vertical_tile_28_23_to_tile_29_23_2),
		.out_wire_1_3(vertical_tile_28_23_to_tile_29_23_3),
		.in_wire_1_0(vertical_tile_29_23_to_tile_28_23_0),
		.in_wire_1_1(vertical_tile_29_23_to_tile_28_23_1),
		.in_wire_1_2(vertical_tile_29_23_to_tile_28_23_2),
		.in_wire_1_3(vertical_tile_29_23_to_tile_28_23_3),
		.out_wire_2_0(horizontal_tile_28_23_to_tile_28_22_0),
		.out_wire_2_1(horizontal_tile_28_23_to_tile_28_22_1),
		.out_wire_2_2(horizontal_tile_28_23_to_tile_28_22_2),
		.out_wire_2_3(horizontal_tile_28_23_to_tile_28_22_3),
		.in_wire_2_0(horizontal_tile_28_22_to_tile_28_23_0),
		.in_wire_2_1(horizontal_tile_28_22_to_tile_28_23_1),
		.in_wire_2_2(horizontal_tile_28_22_to_tile_28_23_2),
		.in_wire_2_3(horizontal_tile_28_22_to_tile_28_23_3),
		.out_wire_0_0(horizontal_tile_28_23_to_tile_28_24_0),
		.out_wire_0_1(horizontal_tile_28_23_to_tile_28_24_1),
		.out_wire_0_2(horizontal_tile_28_23_to_tile_28_24_2),
		.out_wire_0_3(horizontal_tile_28_23_to_tile_28_24_3),
		.in_wire_0_0(horizontal_tile_28_24_to_tile_28_23_0),
		.in_wire_0_1(horizontal_tile_28_24_to_tile_28_23_1),
		.in_wire_0_2(horizontal_tile_28_24_to_tile_28_23_2),
		.in_wire_0_3(horizontal_tile_28_24_to_tile_28_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(920)
	);

	pe_tile pe_tile_28_24(
		.out_wire_3_0(vertical_tile_28_24_to_tile_27_24_0),
		.out_wire_3_1(vertical_tile_28_24_to_tile_27_24_1),
		.out_wire_3_2(vertical_tile_28_24_to_tile_27_24_2),
		.out_wire_3_3(vertical_tile_28_24_to_tile_27_24_3),
		.in_wire_3_0(vertical_tile_27_24_to_tile_28_24_0),
		.in_wire_3_1(vertical_tile_27_24_to_tile_28_24_1),
		.in_wire_3_2(vertical_tile_27_24_to_tile_28_24_2),
		.in_wire_3_3(vertical_tile_27_24_to_tile_28_24_3),
		.out_wire_1_0(vertical_tile_28_24_to_tile_29_24_0),
		.out_wire_1_1(vertical_tile_28_24_to_tile_29_24_1),
		.out_wire_1_2(vertical_tile_28_24_to_tile_29_24_2),
		.out_wire_1_3(vertical_tile_28_24_to_tile_29_24_3),
		.in_wire_1_0(vertical_tile_29_24_to_tile_28_24_0),
		.in_wire_1_1(vertical_tile_29_24_to_tile_28_24_1),
		.in_wire_1_2(vertical_tile_29_24_to_tile_28_24_2),
		.in_wire_1_3(vertical_tile_29_24_to_tile_28_24_3),
		.out_wire_2_0(horizontal_tile_28_24_to_tile_28_23_0),
		.out_wire_2_1(horizontal_tile_28_24_to_tile_28_23_1),
		.out_wire_2_2(horizontal_tile_28_24_to_tile_28_23_2),
		.out_wire_2_3(horizontal_tile_28_24_to_tile_28_23_3),
		.in_wire_2_0(horizontal_tile_28_23_to_tile_28_24_0),
		.in_wire_2_1(horizontal_tile_28_23_to_tile_28_24_1),
		.in_wire_2_2(horizontal_tile_28_23_to_tile_28_24_2),
		.in_wire_2_3(horizontal_tile_28_23_to_tile_28_24_3),
		.out_wire_0_0(horizontal_tile_28_24_to_tile_28_25_0),
		.out_wire_0_1(horizontal_tile_28_24_to_tile_28_25_1),
		.out_wire_0_2(horizontal_tile_28_24_to_tile_28_25_2),
		.out_wire_0_3(horizontal_tile_28_24_to_tile_28_25_3),
		.in_wire_0_0(horizontal_tile_28_25_to_tile_28_24_0),
		.in_wire_0_1(horizontal_tile_28_25_to_tile_28_24_1),
		.in_wire_0_2(horizontal_tile_28_25_to_tile_28_24_2),
		.in_wire_0_3(horizontal_tile_28_25_to_tile_28_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(921)
	);

	pe_tile pe_tile_28_25(
		.out_wire_3_0(vertical_tile_28_25_to_tile_27_25_0),
		.out_wire_3_1(vertical_tile_28_25_to_tile_27_25_1),
		.out_wire_3_2(vertical_tile_28_25_to_tile_27_25_2),
		.out_wire_3_3(vertical_tile_28_25_to_tile_27_25_3),
		.in_wire_3_0(vertical_tile_27_25_to_tile_28_25_0),
		.in_wire_3_1(vertical_tile_27_25_to_tile_28_25_1),
		.in_wire_3_2(vertical_tile_27_25_to_tile_28_25_2),
		.in_wire_3_3(vertical_tile_27_25_to_tile_28_25_3),
		.out_wire_1_0(vertical_tile_28_25_to_tile_29_25_0),
		.out_wire_1_1(vertical_tile_28_25_to_tile_29_25_1),
		.out_wire_1_2(vertical_tile_28_25_to_tile_29_25_2),
		.out_wire_1_3(vertical_tile_28_25_to_tile_29_25_3),
		.in_wire_1_0(vertical_tile_29_25_to_tile_28_25_0),
		.in_wire_1_1(vertical_tile_29_25_to_tile_28_25_1),
		.in_wire_1_2(vertical_tile_29_25_to_tile_28_25_2),
		.in_wire_1_3(vertical_tile_29_25_to_tile_28_25_3),
		.out_wire_2_0(horizontal_tile_28_25_to_tile_28_24_0),
		.out_wire_2_1(horizontal_tile_28_25_to_tile_28_24_1),
		.out_wire_2_2(horizontal_tile_28_25_to_tile_28_24_2),
		.out_wire_2_3(horizontal_tile_28_25_to_tile_28_24_3),
		.in_wire_2_0(horizontal_tile_28_24_to_tile_28_25_0),
		.in_wire_2_1(horizontal_tile_28_24_to_tile_28_25_1),
		.in_wire_2_2(horizontal_tile_28_24_to_tile_28_25_2),
		.in_wire_2_3(horizontal_tile_28_24_to_tile_28_25_3),
		.out_wire_0_0(horizontal_tile_28_25_to_tile_28_26_0),
		.out_wire_0_1(horizontal_tile_28_25_to_tile_28_26_1),
		.out_wire_0_2(horizontal_tile_28_25_to_tile_28_26_2),
		.out_wire_0_3(horizontal_tile_28_25_to_tile_28_26_3),
		.in_wire_0_0(horizontal_tile_28_26_to_tile_28_25_0),
		.in_wire_0_1(horizontal_tile_28_26_to_tile_28_25_1),
		.in_wire_0_2(horizontal_tile_28_26_to_tile_28_25_2),
		.in_wire_0_3(horizontal_tile_28_26_to_tile_28_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(922)
	);

	pe_tile pe_tile_28_26(
		.out_wire_3_0(vertical_tile_28_26_to_tile_27_26_0),
		.out_wire_3_1(vertical_tile_28_26_to_tile_27_26_1),
		.out_wire_3_2(vertical_tile_28_26_to_tile_27_26_2),
		.out_wire_3_3(vertical_tile_28_26_to_tile_27_26_3),
		.in_wire_3_0(vertical_tile_27_26_to_tile_28_26_0),
		.in_wire_3_1(vertical_tile_27_26_to_tile_28_26_1),
		.in_wire_3_2(vertical_tile_27_26_to_tile_28_26_2),
		.in_wire_3_3(vertical_tile_27_26_to_tile_28_26_3),
		.out_wire_1_0(vertical_tile_28_26_to_tile_29_26_0),
		.out_wire_1_1(vertical_tile_28_26_to_tile_29_26_1),
		.out_wire_1_2(vertical_tile_28_26_to_tile_29_26_2),
		.out_wire_1_3(vertical_tile_28_26_to_tile_29_26_3),
		.in_wire_1_0(vertical_tile_29_26_to_tile_28_26_0),
		.in_wire_1_1(vertical_tile_29_26_to_tile_28_26_1),
		.in_wire_1_2(vertical_tile_29_26_to_tile_28_26_2),
		.in_wire_1_3(vertical_tile_29_26_to_tile_28_26_3),
		.out_wire_2_0(horizontal_tile_28_26_to_tile_28_25_0),
		.out_wire_2_1(horizontal_tile_28_26_to_tile_28_25_1),
		.out_wire_2_2(horizontal_tile_28_26_to_tile_28_25_2),
		.out_wire_2_3(horizontal_tile_28_26_to_tile_28_25_3),
		.in_wire_2_0(horizontal_tile_28_25_to_tile_28_26_0),
		.in_wire_2_1(horizontal_tile_28_25_to_tile_28_26_1),
		.in_wire_2_2(horizontal_tile_28_25_to_tile_28_26_2),
		.in_wire_2_3(horizontal_tile_28_25_to_tile_28_26_3),
		.out_wire_0_0(horizontal_tile_28_26_to_tile_28_27_0),
		.out_wire_0_1(horizontal_tile_28_26_to_tile_28_27_1),
		.out_wire_0_2(horizontal_tile_28_26_to_tile_28_27_2),
		.out_wire_0_3(horizontal_tile_28_26_to_tile_28_27_3),
		.in_wire_0_0(horizontal_tile_28_27_to_tile_28_26_0),
		.in_wire_0_1(horizontal_tile_28_27_to_tile_28_26_1),
		.in_wire_0_2(horizontal_tile_28_27_to_tile_28_26_2),
		.in_wire_0_3(horizontal_tile_28_27_to_tile_28_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(923)
	);

	pe_tile pe_tile_28_27(
		.out_wire_3_0(vertical_tile_28_27_to_tile_27_27_0),
		.out_wire_3_1(vertical_tile_28_27_to_tile_27_27_1),
		.out_wire_3_2(vertical_tile_28_27_to_tile_27_27_2),
		.out_wire_3_3(vertical_tile_28_27_to_tile_27_27_3),
		.in_wire_3_0(vertical_tile_27_27_to_tile_28_27_0),
		.in_wire_3_1(vertical_tile_27_27_to_tile_28_27_1),
		.in_wire_3_2(vertical_tile_27_27_to_tile_28_27_2),
		.in_wire_3_3(vertical_tile_27_27_to_tile_28_27_3),
		.out_wire_1_0(vertical_tile_28_27_to_tile_29_27_0),
		.out_wire_1_1(vertical_tile_28_27_to_tile_29_27_1),
		.out_wire_1_2(vertical_tile_28_27_to_tile_29_27_2),
		.out_wire_1_3(vertical_tile_28_27_to_tile_29_27_3),
		.in_wire_1_0(vertical_tile_29_27_to_tile_28_27_0),
		.in_wire_1_1(vertical_tile_29_27_to_tile_28_27_1),
		.in_wire_1_2(vertical_tile_29_27_to_tile_28_27_2),
		.in_wire_1_3(vertical_tile_29_27_to_tile_28_27_3),
		.out_wire_2_0(horizontal_tile_28_27_to_tile_28_26_0),
		.out_wire_2_1(horizontal_tile_28_27_to_tile_28_26_1),
		.out_wire_2_2(horizontal_tile_28_27_to_tile_28_26_2),
		.out_wire_2_3(horizontal_tile_28_27_to_tile_28_26_3),
		.in_wire_2_0(horizontal_tile_28_26_to_tile_28_27_0),
		.in_wire_2_1(horizontal_tile_28_26_to_tile_28_27_1),
		.in_wire_2_2(horizontal_tile_28_26_to_tile_28_27_2),
		.in_wire_2_3(horizontal_tile_28_26_to_tile_28_27_3),
		.out_wire_0_0(horizontal_tile_28_27_to_tile_28_28_0),
		.out_wire_0_1(horizontal_tile_28_27_to_tile_28_28_1),
		.out_wire_0_2(horizontal_tile_28_27_to_tile_28_28_2),
		.out_wire_0_3(horizontal_tile_28_27_to_tile_28_28_3),
		.in_wire_0_0(horizontal_tile_28_28_to_tile_28_27_0),
		.in_wire_0_1(horizontal_tile_28_28_to_tile_28_27_1),
		.in_wire_0_2(horizontal_tile_28_28_to_tile_28_27_2),
		.in_wire_0_3(horizontal_tile_28_28_to_tile_28_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(924)
	);

	pe_tile pe_tile_28_28(
		.out_wire_3_0(vertical_tile_28_28_to_tile_27_28_0),
		.out_wire_3_1(vertical_tile_28_28_to_tile_27_28_1),
		.out_wire_3_2(vertical_tile_28_28_to_tile_27_28_2),
		.out_wire_3_3(vertical_tile_28_28_to_tile_27_28_3),
		.in_wire_3_0(vertical_tile_27_28_to_tile_28_28_0),
		.in_wire_3_1(vertical_tile_27_28_to_tile_28_28_1),
		.in_wire_3_2(vertical_tile_27_28_to_tile_28_28_2),
		.in_wire_3_3(vertical_tile_27_28_to_tile_28_28_3),
		.out_wire_1_0(vertical_tile_28_28_to_tile_29_28_0),
		.out_wire_1_1(vertical_tile_28_28_to_tile_29_28_1),
		.out_wire_1_2(vertical_tile_28_28_to_tile_29_28_2),
		.out_wire_1_3(vertical_tile_28_28_to_tile_29_28_3),
		.in_wire_1_0(vertical_tile_29_28_to_tile_28_28_0),
		.in_wire_1_1(vertical_tile_29_28_to_tile_28_28_1),
		.in_wire_1_2(vertical_tile_29_28_to_tile_28_28_2),
		.in_wire_1_3(vertical_tile_29_28_to_tile_28_28_3),
		.out_wire_2_0(horizontal_tile_28_28_to_tile_28_27_0),
		.out_wire_2_1(horizontal_tile_28_28_to_tile_28_27_1),
		.out_wire_2_2(horizontal_tile_28_28_to_tile_28_27_2),
		.out_wire_2_3(horizontal_tile_28_28_to_tile_28_27_3),
		.in_wire_2_0(horizontal_tile_28_27_to_tile_28_28_0),
		.in_wire_2_1(horizontal_tile_28_27_to_tile_28_28_1),
		.in_wire_2_2(horizontal_tile_28_27_to_tile_28_28_2),
		.in_wire_2_3(horizontal_tile_28_27_to_tile_28_28_3),
		.out_wire_0_0(horizontal_tile_28_28_to_tile_28_29_0),
		.out_wire_0_1(horizontal_tile_28_28_to_tile_28_29_1),
		.out_wire_0_2(horizontal_tile_28_28_to_tile_28_29_2),
		.out_wire_0_3(horizontal_tile_28_28_to_tile_28_29_3),
		.in_wire_0_0(horizontal_tile_28_29_to_tile_28_28_0),
		.in_wire_0_1(horizontal_tile_28_29_to_tile_28_28_1),
		.in_wire_0_2(horizontal_tile_28_29_to_tile_28_28_2),
		.in_wire_0_3(horizontal_tile_28_29_to_tile_28_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(925)
	);

	pe_tile pe_tile_28_29(
		.out_wire_3_0(vertical_tile_28_29_to_tile_27_29_0),
		.out_wire_3_1(vertical_tile_28_29_to_tile_27_29_1),
		.out_wire_3_2(vertical_tile_28_29_to_tile_27_29_2),
		.out_wire_3_3(vertical_tile_28_29_to_tile_27_29_3),
		.in_wire_3_0(vertical_tile_27_29_to_tile_28_29_0),
		.in_wire_3_1(vertical_tile_27_29_to_tile_28_29_1),
		.in_wire_3_2(vertical_tile_27_29_to_tile_28_29_2),
		.in_wire_3_3(vertical_tile_27_29_to_tile_28_29_3),
		.out_wire_1_0(vertical_tile_28_29_to_tile_29_29_0),
		.out_wire_1_1(vertical_tile_28_29_to_tile_29_29_1),
		.out_wire_1_2(vertical_tile_28_29_to_tile_29_29_2),
		.out_wire_1_3(vertical_tile_28_29_to_tile_29_29_3),
		.in_wire_1_0(vertical_tile_29_29_to_tile_28_29_0),
		.in_wire_1_1(vertical_tile_29_29_to_tile_28_29_1),
		.in_wire_1_2(vertical_tile_29_29_to_tile_28_29_2),
		.in_wire_1_3(vertical_tile_29_29_to_tile_28_29_3),
		.out_wire_2_0(horizontal_tile_28_29_to_tile_28_28_0),
		.out_wire_2_1(horizontal_tile_28_29_to_tile_28_28_1),
		.out_wire_2_2(horizontal_tile_28_29_to_tile_28_28_2),
		.out_wire_2_3(horizontal_tile_28_29_to_tile_28_28_3),
		.in_wire_2_0(horizontal_tile_28_28_to_tile_28_29_0),
		.in_wire_2_1(horizontal_tile_28_28_to_tile_28_29_1),
		.in_wire_2_2(horizontal_tile_28_28_to_tile_28_29_2),
		.in_wire_2_3(horizontal_tile_28_28_to_tile_28_29_3),
		.out_wire_0_0(horizontal_tile_28_29_to_tile_28_30_0),
		.out_wire_0_1(horizontal_tile_28_29_to_tile_28_30_1),
		.out_wire_0_2(horizontal_tile_28_29_to_tile_28_30_2),
		.out_wire_0_3(horizontal_tile_28_29_to_tile_28_30_3),
		.in_wire_0_0(horizontal_tile_28_30_to_tile_28_29_0),
		.in_wire_0_1(horizontal_tile_28_30_to_tile_28_29_1),
		.in_wire_0_2(horizontal_tile_28_30_to_tile_28_29_2),
		.in_wire_0_3(horizontal_tile_28_30_to_tile_28_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(926)
	);

	pe_tile pe_tile_28_30(
		.out_wire_3_0(vertical_tile_28_30_to_tile_27_30_0),
		.out_wire_3_1(vertical_tile_28_30_to_tile_27_30_1),
		.out_wire_3_2(vertical_tile_28_30_to_tile_27_30_2),
		.out_wire_3_3(vertical_tile_28_30_to_tile_27_30_3),
		.in_wire_3_0(vertical_tile_27_30_to_tile_28_30_0),
		.in_wire_3_1(vertical_tile_27_30_to_tile_28_30_1),
		.in_wire_3_2(vertical_tile_27_30_to_tile_28_30_2),
		.in_wire_3_3(vertical_tile_27_30_to_tile_28_30_3),
		.out_wire_1_0(vertical_tile_28_30_to_tile_29_30_0),
		.out_wire_1_1(vertical_tile_28_30_to_tile_29_30_1),
		.out_wire_1_2(vertical_tile_28_30_to_tile_29_30_2),
		.out_wire_1_3(vertical_tile_28_30_to_tile_29_30_3),
		.in_wire_1_0(vertical_tile_29_30_to_tile_28_30_0),
		.in_wire_1_1(vertical_tile_29_30_to_tile_28_30_1),
		.in_wire_1_2(vertical_tile_29_30_to_tile_28_30_2),
		.in_wire_1_3(vertical_tile_29_30_to_tile_28_30_3),
		.out_wire_2_0(horizontal_tile_28_30_to_tile_28_29_0),
		.out_wire_2_1(horizontal_tile_28_30_to_tile_28_29_1),
		.out_wire_2_2(horizontal_tile_28_30_to_tile_28_29_2),
		.out_wire_2_3(horizontal_tile_28_30_to_tile_28_29_3),
		.in_wire_2_0(horizontal_tile_28_29_to_tile_28_30_0),
		.in_wire_2_1(horizontal_tile_28_29_to_tile_28_30_1),
		.in_wire_2_2(horizontal_tile_28_29_to_tile_28_30_2),
		.in_wire_2_3(horizontal_tile_28_29_to_tile_28_30_3),
		.out_wire_0_0(horizontal_tile_28_30_to_tile_28_31_0),
		.out_wire_0_1(horizontal_tile_28_30_to_tile_28_31_1),
		.out_wire_0_2(horizontal_tile_28_30_to_tile_28_31_2),
		.out_wire_0_3(horizontal_tile_28_30_to_tile_28_31_3),
		.in_wire_0_0(horizontal_tile_28_31_to_tile_28_30_0),
		.in_wire_0_1(horizontal_tile_28_31_to_tile_28_30_1),
		.in_wire_0_2(horizontal_tile_28_31_to_tile_28_30_2),
		.in_wire_0_3(horizontal_tile_28_31_to_tile_28_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(927)
	);

	pe_tile_right pe_tile_28_31(
		.out_wire_3_0(vertical_tile_28_31_to_tile_27_31_0),
		.out_wire_3_1(vertical_tile_28_31_to_tile_27_31_1),
		.out_wire_3_2(vertical_tile_28_31_to_tile_27_31_2),
		.out_wire_3_3(vertical_tile_28_31_to_tile_27_31_3),
		.in_wire_3_0(vertical_tile_27_31_to_tile_28_31_0),
		.in_wire_3_1(vertical_tile_27_31_to_tile_28_31_1),
		.in_wire_3_2(vertical_tile_27_31_to_tile_28_31_2),
		.in_wire_3_3(vertical_tile_27_31_to_tile_28_31_3),
		.out_wire_1_0(vertical_tile_28_31_to_tile_29_31_0),
		.out_wire_1_1(vertical_tile_28_31_to_tile_29_31_1),
		.out_wire_1_2(vertical_tile_28_31_to_tile_29_31_2),
		.out_wire_1_3(vertical_tile_28_31_to_tile_29_31_3),
		.in_wire_1_0(vertical_tile_29_31_to_tile_28_31_0),
		.in_wire_1_1(vertical_tile_29_31_to_tile_28_31_1),
		.in_wire_1_2(vertical_tile_29_31_to_tile_28_31_2),
		.in_wire_1_3(vertical_tile_29_31_to_tile_28_31_3),
		.out_wire_2_0(horizontal_tile_28_31_to_tile_28_30_0),
		.out_wire_2_1(horizontal_tile_28_31_to_tile_28_30_1),
		.out_wire_2_2(horizontal_tile_28_31_to_tile_28_30_2),
		.out_wire_2_3(horizontal_tile_28_31_to_tile_28_30_3),
		.in_wire_2_0(horizontal_tile_28_30_to_tile_28_31_0),
		.in_wire_2_1(horizontal_tile_28_30_to_tile_28_31_1),
		.in_wire_2_2(horizontal_tile_28_30_to_tile_28_31_2),
		.in_wire_2_3(horizontal_tile_28_30_to_tile_28_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(928)
	);

	pe_tile_left pe_tile_29_0(
		.out_wire_3_0(vertical_tile_29_0_to_tile_28_0_0),
		.out_wire_3_1(vertical_tile_29_0_to_tile_28_0_1),
		.out_wire_3_2(vertical_tile_29_0_to_tile_28_0_2),
		.out_wire_3_3(vertical_tile_29_0_to_tile_28_0_3),
		.in_wire_3_0(vertical_tile_28_0_to_tile_29_0_0),
		.in_wire_3_1(vertical_tile_28_0_to_tile_29_0_1),
		.in_wire_3_2(vertical_tile_28_0_to_tile_29_0_2),
		.in_wire_3_3(vertical_tile_28_0_to_tile_29_0_3),
		.out_wire_1_0(vertical_tile_29_0_to_tile_30_0_0),
		.out_wire_1_1(vertical_tile_29_0_to_tile_30_0_1),
		.out_wire_1_2(vertical_tile_29_0_to_tile_30_0_2),
		.out_wire_1_3(vertical_tile_29_0_to_tile_30_0_3),
		.in_wire_1_0(vertical_tile_30_0_to_tile_29_0_0),
		.in_wire_1_1(vertical_tile_30_0_to_tile_29_0_1),
		.in_wire_1_2(vertical_tile_30_0_to_tile_29_0_2),
		.in_wire_1_3(vertical_tile_30_0_to_tile_29_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_29_0_to_tile_29_1_0),
		.out_wire_0_1(horizontal_tile_29_0_to_tile_29_1_1),
		.out_wire_0_2(horizontal_tile_29_0_to_tile_29_1_2),
		.out_wire_0_3(horizontal_tile_29_0_to_tile_29_1_3),
		.in_wire_0_0(horizontal_tile_29_1_to_tile_29_0_0),
		.in_wire_0_1(horizontal_tile_29_1_to_tile_29_0_1),
		.in_wire_0_2(horizontal_tile_29_1_to_tile_29_0_2),
		.in_wire_0_3(horizontal_tile_29_1_to_tile_29_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(929)
	);

	pe_tile pe_tile_29_1(
		.out_wire_3_0(vertical_tile_29_1_to_tile_28_1_0),
		.out_wire_3_1(vertical_tile_29_1_to_tile_28_1_1),
		.out_wire_3_2(vertical_tile_29_1_to_tile_28_1_2),
		.out_wire_3_3(vertical_tile_29_1_to_tile_28_1_3),
		.in_wire_3_0(vertical_tile_28_1_to_tile_29_1_0),
		.in_wire_3_1(vertical_tile_28_1_to_tile_29_1_1),
		.in_wire_3_2(vertical_tile_28_1_to_tile_29_1_2),
		.in_wire_3_3(vertical_tile_28_1_to_tile_29_1_3),
		.out_wire_1_0(vertical_tile_29_1_to_tile_30_1_0),
		.out_wire_1_1(vertical_tile_29_1_to_tile_30_1_1),
		.out_wire_1_2(vertical_tile_29_1_to_tile_30_1_2),
		.out_wire_1_3(vertical_tile_29_1_to_tile_30_1_3),
		.in_wire_1_0(vertical_tile_30_1_to_tile_29_1_0),
		.in_wire_1_1(vertical_tile_30_1_to_tile_29_1_1),
		.in_wire_1_2(vertical_tile_30_1_to_tile_29_1_2),
		.in_wire_1_3(vertical_tile_30_1_to_tile_29_1_3),
		.out_wire_2_0(horizontal_tile_29_1_to_tile_29_0_0),
		.out_wire_2_1(horizontal_tile_29_1_to_tile_29_0_1),
		.out_wire_2_2(horizontal_tile_29_1_to_tile_29_0_2),
		.out_wire_2_3(horizontal_tile_29_1_to_tile_29_0_3),
		.in_wire_2_0(horizontal_tile_29_0_to_tile_29_1_0),
		.in_wire_2_1(horizontal_tile_29_0_to_tile_29_1_1),
		.in_wire_2_2(horizontal_tile_29_0_to_tile_29_1_2),
		.in_wire_2_3(horizontal_tile_29_0_to_tile_29_1_3),
		.out_wire_0_0(horizontal_tile_29_1_to_tile_29_2_0),
		.out_wire_0_1(horizontal_tile_29_1_to_tile_29_2_1),
		.out_wire_0_2(horizontal_tile_29_1_to_tile_29_2_2),
		.out_wire_0_3(horizontal_tile_29_1_to_tile_29_2_3),
		.in_wire_0_0(horizontal_tile_29_2_to_tile_29_1_0),
		.in_wire_0_1(horizontal_tile_29_2_to_tile_29_1_1),
		.in_wire_0_2(horizontal_tile_29_2_to_tile_29_1_2),
		.in_wire_0_3(horizontal_tile_29_2_to_tile_29_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(930)
	);

	pe_tile pe_tile_29_2(
		.out_wire_3_0(vertical_tile_29_2_to_tile_28_2_0),
		.out_wire_3_1(vertical_tile_29_2_to_tile_28_2_1),
		.out_wire_3_2(vertical_tile_29_2_to_tile_28_2_2),
		.out_wire_3_3(vertical_tile_29_2_to_tile_28_2_3),
		.in_wire_3_0(vertical_tile_28_2_to_tile_29_2_0),
		.in_wire_3_1(vertical_tile_28_2_to_tile_29_2_1),
		.in_wire_3_2(vertical_tile_28_2_to_tile_29_2_2),
		.in_wire_3_3(vertical_tile_28_2_to_tile_29_2_3),
		.out_wire_1_0(vertical_tile_29_2_to_tile_30_2_0),
		.out_wire_1_1(vertical_tile_29_2_to_tile_30_2_1),
		.out_wire_1_2(vertical_tile_29_2_to_tile_30_2_2),
		.out_wire_1_3(vertical_tile_29_2_to_tile_30_2_3),
		.in_wire_1_0(vertical_tile_30_2_to_tile_29_2_0),
		.in_wire_1_1(vertical_tile_30_2_to_tile_29_2_1),
		.in_wire_1_2(vertical_tile_30_2_to_tile_29_2_2),
		.in_wire_1_3(vertical_tile_30_2_to_tile_29_2_3),
		.out_wire_2_0(horizontal_tile_29_2_to_tile_29_1_0),
		.out_wire_2_1(horizontal_tile_29_2_to_tile_29_1_1),
		.out_wire_2_2(horizontal_tile_29_2_to_tile_29_1_2),
		.out_wire_2_3(horizontal_tile_29_2_to_tile_29_1_3),
		.in_wire_2_0(horizontal_tile_29_1_to_tile_29_2_0),
		.in_wire_2_1(horizontal_tile_29_1_to_tile_29_2_1),
		.in_wire_2_2(horizontal_tile_29_1_to_tile_29_2_2),
		.in_wire_2_3(horizontal_tile_29_1_to_tile_29_2_3),
		.out_wire_0_0(horizontal_tile_29_2_to_tile_29_3_0),
		.out_wire_0_1(horizontal_tile_29_2_to_tile_29_3_1),
		.out_wire_0_2(horizontal_tile_29_2_to_tile_29_3_2),
		.out_wire_0_3(horizontal_tile_29_2_to_tile_29_3_3),
		.in_wire_0_0(horizontal_tile_29_3_to_tile_29_2_0),
		.in_wire_0_1(horizontal_tile_29_3_to_tile_29_2_1),
		.in_wire_0_2(horizontal_tile_29_3_to_tile_29_2_2),
		.in_wire_0_3(horizontal_tile_29_3_to_tile_29_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(931)
	);

	pe_tile pe_tile_29_3(
		.out_wire_3_0(vertical_tile_29_3_to_tile_28_3_0),
		.out_wire_3_1(vertical_tile_29_3_to_tile_28_3_1),
		.out_wire_3_2(vertical_tile_29_3_to_tile_28_3_2),
		.out_wire_3_3(vertical_tile_29_3_to_tile_28_3_3),
		.in_wire_3_0(vertical_tile_28_3_to_tile_29_3_0),
		.in_wire_3_1(vertical_tile_28_3_to_tile_29_3_1),
		.in_wire_3_2(vertical_tile_28_3_to_tile_29_3_2),
		.in_wire_3_3(vertical_tile_28_3_to_tile_29_3_3),
		.out_wire_1_0(vertical_tile_29_3_to_tile_30_3_0),
		.out_wire_1_1(vertical_tile_29_3_to_tile_30_3_1),
		.out_wire_1_2(vertical_tile_29_3_to_tile_30_3_2),
		.out_wire_1_3(vertical_tile_29_3_to_tile_30_3_3),
		.in_wire_1_0(vertical_tile_30_3_to_tile_29_3_0),
		.in_wire_1_1(vertical_tile_30_3_to_tile_29_3_1),
		.in_wire_1_2(vertical_tile_30_3_to_tile_29_3_2),
		.in_wire_1_3(vertical_tile_30_3_to_tile_29_3_3),
		.out_wire_2_0(horizontal_tile_29_3_to_tile_29_2_0),
		.out_wire_2_1(horizontal_tile_29_3_to_tile_29_2_1),
		.out_wire_2_2(horizontal_tile_29_3_to_tile_29_2_2),
		.out_wire_2_3(horizontal_tile_29_3_to_tile_29_2_3),
		.in_wire_2_0(horizontal_tile_29_2_to_tile_29_3_0),
		.in_wire_2_1(horizontal_tile_29_2_to_tile_29_3_1),
		.in_wire_2_2(horizontal_tile_29_2_to_tile_29_3_2),
		.in_wire_2_3(horizontal_tile_29_2_to_tile_29_3_3),
		.out_wire_0_0(horizontal_tile_29_3_to_tile_29_4_0),
		.out_wire_0_1(horizontal_tile_29_3_to_tile_29_4_1),
		.out_wire_0_2(horizontal_tile_29_3_to_tile_29_4_2),
		.out_wire_0_3(horizontal_tile_29_3_to_tile_29_4_3),
		.in_wire_0_0(horizontal_tile_29_4_to_tile_29_3_0),
		.in_wire_0_1(horizontal_tile_29_4_to_tile_29_3_1),
		.in_wire_0_2(horizontal_tile_29_4_to_tile_29_3_2),
		.in_wire_0_3(horizontal_tile_29_4_to_tile_29_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(932)
	);

	pe_tile pe_tile_29_4(
		.out_wire_3_0(vertical_tile_29_4_to_tile_28_4_0),
		.out_wire_3_1(vertical_tile_29_4_to_tile_28_4_1),
		.out_wire_3_2(vertical_tile_29_4_to_tile_28_4_2),
		.out_wire_3_3(vertical_tile_29_4_to_tile_28_4_3),
		.in_wire_3_0(vertical_tile_28_4_to_tile_29_4_0),
		.in_wire_3_1(vertical_tile_28_4_to_tile_29_4_1),
		.in_wire_3_2(vertical_tile_28_4_to_tile_29_4_2),
		.in_wire_3_3(vertical_tile_28_4_to_tile_29_4_3),
		.out_wire_1_0(vertical_tile_29_4_to_tile_30_4_0),
		.out_wire_1_1(vertical_tile_29_4_to_tile_30_4_1),
		.out_wire_1_2(vertical_tile_29_4_to_tile_30_4_2),
		.out_wire_1_3(vertical_tile_29_4_to_tile_30_4_3),
		.in_wire_1_0(vertical_tile_30_4_to_tile_29_4_0),
		.in_wire_1_1(vertical_tile_30_4_to_tile_29_4_1),
		.in_wire_1_2(vertical_tile_30_4_to_tile_29_4_2),
		.in_wire_1_3(vertical_tile_30_4_to_tile_29_4_3),
		.out_wire_2_0(horizontal_tile_29_4_to_tile_29_3_0),
		.out_wire_2_1(horizontal_tile_29_4_to_tile_29_3_1),
		.out_wire_2_2(horizontal_tile_29_4_to_tile_29_3_2),
		.out_wire_2_3(horizontal_tile_29_4_to_tile_29_3_3),
		.in_wire_2_0(horizontal_tile_29_3_to_tile_29_4_0),
		.in_wire_2_1(horizontal_tile_29_3_to_tile_29_4_1),
		.in_wire_2_2(horizontal_tile_29_3_to_tile_29_4_2),
		.in_wire_2_3(horizontal_tile_29_3_to_tile_29_4_3),
		.out_wire_0_0(horizontal_tile_29_4_to_tile_29_5_0),
		.out_wire_0_1(horizontal_tile_29_4_to_tile_29_5_1),
		.out_wire_0_2(horizontal_tile_29_4_to_tile_29_5_2),
		.out_wire_0_3(horizontal_tile_29_4_to_tile_29_5_3),
		.in_wire_0_0(horizontal_tile_29_5_to_tile_29_4_0),
		.in_wire_0_1(horizontal_tile_29_5_to_tile_29_4_1),
		.in_wire_0_2(horizontal_tile_29_5_to_tile_29_4_2),
		.in_wire_0_3(horizontal_tile_29_5_to_tile_29_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(933)
	);

	pe_tile pe_tile_29_5(
		.out_wire_3_0(vertical_tile_29_5_to_tile_28_5_0),
		.out_wire_3_1(vertical_tile_29_5_to_tile_28_5_1),
		.out_wire_3_2(vertical_tile_29_5_to_tile_28_5_2),
		.out_wire_3_3(vertical_tile_29_5_to_tile_28_5_3),
		.in_wire_3_0(vertical_tile_28_5_to_tile_29_5_0),
		.in_wire_3_1(vertical_tile_28_5_to_tile_29_5_1),
		.in_wire_3_2(vertical_tile_28_5_to_tile_29_5_2),
		.in_wire_3_3(vertical_tile_28_5_to_tile_29_5_3),
		.out_wire_1_0(vertical_tile_29_5_to_tile_30_5_0),
		.out_wire_1_1(vertical_tile_29_5_to_tile_30_5_1),
		.out_wire_1_2(vertical_tile_29_5_to_tile_30_5_2),
		.out_wire_1_3(vertical_tile_29_5_to_tile_30_5_3),
		.in_wire_1_0(vertical_tile_30_5_to_tile_29_5_0),
		.in_wire_1_1(vertical_tile_30_5_to_tile_29_5_1),
		.in_wire_1_2(vertical_tile_30_5_to_tile_29_5_2),
		.in_wire_1_3(vertical_tile_30_5_to_tile_29_5_3),
		.out_wire_2_0(horizontal_tile_29_5_to_tile_29_4_0),
		.out_wire_2_1(horizontal_tile_29_5_to_tile_29_4_1),
		.out_wire_2_2(horizontal_tile_29_5_to_tile_29_4_2),
		.out_wire_2_3(horizontal_tile_29_5_to_tile_29_4_3),
		.in_wire_2_0(horizontal_tile_29_4_to_tile_29_5_0),
		.in_wire_2_1(horizontal_tile_29_4_to_tile_29_5_1),
		.in_wire_2_2(horizontal_tile_29_4_to_tile_29_5_2),
		.in_wire_2_3(horizontal_tile_29_4_to_tile_29_5_3),
		.out_wire_0_0(horizontal_tile_29_5_to_tile_29_6_0),
		.out_wire_0_1(horizontal_tile_29_5_to_tile_29_6_1),
		.out_wire_0_2(horizontal_tile_29_5_to_tile_29_6_2),
		.out_wire_0_3(horizontal_tile_29_5_to_tile_29_6_3),
		.in_wire_0_0(horizontal_tile_29_6_to_tile_29_5_0),
		.in_wire_0_1(horizontal_tile_29_6_to_tile_29_5_1),
		.in_wire_0_2(horizontal_tile_29_6_to_tile_29_5_2),
		.in_wire_0_3(horizontal_tile_29_6_to_tile_29_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(934)
	);

	pe_tile pe_tile_29_6(
		.out_wire_3_0(vertical_tile_29_6_to_tile_28_6_0),
		.out_wire_3_1(vertical_tile_29_6_to_tile_28_6_1),
		.out_wire_3_2(vertical_tile_29_6_to_tile_28_6_2),
		.out_wire_3_3(vertical_tile_29_6_to_tile_28_6_3),
		.in_wire_3_0(vertical_tile_28_6_to_tile_29_6_0),
		.in_wire_3_1(vertical_tile_28_6_to_tile_29_6_1),
		.in_wire_3_2(vertical_tile_28_6_to_tile_29_6_2),
		.in_wire_3_3(vertical_tile_28_6_to_tile_29_6_3),
		.out_wire_1_0(vertical_tile_29_6_to_tile_30_6_0),
		.out_wire_1_1(vertical_tile_29_6_to_tile_30_6_1),
		.out_wire_1_2(vertical_tile_29_6_to_tile_30_6_2),
		.out_wire_1_3(vertical_tile_29_6_to_tile_30_6_3),
		.in_wire_1_0(vertical_tile_30_6_to_tile_29_6_0),
		.in_wire_1_1(vertical_tile_30_6_to_tile_29_6_1),
		.in_wire_1_2(vertical_tile_30_6_to_tile_29_6_2),
		.in_wire_1_3(vertical_tile_30_6_to_tile_29_6_3),
		.out_wire_2_0(horizontal_tile_29_6_to_tile_29_5_0),
		.out_wire_2_1(horizontal_tile_29_6_to_tile_29_5_1),
		.out_wire_2_2(horizontal_tile_29_6_to_tile_29_5_2),
		.out_wire_2_3(horizontal_tile_29_6_to_tile_29_5_3),
		.in_wire_2_0(horizontal_tile_29_5_to_tile_29_6_0),
		.in_wire_2_1(horizontal_tile_29_5_to_tile_29_6_1),
		.in_wire_2_2(horizontal_tile_29_5_to_tile_29_6_2),
		.in_wire_2_3(horizontal_tile_29_5_to_tile_29_6_3),
		.out_wire_0_0(horizontal_tile_29_6_to_tile_29_7_0),
		.out_wire_0_1(horizontal_tile_29_6_to_tile_29_7_1),
		.out_wire_0_2(horizontal_tile_29_6_to_tile_29_7_2),
		.out_wire_0_3(horizontal_tile_29_6_to_tile_29_7_3),
		.in_wire_0_0(horizontal_tile_29_7_to_tile_29_6_0),
		.in_wire_0_1(horizontal_tile_29_7_to_tile_29_6_1),
		.in_wire_0_2(horizontal_tile_29_7_to_tile_29_6_2),
		.in_wire_0_3(horizontal_tile_29_7_to_tile_29_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(935)
	);

	pe_tile pe_tile_29_7(
		.out_wire_3_0(vertical_tile_29_7_to_tile_28_7_0),
		.out_wire_3_1(vertical_tile_29_7_to_tile_28_7_1),
		.out_wire_3_2(vertical_tile_29_7_to_tile_28_7_2),
		.out_wire_3_3(vertical_tile_29_7_to_tile_28_7_3),
		.in_wire_3_0(vertical_tile_28_7_to_tile_29_7_0),
		.in_wire_3_1(vertical_tile_28_7_to_tile_29_7_1),
		.in_wire_3_2(vertical_tile_28_7_to_tile_29_7_2),
		.in_wire_3_3(vertical_tile_28_7_to_tile_29_7_3),
		.out_wire_1_0(vertical_tile_29_7_to_tile_30_7_0),
		.out_wire_1_1(vertical_tile_29_7_to_tile_30_7_1),
		.out_wire_1_2(vertical_tile_29_7_to_tile_30_7_2),
		.out_wire_1_3(vertical_tile_29_7_to_tile_30_7_3),
		.in_wire_1_0(vertical_tile_30_7_to_tile_29_7_0),
		.in_wire_1_1(vertical_tile_30_7_to_tile_29_7_1),
		.in_wire_1_2(vertical_tile_30_7_to_tile_29_7_2),
		.in_wire_1_3(vertical_tile_30_7_to_tile_29_7_3),
		.out_wire_2_0(horizontal_tile_29_7_to_tile_29_6_0),
		.out_wire_2_1(horizontal_tile_29_7_to_tile_29_6_1),
		.out_wire_2_2(horizontal_tile_29_7_to_tile_29_6_2),
		.out_wire_2_3(horizontal_tile_29_7_to_tile_29_6_3),
		.in_wire_2_0(horizontal_tile_29_6_to_tile_29_7_0),
		.in_wire_2_1(horizontal_tile_29_6_to_tile_29_7_1),
		.in_wire_2_2(horizontal_tile_29_6_to_tile_29_7_2),
		.in_wire_2_3(horizontal_tile_29_6_to_tile_29_7_3),
		.out_wire_0_0(horizontal_tile_29_7_to_tile_29_8_0),
		.out_wire_0_1(horizontal_tile_29_7_to_tile_29_8_1),
		.out_wire_0_2(horizontal_tile_29_7_to_tile_29_8_2),
		.out_wire_0_3(horizontal_tile_29_7_to_tile_29_8_3),
		.in_wire_0_0(horizontal_tile_29_8_to_tile_29_7_0),
		.in_wire_0_1(horizontal_tile_29_8_to_tile_29_7_1),
		.in_wire_0_2(horizontal_tile_29_8_to_tile_29_7_2),
		.in_wire_0_3(horizontal_tile_29_8_to_tile_29_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(936)
	);

	pe_tile pe_tile_29_8(
		.out_wire_3_0(vertical_tile_29_8_to_tile_28_8_0),
		.out_wire_3_1(vertical_tile_29_8_to_tile_28_8_1),
		.out_wire_3_2(vertical_tile_29_8_to_tile_28_8_2),
		.out_wire_3_3(vertical_tile_29_8_to_tile_28_8_3),
		.in_wire_3_0(vertical_tile_28_8_to_tile_29_8_0),
		.in_wire_3_1(vertical_tile_28_8_to_tile_29_8_1),
		.in_wire_3_2(vertical_tile_28_8_to_tile_29_8_2),
		.in_wire_3_3(vertical_tile_28_8_to_tile_29_8_3),
		.out_wire_1_0(vertical_tile_29_8_to_tile_30_8_0),
		.out_wire_1_1(vertical_tile_29_8_to_tile_30_8_1),
		.out_wire_1_2(vertical_tile_29_8_to_tile_30_8_2),
		.out_wire_1_3(vertical_tile_29_8_to_tile_30_8_3),
		.in_wire_1_0(vertical_tile_30_8_to_tile_29_8_0),
		.in_wire_1_1(vertical_tile_30_8_to_tile_29_8_1),
		.in_wire_1_2(vertical_tile_30_8_to_tile_29_8_2),
		.in_wire_1_3(vertical_tile_30_8_to_tile_29_8_3),
		.out_wire_2_0(horizontal_tile_29_8_to_tile_29_7_0),
		.out_wire_2_1(horizontal_tile_29_8_to_tile_29_7_1),
		.out_wire_2_2(horizontal_tile_29_8_to_tile_29_7_2),
		.out_wire_2_3(horizontal_tile_29_8_to_tile_29_7_3),
		.in_wire_2_0(horizontal_tile_29_7_to_tile_29_8_0),
		.in_wire_2_1(horizontal_tile_29_7_to_tile_29_8_1),
		.in_wire_2_2(horizontal_tile_29_7_to_tile_29_8_2),
		.in_wire_2_3(horizontal_tile_29_7_to_tile_29_8_3),
		.out_wire_0_0(horizontal_tile_29_8_to_tile_29_9_0),
		.out_wire_0_1(horizontal_tile_29_8_to_tile_29_9_1),
		.out_wire_0_2(horizontal_tile_29_8_to_tile_29_9_2),
		.out_wire_0_3(horizontal_tile_29_8_to_tile_29_9_3),
		.in_wire_0_0(horizontal_tile_29_9_to_tile_29_8_0),
		.in_wire_0_1(horizontal_tile_29_9_to_tile_29_8_1),
		.in_wire_0_2(horizontal_tile_29_9_to_tile_29_8_2),
		.in_wire_0_3(horizontal_tile_29_9_to_tile_29_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(937)
	);

	pe_tile pe_tile_29_9(
		.out_wire_3_0(vertical_tile_29_9_to_tile_28_9_0),
		.out_wire_3_1(vertical_tile_29_9_to_tile_28_9_1),
		.out_wire_3_2(vertical_tile_29_9_to_tile_28_9_2),
		.out_wire_3_3(vertical_tile_29_9_to_tile_28_9_3),
		.in_wire_3_0(vertical_tile_28_9_to_tile_29_9_0),
		.in_wire_3_1(vertical_tile_28_9_to_tile_29_9_1),
		.in_wire_3_2(vertical_tile_28_9_to_tile_29_9_2),
		.in_wire_3_3(vertical_tile_28_9_to_tile_29_9_3),
		.out_wire_1_0(vertical_tile_29_9_to_tile_30_9_0),
		.out_wire_1_1(vertical_tile_29_9_to_tile_30_9_1),
		.out_wire_1_2(vertical_tile_29_9_to_tile_30_9_2),
		.out_wire_1_3(vertical_tile_29_9_to_tile_30_9_3),
		.in_wire_1_0(vertical_tile_30_9_to_tile_29_9_0),
		.in_wire_1_1(vertical_tile_30_9_to_tile_29_9_1),
		.in_wire_1_2(vertical_tile_30_9_to_tile_29_9_2),
		.in_wire_1_3(vertical_tile_30_9_to_tile_29_9_3),
		.out_wire_2_0(horizontal_tile_29_9_to_tile_29_8_0),
		.out_wire_2_1(horizontal_tile_29_9_to_tile_29_8_1),
		.out_wire_2_2(horizontal_tile_29_9_to_tile_29_8_2),
		.out_wire_2_3(horizontal_tile_29_9_to_tile_29_8_3),
		.in_wire_2_0(horizontal_tile_29_8_to_tile_29_9_0),
		.in_wire_2_1(horizontal_tile_29_8_to_tile_29_9_1),
		.in_wire_2_2(horizontal_tile_29_8_to_tile_29_9_2),
		.in_wire_2_3(horizontal_tile_29_8_to_tile_29_9_3),
		.out_wire_0_0(horizontal_tile_29_9_to_tile_29_10_0),
		.out_wire_0_1(horizontal_tile_29_9_to_tile_29_10_1),
		.out_wire_0_2(horizontal_tile_29_9_to_tile_29_10_2),
		.out_wire_0_3(horizontal_tile_29_9_to_tile_29_10_3),
		.in_wire_0_0(horizontal_tile_29_10_to_tile_29_9_0),
		.in_wire_0_1(horizontal_tile_29_10_to_tile_29_9_1),
		.in_wire_0_2(horizontal_tile_29_10_to_tile_29_9_2),
		.in_wire_0_3(horizontal_tile_29_10_to_tile_29_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(938)
	);

	pe_tile pe_tile_29_10(
		.out_wire_3_0(vertical_tile_29_10_to_tile_28_10_0),
		.out_wire_3_1(vertical_tile_29_10_to_tile_28_10_1),
		.out_wire_3_2(vertical_tile_29_10_to_tile_28_10_2),
		.out_wire_3_3(vertical_tile_29_10_to_tile_28_10_3),
		.in_wire_3_0(vertical_tile_28_10_to_tile_29_10_0),
		.in_wire_3_1(vertical_tile_28_10_to_tile_29_10_1),
		.in_wire_3_2(vertical_tile_28_10_to_tile_29_10_2),
		.in_wire_3_3(vertical_tile_28_10_to_tile_29_10_3),
		.out_wire_1_0(vertical_tile_29_10_to_tile_30_10_0),
		.out_wire_1_1(vertical_tile_29_10_to_tile_30_10_1),
		.out_wire_1_2(vertical_tile_29_10_to_tile_30_10_2),
		.out_wire_1_3(vertical_tile_29_10_to_tile_30_10_3),
		.in_wire_1_0(vertical_tile_30_10_to_tile_29_10_0),
		.in_wire_1_1(vertical_tile_30_10_to_tile_29_10_1),
		.in_wire_1_2(vertical_tile_30_10_to_tile_29_10_2),
		.in_wire_1_3(vertical_tile_30_10_to_tile_29_10_3),
		.out_wire_2_0(horizontal_tile_29_10_to_tile_29_9_0),
		.out_wire_2_1(horizontal_tile_29_10_to_tile_29_9_1),
		.out_wire_2_2(horizontal_tile_29_10_to_tile_29_9_2),
		.out_wire_2_3(horizontal_tile_29_10_to_tile_29_9_3),
		.in_wire_2_0(horizontal_tile_29_9_to_tile_29_10_0),
		.in_wire_2_1(horizontal_tile_29_9_to_tile_29_10_1),
		.in_wire_2_2(horizontal_tile_29_9_to_tile_29_10_2),
		.in_wire_2_3(horizontal_tile_29_9_to_tile_29_10_3),
		.out_wire_0_0(horizontal_tile_29_10_to_tile_29_11_0),
		.out_wire_0_1(horizontal_tile_29_10_to_tile_29_11_1),
		.out_wire_0_2(horizontal_tile_29_10_to_tile_29_11_2),
		.out_wire_0_3(horizontal_tile_29_10_to_tile_29_11_3),
		.in_wire_0_0(horizontal_tile_29_11_to_tile_29_10_0),
		.in_wire_0_1(horizontal_tile_29_11_to_tile_29_10_1),
		.in_wire_0_2(horizontal_tile_29_11_to_tile_29_10_2),
		.in_wire_0_3(horizontal_tile_29_11_to_tile_29_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(939)
	);

	pe_tile pe_tile_29_11(
		.out_wire_3_0(vertical_tile_29_11_to_tile_28_11_0),
		.out_wire_3_1(vertical_tile_29_11_to_tile_28_11_1),
		.out_wire_3_2(vertical_tile_29_11_to_tile_28_11_2),
		.out_wire_3_3(vertical_tile_29_11_to_tile_28_11_3),
		.in_wire_3_0(vertical_tile_28_11_to_tile_29_11_0),
		.in_wire_3_1(vertical_tile_28_11_to_tile_29_11_1),
		.in_wire_3_2(vertical_tile_28_11_to_tile_29_11_2),
		.in_wire_3_3(vertical_tile_28_11_to_tile_29_11_3),
		.out_wire_1_0(vertical_tile_29_11_to_tile_30_11_0),
		.out_wire_1_1(vertical_tile_29_11_to_tile_30_11_1),
		.out_wire_1_2(vertical_tile_29_11_to_tile_30_11_2),
		.out_wire_1_3(vertical_tile_29_11_to_tile_30_11_3),
		.in_wire_1_0(vertical_tile_30_11_to_tile_29_11_0),
		.in_wire_1_1(vertical_tile_30_11_to_tile_29_11_1),
		.in_wire_1_2(vertical_tile_30_11_to_tile_29_11_2),
		.in_wire_1_3(vertical_tile_30_11_to_tile_29_11_3),
		.out_wire_2_0(horizontal_tile_29_11_to_tile_29_10_0),
		.out_wire_2_1(horizontal_tile_29_11_to_tile_29_10_1),
		.out_wire_2_2(horizontal_tile_29_11_to_tile_29_10_2),
		.out_wire_2_3(horizontal_tile_29_11_to_tile_29_10_3),
		.in_wire_2_0(horizontal_tile_29_10_to_tile_29_11_0),
		.in_wire_2_1(horizontal_tile_29_10_to_tile_29_11_1),
		.in_wire_2_2(horizontal_tile_29_10_to_tile_29_11_2),
		.in_wire_2_3(horizontal_tile_29_10_to_tile_29_11_3),
		.out_wire_0_0(horizontal_tile_29_11_to_tile_29_12_0),
		.out_wire_0_1(horizontal_tile_29_11_to_tile_29_12_1),
		.out_wire_0_2(horizontal_tile_29_11_to_tile_29_12_2),
		.out_wire_0_3(horizontal_tile_29_11_to_tile_29_12_3),
		.in_wire_0_0(horizontal_tile_29_12_to_tile_29_11_0),
		.in_wire_0_1(horizontal_tile_29_12_to_tile_29_11_1),
		.in_wire_0_2(horizontal_tile_29_12_to_tile_29_11_2),
		.in_wire_0_3(horizontal_tile_29_12_to_tile_29_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(940)
	);

	pe_tile pe_tile_29_12(
		.out_wire_3_0(vertical_tile_29_12_to_tile_28_12_0),
		.out_wire_3_1(vertical_tile_29_12_to_tile_28_12_1),
		.out_wire_3_2(vertical_tile_29_12_to_tile_28_12_2),
		.out_wire_3_3(vertical_tile_29_12_to_tile_28_12_3),
		.in_wire_3_0(vertical_tile_28_12_to_tile_29_12_0),
		.in_wire_3_1(vertical_tile_28_12_to_tile_29_12_1),
		.in_wire_3_2(vertical_tile_28_12_to_tile_29_12_2),
		.in_wire_3_3(vertical_tile_28_12_to_tile_29_12_3),
		.out_wire_1_0(vertical_tile_29_12_to_tile_30_12_0),
		.out_wire_1_1(vertical_tile_29_12_to_tile_30_12_1),
		.out_wire_1_2(vertical_tile_29_12_to_tile_30_12_2),
		.out_wire_1_3(vertical_tile_29_12_to_tile_30_12_3),
		.in_wire_1_0(vertical_tile_30_12_to_tile_29_12_0),
		.in_wire_1_1(vertical_tile_30_12_to_tile_29_12_1),
		.in_wire_1_2(vertical_tile_30_12_to_tile_29_12_2),
		.in_wire_1_3(vertical_tile_30_12_to_tile_29_12_3),
		.out_wire_2_0(horizontal_tile_29_12_to_tile_29_11_0),
		.out_wire_2_1(horizontal_tile_29_12_to_tile_29_11_1),
		.out_wire_2_2(horizontal_tile_29_12_to_tile_29_11_2),
		.out_wire_2_3(horizontal_tile_29_12_to_tile_29_11_3),
		.in_wire_2_0(horizontal_tile_29_11_to_tile_29_12_0),
		.in_wire_2_1(horizontal_tile_29_11_to_tile_29_12_1),
		.in_wire_2_2(horizontal_tile_29_11_to_tile_29_12_2),
		.in_wire_2_3(horizontal_tile_29_11_to_tile_29_12_3),
		.out_wire_0_0(horizontal_tile_29_12_to_tile_29_13_0),
		.out_wire_0_1(horizontal_tile_29_12_to_tile_29_13_1),
		.out_wire_0_2(horizontal_tile_29_12_to_tile_29_13_2),
		.out_wire_0_3(horizontal_tile_29_12_to_tile_29_13_3),
		.in_wire_0_0(horizontal_tile_29_13_to_tile_29_12_0),
		.in_wire_0_1(horizontal_tile_29_13_to_tile_29_12_1),
		.in_wire_0_2(horizontal_tile_29_13_to_tile_29_12_2),
		.in_wire_0_3(horizontal_tile_29_13_to_tile_29_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(941)
	);

	pe_tile pe_tile_29_13(
		.out_wire_3_0(vertical_tile_29_13_to_tile_28_13_0),
		.out_wire_3_1(vertical_tile_29_13_to_tile_28_13_1),
		.out_wire_3_2(vertical_tile_29_13_to_tile_28_13_2),
		.out_wire_3_3(vertical_tile_29_13_to_tile_28_13_3),
		.in_wire_3_0(vertical_tile_28_13_to_tile_29_13_0),
		.in_wire_3_1(vertical_tile_28_13_to_tile_29_13_1),
		.in_wire_3_2(vertical_tile_28_13_to_tile_29_13_2),
		.in_wire_3_3(vertical_tile_28_13_to_tile_29_13_3),
		.out_wire_1_0(vertical_tile_29_13_to_tile_30_13_0),
		.out_wire_1_1(vertical_tile_29_13_to_tile_30_13_1),
		.out_wire_1_2(vertical_tile_29_13_to_tile_30_13_2),
		.out_wire_1_3(vertical_tile_29_13_to_tile_30_13_3),
		.in_wire_1_0(vertical_tile_30_13_to_tile_29_13_0),
		.in_wire_1_1(vertical_tile_30_13_to_tile_29_13_1),
		.in_wire_1_2(vertical_tile_30_13_to_tile_29_13_2),
		.in_wire_1_3(vertical_tile_30_13_to_tile_29_13_3),
		.out_wire_2_0(horizontal_tile_29_13_to_tile_29_12_0),
		.out_wire_2_1(horizontal_tile_29_13_to_tile_29_12_1),
		.out_wire_2_2(horizontal_tile_29_13_to_tile_29_12_2),
		.out_wire_2_3(horizontal_tile_29_13_to_tile_29_12_3),
		.in_wire_2_0(horizontal_tile_29_12_to_tile_29_13_0),
		.in_wire_2_1(horizontal_tile_29_12_to_tile_29_13_1),
		.in_wire_2_2(horizontal_tile_29_12_to_tile_29_13_2),
		.in_wire_2_3(horizontal_tile_29_12_to_tile_29_13_3),
		.out_wire_0_0(horizontal_tile_29_13_to_tile_29_14_0),
		.out_wire_0_1(horizontal_tile_29_13_to_tile_29_14_1),
		.out_wire_0_2(horizontal_tile_29_13_to_tile_29_14_2),
		.out_wire_0_3(horizontal_tile_29_13_to_tile_29_14_3),
		.in_wire_0_0(horizontal_tile_29_14_to_tile_29_13_0),
		.in_wire_0_1(horizontal_tile_29_14_to_tile_29_13_1),
		.in_wire_0_2(horizontal_tile_29_14_to_tile_29_13_2),
		.in_wire_0_3(horizontal_tile_29_14_to_tile_29_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(942)
	);

	pe_tile pe_tile_29_14(
		.out_wire_3_0(vertical_tile_29_14_to_tile_28_14_0),
		.out_wire_3_1(vertical_tile_29_14_to_tile_28_14_1),
		.out_wire_3_2(vertical_tile_29_14_to_tile_28_14_2),
		.out_wire_3_3(vertical_tile_29_14_to_tile_28_14_3),
		.in_wire_3_0(vertical_tile_28_14_to_tile_29_14_0),
		.in_wire_3_1(vertical_tile_28_14_to_tile_29_14_1),
		.in_wire_3_2(vertical_tile_28_14_to_tile_29_14_2),
		.in_wire_3_3(vertical_tile_28_14_to_tile_29_14_3),
		.out_wire_1_0(vertical_tile_29_14_to_tile_30_14_0),
		.out_wire_1_1(vertical_tile_29_14_to_tile_30_14_1),
		.out_wire_1_2(vertical_tile_29_14_to_tile_30_14_2),
		.out_wire_1_3(vertical_tile_29_14_to_tile_30_14_3),
		.in_wire_1_0(vertical_tile_30_14_to_tile_29_14_0),
		.in_wire_1_1(vertical_tile_30_14_to_tile_29_14_1),
		.in_wire_1_2(vertical_tile_30_14_to_tile_29_14_2),
		.in_wire_1_3(vertical_tile_30_14_to_tile_29_14_3),
		.out_wire_2_0(horizontal_tile_29_14_to_tile_29_13_0),
		.out_wire_2_1(horizontal_tile_29_14_to_tile_29_13_1),
		.out_wire_2_2(horizontal_tile_29_14_to_tile_29_13_2),
		.out_wire_2_3(horizontal_tile_29_14_to_tile_29_13_3),
		.in_wire_2_0(horizontal_tile_29_13_to_tile_29_14_0),
		.in_wire_2_1(horizontal_tile_29_13_to_tile_29_14_1),
		.in_wire_2_2(horizontal_tile_29_13_to_tile_29_14_2),
		.in_wire_2_3(horizontal_tile_29_13_to_tile_29_14_3),
		.out_wire_0_0(horizontal_tile_29_14_to_tile_29_15_0),
		.out_wire_0_1(horizontal_tile_29_14_to_tile_29_15_1),
		.out_wire_0_2(horizontal_tile_29_14_to_tile_29_15_2),
		.out_wire_0_3(horizontal_tile_29_14_to_tile_29_15_3),
		.in_wire_0_0(horizontal_tile_29_15_to_tile_29_14_0),
		.in_wire_0_1(horizontal_tile_29_15_to_tile_29_14_1),
		.in_wire_0_2(horizontal_tile_29_15_to_tile_29_14_2),
		.in_wire_0_3(horizontal_tile_29_15_to_tile_29_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(943)
	);

	pe_tile pe_tile_29_15(
		.out_wire_3_0(vertical_tile_29_15_to_tile_28_15_0),
		.out_wire_3_1(vertical_tile_29_15_to_tile_28_15_1),
		.out_wire_3_2(vertical_tile_29_15_to_tile_28_15_2),
		.out_wire_3_3(vertical_tile_29_15_to_tile_28_15_3),
		.in_wire_3_0(vertical_tile_28_15_to_tile_29_15_0),
		.in_wire_3_1(vertical_tile_28_15_to_tile_29_15_1),
		.in_wire_3_2(vertical_tile_28_15_to_tile_29_15_2),
		.in_wire_3_3(vertical_tile_28_15_to_tile_29_15_3),
		.out_wire_1_0(vertical_tile_29_15_to_tile_30_15_0),
		.out_wire_1_1(vertical_tile_29_15_to_tile_30_15_1),
		.out_wire_1_2(vertical_tile_29_15_to_tile_30_15_2),
		.out_wire_1_3(vertical_tile_29_15_to_tile_30_15_3),
		.in_wire_1_0(vertical_tile_30_15_to_tile_29_15_0),
		.in_wire_1_1(vertical_tile_30_15_to_tile_29_15_1),
		.in_wire_1_2(vertical_tile_30_15_to_tile_29_15_2),
		.in_wire_1_3(vertical_tile_30_15_to_tile_29_15_3),
		.out_wire_2_0(horizontal_tile_29_15_to_tile_29_14_0),
		.out_wire_2_1(horizontal_tile_29_15_to_tile_29_14_1),
		.out_wire_2_2(horizontal_tile_29_15_to_tile_29_14_2),
		.out_wire_2_3(horizontal_tile_29_15_to_tile_29_14_3),
		.in_wire_2_0(horizontal_tile_29_14_to_tile_29_15_0),
		.in_wire_2_1(horizontal_tile_29_14_to_tile_29_15_1),
		.in_wire_2_2(horizontal_tile_29_14_to_tile_29_15_2),
		.in_wire_2_3(horizontal_tile_29_14_to_tile_29_15_3),
		.out_wire_0_0(horizontal_tile_29_15_to_tile_29_16_0),
		.out_wire_0_1(horizontal_tile_29_15_to_tile_29_16_1),
		.out_wire_0_2(horizontal_tile_29_15_to_tile_29_16_2),
		.out_wire_0_3(horizontal_tile_29_15_to_tile_29_16_3),
		.in_wire_0_0(horizontal_tile_29_16_to_tile_29_15_0),
		.in_wire_0_1(horizontal_tile_29_16_to_tile_29_15_1),
		.in_wire_0_2(horizontal_tile_29_16_to_tile_29_15_2),
		.in_wire_0_3(horizontal_tile_29_16_to_tile_29_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(944)
	);

	pe_tile pe_tile_29_16(
		.out_wire_3_0(vertical_tile_29_16_to_tile_28_16_0),
		.out_wire_3_1(vertical_tile_29_16_to_tile_28_16_1),
		.out_wire_3_2(vertical_tile_29_16_to_tile_28_16_2),
		.out_wire_3_3(vertical_tile_29_16_to_tile_28_16_3),
		.in_wire_3_0(vertical_tile_28_16_to_tile_29_16_0),
		.in_wire_3_1(vertical_tile_28_16_to_tile_29_16_1),
		.in_wire_3_2(vertical_tile_28_16_to_tile_29_16_2),
		.in_wire_3_3(vertical_tile_28_16_to_tile_29_16_3),
		.out_wire_1_0(vertical_tile_29_16_to_tile_30_16_0),
		.out_wire_1_1(vertical_tile_29_16_to_tile_30_16_1),
		.out_wire_1_2(vertical_tile_29_16_to_tile_30_16_2),
		.out_wire_1_3(vertical_tile_29_16_to_tile_30_16_3),
		.in_wire_1_0(vertical_tile_30_16_to_tile_29_16_0),
		.in_wire_1_1(vertical_tile_30_16_to_tile_29_16_1),
		.in_wire_1_2(vertical_tile_30_16_to_tile_29_16_2),
		.in_wire_1_3(vertical_tile_30_16_to_tile_29_16_3),
		.out_wire_2_0(horizontal_tile_29_16_to_tile_29_15_0),
		.out_wire_2_1(horizontal_tile_29_16_to_tile_29_15_1),
		.out_wire_2_2(horizontal_tile_29_16_to_tile_29_15_2),
		.out_wire_2_3(horizontal_tile_29_16_to_tile_29_15_3),
		.in_wire_2_0(horizontal_tile_29_15_to_tile_29_16_0),
		.in_wire_2_1(horizontal_tile_29_15_to_tile_29_16_1),
		.in_wire_2_2(horizontal_tile_29_15_to_tile_29_16_2),
		.in_wire_2_3(horizontal_tile_29_15_to_tile_29_16_3),
		.out_wire_0_0(horizontal_tile_29_16_to_tile_29_17_0),
		.out_wire_0_1(horizontal_tile_29_16_to_tile_29_17_1),
		.out_wire_0_2(horizontal_tile_29_16_to_tile_29_17_2),
		.out_wire_0_3(horizontal_tile_29_16_to_tile_29_17_3),
		.in_wire_0_0(horizontal_tile_29_17_to_tile_29_16_0),
		.in_wire_0_1(horizontal_tile_29_17_to_tile_29_16_1),
		.in_wire_0_2(horizontal_tile_29_17_to_tile_29_16_2),
		.in_wire_0_3(horizontal_tile_29_17_to_tile_29_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(945)
	);

	pe_tile pe_tile_29_17(
		.out_wire_3_0(vertical_tile_29_17_to_tile_28_17_0),
		.out_wire_3_1(vertical_tile_29_17_to_tile_28_17_1),
		.out_wire_3_2(vertical_tile_29_17_to_tile_28_17_2),
		.out_wire_3_3(vertical_tile_29_17_to_tile_28_17_3),
		.in_wire_3_0(vertical_tile_28_17_to_tile_29_17_0),
		.in_wire_3_1(vertical_tile_28_17_to_tile_29_17_1),
		.in_wire_3_2(vertical_tile_28_17_to_tile_29_17_2),
		.in_wire_3_3(vertical_tile_28_17_to_tile_29_17_3),
		.out_wire_1_0(vertical_tile_29_17_to_tile_30_17_0),
		.out_wire_1_1(vertical_tile_29_17_to_tile_30_17_1),
		.out_wire_1_2(vertical_tile_29_17_to_tile_30_17_2),
		.out_wire_1_3(vertical_tile_29_17_to_tile_30_17_3),
		.in_wire_1_0(vertical_tile_30_17_to_tile_29_17_0),
		.in_wire_1_1(vertical_tile_30_17_to_tile_29_17_1),
		.in_wire_1_2(vertical_tile_30_17_to_tile_29_17_2),
		.in_wire_1_3(vertical_tile_30_17_to_tile_29_17_3),
		.out_wire_2_0(horizontal_tile_29_17_to_tile_29_16_0),
		.out_wire_2_1(horizontal_tile_29_17_to_tile_29_16_1),
		.out_wire_2_2(horizontal_tile_29_17_to_tile_29_16_2),
		.out_wire_2_3(horizontal_tile_29_17_to_tile_29_16_3),
		.in_wire_2_0(horizontal_tile_29_16_to_tile_29_17_0),
		.in_wire_2_1(horizontal_tile_29_16_to_tile_29_17_1),
		.in_wire_2_2(horizontal_tile_29_16_to_tile_29_17_2),
		.in_wire_2_3(horizontal_tile_29_16_to_tile_29_17_3),
		.out_wire_0_0(horizontal_tile_29_17_to_tile_29_18_0),
		.out_wire_0_1(horizontal_tile_29_17_to_tile_29_18_1),
		.out_wire_0_2(horizontal_tile_29_17_to_tile_29_18_2),
		.out_wire_0_3(horizontal_tile_29_17_to_tile_29_18_3),
		.in_wire_0_0(horizontal_tile_29_18_to_tile_29_17_0),
		.in_wire_0_1(horizontal_tile_29_18_to_tile_29_17_1),
		.in_wire_0_2(horizontal_tile_29_18_to_tile_29_17_2),
		.in_wire_0_3(horizontal_tile_29_18_to_tile_29_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(946)
	);

	pe_tile pe_tile_29_18(
		.out_wire_3_0(vertical_tile_29_18_to_tile_28_18_0),
		.out_wire_3_1(vertical_tile_29_18_to_tile_28_18_1),
		.out_wire_3_2(vertical_tile_29_18_to_tile_28_18_2),
		.out_wire_3_3(vertical_tile_29_18_to_tile_28_18_3),
		.in_wire_3_0(vertical_tile_28_18_to_tile_29_18_0),
		.in_wire_3_1(vertical_tile_28_18_to_tile_29_18_1),
		.in_wire_3_2(vertical_tile_28_18_to_tile_29_18_2),
		.in_wire_3_3(vertical_tile_28_18_to_tile_29_18_3),
		.out_wire_1_0(vertical_tile_29_18_to_tile_30_18_0),
		.out_wire_1_1(vertical_tile_29_18_to_tile_30_18_1),
		.out_wire_1_2(vertical_tile_29_18_to_tile_30_18_2),
		.out_wire_1_3(vertical_tile_29_18_to_tile_30_18_3),
		.in_wire_1_0(vertical_tile_30_18_to_tile_29_18_0),
		.in_wire_1_1(vertical_tile_30_18_to_tile_29_18_1),
		.in_wire_1_2(vertical_tile_30_18_to_tile_29_18_2),
		.in_wire_1_3(vertical_tile_30_18_to_tile_29_18_3),
		.out_wire_2_0(horizontal_tile_29_18_to_tile_29_17_0),
		.out_wire_2_1(horizontal_tile_29_18_to_tile_29_17_1),
		.out_wire_2_2(horizontal_tile_29_18_to_tile_29_17_2),
		.out_wire_2_3(horizontal_tile_29_18_to_tile_29_17_3),
		.in_wire_2_0(horizontal_tile_29_17_to_tile_29_18_0),
		.in_wire_2_1(horizontal_tile_29_17_to_tile_29_18_1),
		.in_wire_2_2(horizontal_tile_29_17_to_tile_29_18_2),
		.in_wire_2_3(horizontal_tile_29_17_to_tile_29_18_3),
		.out_wire_0_0(horizontal_tile_29_18_to_tile_29_19_0),
		.out_wire_0_1(horizontal_tile_29_18_to_tile_29_19_1),
		.out_wire_0_2(horizontal_tile_29_18_to_tile_29_19_2),
		.out_wire_0_3(horizontal_tile_29_18_to_tile_29_19_3),
		.in_wire_0_0(horizontal_tile_29_19_to_tile_29_18_0),
		.in_wire_0_1(horizontal_tile_29_19_to_tile_29_18_1),
		.in_wire_0_2(horizontal_tile_29_19_to_tile_29_18_2),
		.in_wire_0_3(horizontal_tile_29_19_to_tile_29_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(947)
	);

	pe_tile pe_tile_29_19(
		.out_wire_3_0(vertical_tile_29_19_to_tile_28_19_0),
		.out_wire_3_1(vertical_tile_29_19_to_tile_28_19_1),
		.out_wire_3_2(vertical_tile_29_19_to_tile_28_19_2),
		.out_wire_3_3(vertical_tile_29_19_to_tile_28_19_3),
		.in_wire_3_0(vertical_tile_28_19_to_tile_29_19_0),
		.in_wire_3_1(vertical_tile_28_19_to_tile_29_19_1),
		.in_wire_3_2(vertical_tile_28_19_to_tile_29_19_2),
		.in_wire_3_3(vertical_tile_28_19_to_tile_29_19_3),
		.out_wire_1_0(vertical_tile_29_19_to_tile_30_19_0),
		.out_wire_1_1(vertical_tile_29_19_to_tile_30_19_1),
		.out_wire_1_2(vertical_tile_29_19_to_tile_30_19_2),
		.out_wire_1_3(vertical_tile_29_19_to_tile_30_19_3),
		.in_wire_1_0(vertical_tile_30_19_to_tile_29_19_0),
		.in_wire_1_1(vertical_tile_30_19_to_tile_29_19_1),
		.in_wire_1_2(vertical_tile_30_19_to_tile_29_19_2),
		.in_wire_1_3(vertical_tile_30_19_to_tile_29_19_3),
		.out_wire_2_0(horizontal_tile_29_19_to_tile_29_18_0),
		.out_wire_2_1(horizontal_tile_29_19_to_tile_29_18_1),
		.out_wire_2_2(horizontal_tile_29_19_to_tile_29_18_2),
		.out_wire_2_3(horizontal_tile_29_19_to_tile_29_18_3),
		.in_wire_2_0(horizontal_tile_29_18_to_tile_29_19_0),
		.in_wire_2_1(horizontal_tile_29_18_to_tile_29_19_1),
		.in_wire_2_2(horizontal_tile_29_18_to_tile_29_19_2),
		.in_wire_2_3(horizontal_tile_29_18_to_tile_29_19_3),
		.out_wire_0_0(horizontal_tile_29_19_to_tile_29_20_0),
		.out_wire_0_1(horizontal_tile_29_19_to_tile_29_20_1),
		.out_wire_0_2(horizontal_tile_29_19_to_tile_29_20_2),
		.out_wire_0_3(horizontal_tile_29_19_to_tile_29_20_3),
		.in_wire_0_0(horizontal_tile_29_20_to_tile_29_19_0),
		.in_wire_0_1(horizontal_tile_29_20_to_tile_29_19_1),
		.in_wire_0_2(horizontal_tile_29_20_to_tile_29_19_2),
		.in_wire_0_3(horizontal_tile_29_20_to_tile_29_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(948)
	);

	pe_tile pe_tile_29_20(
		.out_wire_3_0(vertical_tile_29_20_to_tile_28_20_0),
		.out_wire_3_1(vertical_tile_29_20_to_tile_28_20_1),
		.out_wire_3_2(vertical_tile_29_20_to_tile_28_20_2),
		.out_wire_3_3(vertical_tile_29_20_to_tile_28_20_3),
		.in_wire_3_0(vertical_tile_28_20_to_tile_29_20_0),
		.in_wire_3_1(vertical_tile_28_20_to_tile_29_20_1),
		.in_wire_3_2(vertical_tile_28_20_to_tile_29_20_2),
		.in_wire_3_3(vertical_tile_28_20_to_tile_29_20_3),
		.out_wire_1_0(vertical_tile_29_20_to_tile_30_20_0),
		.out_wire_1_1(vertical_tile_29_20_to_tile_30_20_1),
		.out_wire_1_2(vertical_tile_29_20_to_tile_30_20_2),
		.out_wire_1_3(vertical_tile_29_20_to_tile_30_20_3),
		.in_wire_1_0(vertical_tile_30_20_to_tile_29_20_0),
		.in_wire_1_1(vertical_tile_30_20_to_tile_29_20_1),
		.in_wire_1_2(vertical_tile_30_20_to_tile_29_20_2),
		.in_wire_1_3(vertical_tile_30_20_to_tile_29_20_3),
		.out_wire_2_0(horizontal_tile_29_20_to_tile_29_19_0),
		.out_wire_2_1(horizontal_tile_29_20_to_tile_29_19_1),
		.out_wire_2_2(horizontal_tile_29_20_to_tile_29_19_2),
		.out_wire_2_3(horizontal_tile_29_20_to_tile_29_19_3),
		.in_wire_2_0(horizontal_tile_29_19_to_tile_29_20_0),
		.in_wire_2_1(horizontal_tile_29_19_to_tile_29_20_1),
		.in_wire_2_2(horizontal_tile_29_19_to_tile_29_20_2),
		.in_wire_2_3(horizontal_tile_29_19_to_tile_29_20_3),
		.out_wire_0_0(horizontal_tile_29_20_to_tile_29_21_0),
		.out_wire_0_1(horizontal_tile_29_20_to_tile_29_21_1),
		.out_wire_0_2(horizontal_tile_29_20_to_tile_29_21_2),
		.out_wire_0_3(horizontal_tile_29_20_to_tile_29_21_3),
		.in_wire_0_0(horizontal_tile_29_21_to_tile_29_20_0),
		.in_wire_0_1(horizontal_tile_29_21_to_tile_29_20_1),
		.in_wire_0_2(horizontal_tile_29_21_to_tile_29_20_2),
		.in_wire_0_3(horizontal_tile_29_21_to_tile_29_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(949)
	);

	pe_tile pe_tile_29_21(
		.out_wire_3_0(vertical_tile_29_21_to_tile_28_21_0),
		.out_wire_3_1(vertical_tile_29_21_to_tile_28_21_1),
		.out_wire_3_2(vertical_tile_29_21_to_tile_28_21_2),
		.out_wire_3_3(vertical_tile_29_21_to_tile_28_21_3),
		.in_wire_3_0(vertical_tile_28_21_to_tile_29_21_0),
		.in_wire_3_1(vertical_tile_28_21_to_tile_29_21_1),
		.in_wire_3_2(vertical_tile_28_21_to_tile_29_21_2),
		.in_wire_3_3(vertical_tile_28_21_to_tile_29_21_3),
		.out_wire_1_0(vertical_tile_29_21_to_tile_30_21_0),
		.out_wire_1_1(vertical_tile_29_21_to_tile_30_21_1),
		.out_wire_1_2(vertical_tile_29_21_to_tile_30_21_2),
		.out_wire_1_3(vertical_tile_29_21_to_tile_30_21_3),
		.in_wire_1_0(vertical_tile_30_21_to_tile_29_21_0),
		.in_wire_1_1(vertical_tile_30_21_to_tile_29_21_1),
		.in_wire_1_2(vertical_tile_30_21_to_tile_29_21_2),
		.in_wire_1_3(vertical_tile_30_21_to_tile_29_21_3),
		.out_wire_2_0(horizontal_tile_29_21_to_tile_29_20_0),
		.out_wire_2_1(horizontal_tile_29_21_to_tile_29_20_1),
		.out_wire_2_2(horizontal_tile_29_21_to_tile_29_20_2),
		.out_wire_2_3(horizontal_tile_29_21_to_tile_29_20_3),
		.in_wire_2_0(horizontal_tile_29_20_to_tile_29_21_0),
		.in_wire_2_1(horizontal_tile_29_20_to_tile_29_21_1),
		.in_wire_2_2(horizontal_tile_29_20_to_tile_29_21_2),
		.in_wire_2_3(horizontal_tile_29_20_to_tile_29_21_3),
		.out_wire_0_0(horizontal_tile_29_21_to_tile_29_22_0),
		.out_wire_0_1(horizontal_tile_29_21_to_tile_29_22_1),
		.out_wire_0_2(horizontal_tile_29_21_to_tile_29_22_2),
		.out_wire_0_3(horizontal_tile_29_21_to_tile_29_22_3),
		.in_wire_0_0(horizontal_tile_29_22_to_tile_29_21_0),
		.in_wire_0_1(horizontal_tile_29_22_to_tile_29_21_1),
		.in_wire_0_2(horizontal_tile_29_22_to_tile_29_21_2),
		.in_wire_0_3(horizontal_tile_29_22_to_tile_29_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(950)
	);

	pe_tile pe_tile_29_22(
		.out_wire_3_0(vertical_tile_29_22_to_tile_28_22_0),
		.out_wire_3_1(vertical_tile_29_22_to_tile_28_22_1),
		.out_wire_3_2(vertical_tile_29_22_to_tile_28_22_2),
		.out_wire_3_3(vertical_tile_29_22_to_tile_28_22_3),
		.in_wire_3_0(vertical_tile_28_22_to_tile_29_22_0),
		.in_wire_3_1(vertical_tile_28_22_to_tile_29_22_1),
		.in_wire_3_2(vertical_tile_28_22_to_tile_29_22_2),
		.in_wire_3_3(vertical_tile_28_22_to_tile_29_22_3),
		.out_wire_1_0(vertical_tile_29_22_to_tile_30_22_0),
		.out_wire_1_1(vertical_tile_29_22_to_tile_30_22_1),
		.out_wire_1_2(vertical_tile_29_22_to_tile_30_22_2),
		.out_wire_1_3(vertical_tile_29_22_to_tile_30_22_3),
		.in_wire_1_0(vertical_tile_30_22_to_tile_29_22_0),
		.in_wire_1_1(vertical_tile_30_22_to_tile_29_22_1),
		.in_wire_1_2(vertical_tile_30_22_to_tile_29_22_2),
		.in_wire_1_3(vertical_tile_30_22_to_tile_29_22_3),
		.out_wire_2_0(horizontal_tile_29_22_to_tile_29_21_0),
		.out_wire_2_1(horizontal_tile_29_22_to_tile_29_21_1),
		.out_wire_2_2(horizontal_tile_29_22_to_tile_29_21_2),
		.out_wire_2_3(horizontal_tile_29_22_to_tile_29_21_3),
		.in_wire_2_0(horizontal_tile_29_21_to_tile_29_22_0),
		.in_wire_2_1(horizontal_tile_29_21_to_tile_29_22_1),
		.in_wire_2_2(horizontal_tile_29_21_to_tile_29_22_2),
		.in_wire_2_3(horizontal_tile_29_21_to_tile_29_22_3),
		.out_wire_0_0(horizontal_tile_29_22_to_tile_29_23_0),
		.out_wire_0_1(horizontal_tile_29_22_to_tile_29_23_1),
		.out_wire_0_2(horizontal_tile_29_22_to_tile_29_23_2),
		.out_wire_0_3(horizontal_tile_29_22_to_tile_29_23_3),
		.in_wire_0_0(horizontal_tile_29_23_to_tile_29_22_0),
		.in_wire_0_1(horizontal_tile_29_23_to_tile_29_22_1),
		.in_wire_0_2(horizontal_tile_29_23_to_tile_29_22_2),
		.in_wire_0_3(horizontal_tile_29_23_to_tile_29_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(951)
	);

	pe_tile pe_tile_29_23(
		.out_wire_3_0(vertical_tile_29_23_to_tile_28_23_0),
		.out_wire_3_1(vertical_tile_29_23_to_tile_28_23_1),
		.out_wire_3_2(vertical_tile_29_23_to_tile_28_23_2),
		.out_wire_3_3(vertical_tile_29_23_to_tile_28_23_3),
		.in_wire_3_0(vertical_tile_28_23_to_tile_29_23_0),
		.in_wire_3_1(vertical_tile_28_23_to_tile_29_23_1),
		.in_wire_3_2(vertical_tile_28_23_to_tile_29_23_2),
		.in_wire_3_3(vertical_tile_28_23_to_tile_29_23_3),
		.out_wire_1_0(vertical_tile_29_23_to_tile_30_23_0),
		.out_wire_1_1(vertical_tile_29_23_to_tile_30_23_1),
		.out_wire_1_2(vertical_tile_29_23_to_tile_30_23_2),
		.out_wire_1_3(vertical_tile_29_23_to_tile_30_23_3),
		.in_wire_1_0(vertical_tile_30_23_to_tile_29_23_0),
		.in_wire_1_1(vertical_tile_30_23_to_tile_29_23_1),
		.in_wire_1_2(vertical_tile_30_23_to_tile_29_23_2),
		.in_wire_1_3(vertical_tile_30_23_to_tile_29_23_3),
		.out_wire_2_0(horizontal_tile_29_23_to_tile_29_22_0),
		.out_wire_2_1(horizontal_tile_29_23_to_tile_29_22_1),
		.out_wire_2_2(horizontal_tile_29_23_to_tile_29_22_2),
		.out_wire_2_3(horizontal_tile_29_23_to_tile_29_22_3),
		.in_wire_2_0(horizontal_tile_29_22_to_tile_29_23_0),
		.in_wire_2_1(horizontal_tile_29_22_to_tile_29_23_1),
		.in_wire_2_2(horizontal_tile_29_22_to_tile_29_23_2),
		.in_wire_2_3(horizontal_tile_29_22_to_tile_29_23_3),
		.out_wire_0_0(horizontal_tile_29_23_to_tile_29_24_0),
		.out_wire_0_1(horizontal_tile_29_23_to_tile_29_24_1),
		.out_wire_0_2(horizontal_tile_29_23_to_tile_29_24_2),
		.out_wire_0_3(horizontal_tile_29_23_to_tile_29_24_3),
		.in_wire_0_0(horizontal_tile_29_24_to_tile_29_23_0),
		.in_wire_0_1(horizontal_tile_29_24_to_tile_29_23_1),
		.in_wire_0_2(horizontal_tile_29_24_to_tile_29_23_2),
		.in_wire_0_3(horizontal_tile_29_24_to_tile_29_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(952)
	);

	pe_tile pe_tile_29_24(
		.out_wire_3_0(vertical_tile_29_24_to_tile_28_24_0),
		.out_wire_3_1(vertical_tile_29_24_to_tile_28_24_1),
		.out_wire_3_2(vertical_tile_29_24_to_tile_28_24_2),
		.out_wire_3_3(vertical_tile_29_24_to_tile_28_24_3),
		.in_wire_3_0(vertical_tile_28_24_to_tile_29_24_0),
		.in_wire_3_1(vertical_tile_28_24_to_tile_29_24_1),
		.in_wire_3_2(vertical_tile_28_24_to_tile_29_24_2),
		.in_wire_3_3(vertical_tile_28_24_to_tile_29_24_3),
		.out_wire_1_0(vertical_tile_29_24_to_tile_30_24_0),
		.out_wire_1_1(vertical_tile_29_24_to_tile_30_24_1),
		.out_wire_1_2(vertical_tile_29_24_to_tile_30_24_2),
		.out_wire_1_3(vertical_tile_29_24_to_tile_30_24_3),
		.in_wire_1_0(vertical_tile_30_24_to_tile_29_24_0),
		.in_wire_1_1(vertical_tile_30_24_to_tile_29_24_1),
		.in_wire_1_2(vertical_tile_30_24_to_tile_29_24_2),
		.in_wire_1_3(vertical_tile_30_24_to_tile_29_24_3),
		.out_wire_2_0(horizontal_tile_29_24_to_tile_29_23_0),
		.out_wire_2_1(horizontal_tile_29_24_to_tile_29_23_1),
		.out_wire_2_2(horizontal_tile_29_24_to_tile_29_23_2),
		.out_wire_2_3(horizontal_tile_29_24_to_tile_29_23_3),
		.in_wire_2_0(horizontal_tile_29_23_to_tile_29_24_0),
		.in_wire_2_1(horizontal_tile_29_23_to_tile_29_24_1),
		.in_wire_2_2(horizontal_tile_29_23_to_tile_29_24_2),
		.in_wire_2_3(horizontal_tile_29_23_to_tile_29_24_3),
		.out_wire_0_0(horizontal_tile_29_24_to_tile_29_25_0),
		.out_wire_0_1(horizontal_tile_29_24_to_tile_29_25_1),
		.out_wire_0_2(horizontal_tile_29_24_to_tile_29_25_2),
		.out_wire_0_3(horizontal_tile_29_24_to_tile_29_25_3),
		.in_wire_0_0(horizontal_tile_29_25_to_tile_29_24_0),
		.in_wire_0_1(horizontal_tile_29_25_to_tile_29_24_1),
		.in_wire_0_2(horizontal_tile_29_25_to_tile_29_24_2),
		.in_wire_0_3(horizontal_tile_29_25_to_tile_29_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(953)
	);

	pe_tile pe_tile_29_25(
		.out_wire_3_0(vertical_tile_29_25_to_tile_28_25_0),
		.out_wire_3_1(vertical_tile_29_25_to_tile_28_25_1),
		.out_wire_3_2(vertical_tile_29_25_to_tile_28_25_2),
		.out_wire_3_3(vertical_tile_29_25_to_tile_28_25_3),
		.in_wire_3_0(vertical_tile_28_25_to_tile_29_25_0),
		.in_wire_3_1(vertical_tile_28_25_to_tile_29_25_1),
		.in_wire_3_2(vertical_tile_28_25_to_tile_29_25_2),
		.in_wire_3_3(vertical_tile_28_25_to_tile_29_25_3),
		.out_wire_1_0(vertical_tile_29_25_to_tile_30_25_0),
		.out_wire_1_1(vertical_tile_29_25_to_tile_30_25_1),
		.out_wire_1_2(vertical_tile_29_25_to_tile_30_25_2),
		.out_wire_1_3(vertical_tile_29_25_to_tile_30_25_3),
		.in_wire_1_0(vertical_tile_30_25_to_tile_29_25_0),
		.in_wire_1_1(vertical_tile_30_25_to_tile_29_25_1),
		.in_wire_1_2(vertical_tile_30_25_to_tile_29_25_2),
		.in_wire_1_3(vertical_tile_30_25_to_tile_29_25_3),
		.out_wire_2_0(horizontal_tile_29_25_to_tile_29_24_0),
		.out_wire_2_1(horizontal_tile_29_25_to_tile_29_24_1),
		.out_wire_2_2(horizontal_tile_29_25_to_tile_29_24_2),
		.out_wire_2_3(horizontal_tile_29_25_to_tile_29_24_3),
		.in_wire_2_0(horizontal_tile_29_24_to_tile_29_25_0),
		.in_wire_2_1(horizontal_tile_29_24_to_tile_29_25_1),
		.in_wire_2_2(horizontal_tile_29_24_to_tile_29_25_2),
		.in_wire_2_3(horizontal_tile_29_24_to_tile_29_25_3),
		.out_wire_0_0(horizontal_tile_29_25_to_tile_29_26_0),
		.out_wire_0_1(horizontal_tile_29_25_to_tile_29_26_1),
		.out_wire_0_2(horizontal_tile_29_25_to_tile_29_26_2),
		.out_wire_0_3(horizontal_tile_29_25_to_tile_29_26_3),
		.in_wire_0_0(horizontal_tile_29_26_to_tile_29_25_0),
		.in_wire_0_1(horizontal_tile_29_26_to_tile_29_25_1),
		.in_wire_0_2(horizontal_tile_29_26_to_tile_29_25_2),
		.in_wire_0_3(horizontal_tile_29_26_to_tile_29_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(954)
	);

	pe_tile pe_tile_29_26(
		.out_wire_3_0(vertical_tile_29_26_to_tile_28_26_0),
		.out_wire_3_1(vertical_tile_29_26_to_tile_28_26_1),
		.out_wire_3_2(vertical_tile_29_26_to_tile_28_26_2),
		.out_wire_3_3(vertical_tile_29_26_to_tile_28_26_3),
		.in_wire_3_0(vertical_tile_28_26_to_tile_29_26_0),
		.in_wire_3_1(vertical_tile_28_26_to_tile_29_26_1),
		.in_wire_3_2(vertical_tile_28_26_to_tile_29_26_2),
		.in_wire_3_3(vertical_tile_28_26_to_tile_29_26_3),
		.out_wire_1_0(vertical_tile_29_26_to_tile_30_26_0),
		.out_wire_1_1(vertical_tile_29_26_to_tile_30_26_1),
		.out_wire_1_2(vertical_tile_29_26_to_tile_30_26_2),
		.out_wire_1_3(vertical_tile_29_26_to_tile_30_26_3),
		.in_wire_1_0(vertical_tile_30_26_to_tile_29_26_0),
		.in_wire_1_1(vertical_tile_30_26_to_tile_29_26_1),
		.in_wire_1_2(vertical_tile_30_26_to_tile_29_26_2),
		.in_wire_1_3(vertical_tile_30_26_to_tile_29_26_3),
		.out_wire_2_0(horizontal_tile_29_26_to_tile_29_25_0),
		.out_wire_2_1(horizontal_tile_29_26_to_tile_29_25_1),
		.out_wire_2_2(horizontal_tile_29_26_to_tile_29_25_2),
		.out_wire_2_3(horizontal_tile_29_26_to_tile_29_25_3),
		.in_wire_2_0(horizontal_tile_29_25_to_tile_29_26_0),
		.in_wire_2_1(horizontal_tile_29_25_to_tile_29_26_1),
		.in_wire_2_2(horizontal_tile_29_25_to_tile_29_26_2),
		.in_wire_2_3(horizontal_tile_29_25_to_tile_29_26_3),
		.out_wire_0_0(horizontal_tile_29_26_to_tile_29_27_0),
		.out_wire_0_1(horizontal_tile_29_26_to_tile_29_27_1),
		.out_wire_0_2(horizontal_tile_29_26_to_tile_29_27_2),
		.out_wire_0_3(horizontal_tile_29_26_to_tile_29_27_3),
		.in_wire_0_0(horizontal_tile_29_27_to_tile_29_26_0),
		.in_wire_0_1(horizontal_tile_29_27_to_tile_29_26_1),
		.in_wire_0_2(horizontal_tile_29_27_to_tile_29_26_2),
		.in_wire_0_3(horizontal_tile_29_27_to_tile_29_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(955)
	);

	pe_tile pe_tile_29_27(
		.out_wire_3_0(vertical_tile_29_27_to_tile_28_27_0),
		.out_wire_3_1(vertical_tile_29_27_to_tile_28_27_1),
		.out_wire_3_2(vertical_tile_29_27_to_tile_28_27_2),
		.out_wire_3_3(vertical_tile_29_27_to_tile_28_27_3),
		.in_wire_3_0(vertical_tile_28_27_to_tile_29_27_0),
		.in_wire_3_1(vertical_tile_28_27_to_tile_29_27_1),
		.in_wire_3_2(vertical_tile_28_27_to_tile_29_27_2),
		.in_wire_3_3(vertical_tile_28_27_to_tile_29_27_3),
		.out_wire_1_0(vertical_tile_29_27_to_tile_30_27_0),
		.out_wire_1_1(vertical_tile_29_27_to_tile_30_27_1),
		.out_wire_1_2(vertical_tile_29_27_to_tile_30_27_2),
		.out_wire_1_3(vertical_tile_29_27_to_tile_30_27_3),
		.in_wire_1_0(vertical_tile_30_27_to_tile_29_27_0),
		.in_wire_1_1(vertical_tile_30_27_to_tile_29_27_1),
		.in_wire_1_2(vertical_tile_30_27_to_tile_29_27_2),
		.in_wire_1_3(vertical_tile_30_27_to_tile_29_27_3),
		.out_wire_2_0(horizontal_tile_29_27_to_tile_29_26_0),
		.out_wire_2_1(horizontal_tile_29_27_to_tile_29_26_1),
		.out_wire_2_2(horizontal_tile_29_27_to_tile_29_26_2),
		.out_wire_2_3(horizontal_tile_29_27_to_tile_29_26_3),
		.in_wire_2_0(horizontal_tile_29_26_to_tile_29_27_0),
		.in_wire_2_1(horizontal_tile_29_26_to_tile_29_27_1),
		.in_wire_2_2(horizontal_tile_29_26_to_tile_29_27_2),
		.in_wire_2_3(horizontal_tile_29_26_to_tile_29_27_3),
		.out_wire_0_0(horizontal_tile_29_27_to_tile_29_28_0),
		.out_wire_0_1(horizontal_tile_29_27_to_tile_29_28_1),
		.out_wire_0_2(horizontal_tile_29_27_to_tile_29_28_2),
		.out_wire_0_3(horizontal_tile_29_27_to_tile_29_28_3),
		.in_wire_0_0(horizontal_tile_29_28_to_tile_29_27_0),
		.in_wire_0_1(horizontal_tile_29_28_to_tile_29_27_1),
		.in_wire_0_2(horizontal_tile_29_28_to_tile_29_27_2),
		.in_wire_0_3(horizontal_tile_29_28_to_tile_29_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(956)
	);

	pe_tile pe_tile_29_28(
		.out_wire_3_0(vertical_tile_29_28_to_tile_28_28_0),
		.out_wire_3_1(vertical_tile_29_28_to_tile_28_28_1),
		.out_wire_3_2(vertical_tile_29_28_to_tile_28_28_2),
		.out_wire_3_3(vertical_tile_29_28_to_tile_28_28_3),
		.in_wire_3_0(vertical_tile_28_28_to_tile_29_28_0),
		.in_wire_3_1(vertical_tile_28_28_to_tile_29_28_1),
		.in_wire_3_2(vertical_tile_28_28_to_tile_29_28_2),
		.in_wire_3_3(vertical_tile_28_28_to_tile_29_28_3),
		.out_wire_1_0(vertical_tile_29_28_to_tile_30_28_0),
		.out_wire_1_1(vertical_tile_29_28_to_tile_30_28_1),
		.out_wire_1_2(vertical_tile_29_28_to_tile_30_28_2),
		.out_wire_1_3(vertical_tile_29_28_to_tile_30_28_3),
		.in_wire_1_0(vertical_tile_30_28_to_tile_29_28_0),
		.in_wire_1_1(vertical_tile_30_28_to_tile_29_28_1),
		.in_wire_1_2(vertical_tile_30_28_to_tile_29_28_2),
		.in_wire_1_3(vertical_tile_30_28_to_tile_29_28_3),
		.out_wire_2_0(horizontal_tile_29_28_to_tile_29_27_0),
		.out_wire_2_1(horizontal_tile_29_28_to_tile_29_27_1),
		.out_wire_2_2(horizontal_tile_29_28_to_tile_29_27_2),
		.out_wire_2_3(horizontal_tile_29_28_to_tile_29_27_3),
		.in_wire_2_0(horizontal_tile_29_27_to_tile_29_28_0),
		.in_wire_2_1(horizontal_tile_29_27_to_tile_29_28_1),
		.in_wire_2_2(horizontal_tile_29_27_to_tile_29_28_2),
		.in_wire_2_3(horizontal_tile_29_27_to_tile_29_28_3),
		.out_wire_0_0(horizontal_tile_29_28_to_tile_29_29_0),
		.out_wire_0_1(horizontal_tile_29_28_to_tile_29_29_1),
		.out_wire_0_2(horizontal_tile_29_28_to_tile_29_29_2),
		.out_wire_0_3(horizontal_tile_29_28_to_tile_29_29_3),
		.in_wire_0_0(horizontal_tile_29_29_to_tile_29_28_0),
		.in_wire_0_1(horizontal_tile_29_29_to_tile_29_28_1),
		.in_wire_0_2(horizontal_tile_29_29_to_tile_29_28_2),
		.in_wire_0_3(horizontal_tile_29_29_to_tile_29_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(957)
	);

	pe_tile pe_tile_29_29(
		.out_wire_3_0(vertical_tile_29_29_to_tile_28_29_0),
		.out_wire_3_1(vertical_tile_29_29_to_tile_28_29_1),
		.out_wire_3_2(vertical_tile_29_29_to_tile_28_29_2),
		.out_wire_3_3(vertical_tile_29_29_to_tile_28_29_3),
		.in_wire_3_0(vertical_tile_28_29_to_tile_29_29_0),
		.in_wire_3_1(vertical_tile_28_29_to_tile_29_29_1),
		.in_wire_3_2(vertical_tile_28_29_to_tile_29_29_2),
		.in_wire_3_3(vertical_tile_28_29_to_tile_29_29_3),
		.out_wire_1_0(vertical_tile_29_29_to_tile_30_29_0),
		.out_wire_1_1(vertical_tile_29_29_to_tile_30_29_1),
		.out_wire_1_2(vertical_tile_29_29_to_tile_30_29_2),
		.out_wire_1_3(vertical_tile_29_29_to_tile_30_29_3),
		.in_wire_1_0(vertical_tile_30_29_to_tile_29_29_0),
		.in_wire_1_1(vertical_tile_30_29_to_tile_29_29_1),
		.in_wire_1_2(vertical_tile_30_29_to_tile_29_29_2),
		.in_wire_1_3(vertical_tile_30_29_to_tile_29_29_3),
		.out_wire_2_0(horizontal_tile_29_29_to_tile_29_28_0),
		.out_wire_2_1(horizontal_tile_29_29_to_tile_29_28_1),
		.out_wire_2_2(horizontal_tile_29_29_to_tile_29_28_2),
		.out_wire_2_3(horizontal_tile_29_29_to_tile_29_28_3),
		.in_wire_2_0(horizontal_tile_29_28_to_tile_29_29_0),
		.in_wire_2_1(horizontal_tile_29_28_to_tile_29_29_1),
		.in_wire_2_2(horizontal_tile_29_28_to_tile_29_29_2),
		.in_wire_2_3(horizontal_tile_29_28_to_tile_29_29_3),
		.out_wire_0_0(horizontal_tile_29_29_to_tile_29_30_0),
		.out_wire_0_1(horizontal_tile_29_29_to_tile_29_30_1),
		.out_wire_0_2(horizontal_tile_29_29_to_tile_29_30_2),
		.out_wire_0_3(horizontal_tile_29_29_to_tile_29_30_3),
		.in_wire_0_0(horizontal_tile_29_30_to_tile_29_29_0),
		.in_wire_0_1(horizontal_tile_29_30_to_tile_29_29_1),
		.in_wire_0_2(horizontal_tile_29_30_to_tile_29_29_2),
		.in_wire_0_3(horizontal_tile_29_30_to_tile_29_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(958)
	);

	pe_tile pe_tile_29_30(
		.out_wire_3_0(vertical_tile_29_30_to_tile_28_30_0),
		.out_wire_3_1(vertical_tile_29_30_to_tile_28_30_1),
		.out_wire_3_2(vertical_tile_29_30_to_tile_28_30_2),
		.out_wire_3_3(vertical_tile_29_30_to_tile_28_30_3),
		.in_wire_3_0(vertical_tile_28_30_to_tile_29_30_0),
		.in_wire_3_1(vertical_tile_28_30_to_tile_29_30_1),
		.in_wire_3_2(vertical_tile_28_30_to_tile_29_30_2),
		.in_wire_3_3(vertical_tile_28_30_to_tile_29_30_3),
		.out_wire_1_0(vertical_tile_29_30_to_tile_30_30_0),
		.out_wire_1_1(vertical_tile_29_30_to_tile_30_30_1),
		.out_wire_1_2(vertical_tile_29_30_to_tile_30_30_2),
		.out_wire_1_3(vertical_tile_29_30_to_tile_30_30_3),
		.in_wire_1_0(vertical_tile_30_30_to_tile_29_30_0),
		.in_wire_1_1(vertical_tile_30_30_to_tile_29_30_1),
		.in_wire_1_2(vertical_tile_30_30_to_tile_29_30_2),
		.in_wire_1_3(vertical_tile_30_30_to_tile_29_30_3),
		.out_wire_2_0(horizontal_tile_29_30_to_tile_29_29_0),
		.out_wire_2_1(horizontal_tile_29_30_to_tile_29_29_1),
		.out_wire_2_2(horizontal_tile_29_30_to_tile_29_29_2),
		.out_wire_2_3(horizontal_tile_29_30_to_tile_29_29_3),
		.in_wire_2_0(horizontal_tile_29_29_to_tile_29_30_0),
		.in_wire_2_1(horizontal_tile_29_29_to_tile_29_30_1),
		.in_wire_2_2(horizontal_tile_29_29_to_tile_29_30_2),
		.in_wire_2_3(horizontal_tile_29_29_to_tile_29_30_3),
		.out_wire_0_0(horizontal_tile_29_30_to_tile_29_31_0),
		.out_wire_0_1(horizontal_tile_29_30_to_tile_29_31_1),
		.out_wire_0_2(horizontal_tile_29_30_to_tile_29_31_2),
		.out_wire_0_3(horizontal_tile_29_30_to_tile_29_31_3),
		.in_wire_0_0(horizontal_tile_29_31_to_tile_29_30_0),
		.in_wire_0_1(horizontal_tile_29_31_to_tile_29_30_1),
		.in_wire_0_2(horizontal_tile_29_31_to_tile_29_30_2),
		.in_wire_0_3(horizontal_tile_29_31_to_tile_29_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(959)
	);

	pe_tile_right pe_tile_29_31(
		.out_wire_3_0(vertical_tile_29_31_to_tile_28_31_0),
		.out_wire_3_1(vertical_tile_29_31_to_tile_28_31_1),
		.out_wire_3_2(vertical_tile_29_31_to_tile_28_31_2),
		.out_wire_3_3(vertical_tile_29_31_to_tile_28_31_3),
		.in_wire_3_0(vertical_tile_28_31_to_tile_29_31_0),
		.in_wire_3_1(vertical_tile_28_31_to_tile_29_31_1),
		.in_wire_3_2(vertical_tile_28_31_to_tile_29_31_2),
		.in_wire_3_3(vertical_tile_28_31_to_tile_29_31_3),
		.out_wire_1_0(vertical_tile_29_31_to_tile_30_31_0),
		.out_wire_1_1(vertical_tile_29_31_to_tile_30_31_1),
		.out_wire_1_2(vertical_tile_29_31_to_tile_30_31_2),
		.out_wire_1_3(vertical_tile_29_31_to_tile_30_31_3),
		.in_wire_1_0(vertical_tile_30_31_to_tile_29_31_0),
		.in_wire_1_1(vertical_tile_30_31_to_tile_29_31_1),
		.in_wire_1_2(vertical_tile_30_31_to_tile_29_31_2),
		.in_wire_1_3(vertical_tile_30_31_to_tile_29_31_3),
		.out_wire_2_0(horizontal_tile_29_31_to_tile_29_30_0),
		.out_wire_2_1(horizontal_tile_29_31_to_tile_29_30_1),
		.out_wire_2_2(horizontal_tile_29_31_to_tile_29_30_2),
		.out_wire_2_3(horizontal_tile_29_31_to_tile_29_30_3),
		.in_wire_2_0(horizontal_tile_29_30_to_tile_29_31_0),
		.in_wire_2_1(horizontal_tile_29_30_to_tile_29_31_1),
		.in_wire_2_2(horizontal_tile_29_30_to_tile_29_31_2),
		.in_wire_2_3(horizontal_tile_29_30_to_tile_29_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(960)
	);

	pe_tile_left pe_tile_30_0(
		.out_wire_3_0(vertical_tile_30_0_to_tile_29_0_0),
		.out_wire_3_1(vertical_tile_30_0_to_tile_29_0_1),
		.out_wire_3_2(vertical_tile_30_0_to_tile_29_0_2),
		.out_wire_3_3(vertical_tile_30_0_to_tile_29_0_3),
		.in_wire_3_0(vertical_tile_29_0_to_tile_30_0_0),
		.in_wire_3_1(vertical_tile_29_0_to_tile_30_0_1),
		.in_wire_3_2(vertical_tile_29_0_to_tile_30_0_2),
		.in_wire_3_3(vertical_tile_29_0_to_tile_30_0_3),
		.out_wire_1_0(vertical_tile_30_0_to_tile_31_0_0),
		.out_wire_1_1(vertical_tile_30_0_to_tile_31_0_1),
		.out_wire_1_2(vertical_tile_30_0_to_tile_31_0_2),
		.out_wire_1_3(vertical_tile_30_0_to_tile_31_0_3),
		.in_wire_1_0(vertical_tile_31_0_to_tile_30_0_0),
		.in_wire_1_1(vertical_tile_31_0_to_tile_30_0_1),
		.in_wire_1_2(vertical_tile_31_0_to_tile_30_0_2),
		.in_wire_1_3(vertical_tile_31_0_to_tile_30_0_3),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_30_0_to_tile_30_1_0),
		.out_wire_0_1(horizontal_tile_30_0_to_tile_30_1_1),
		.out_wire_0_2(horizontal_tile_30_0_to_tile_30_1_2),
		.out_wire_0_3(horizontal_tile_30_0_to_tile_30_1_3),
		.in_wire_0_0(horizontal_tile_30_1_to_tile_30_0_0),
		.in_wire_0_1(horizontal_tile_30_1_to_tile_30_0_1),
		.in_wire_0_2(horizontal_tile_30_1_to_tile_30_0_2),
		.in_wire_0_3(horizontal_tile_30_1_to_tile_30_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(961)
	);

	pe_tile pe_tile_30_1(
		.out_wire_3_0(vertical_tile_30_1_to_tile_29_1_0),
		.out_wire_3_1(vertical_tile_30_1_to_tile_29_1_1),
		.out_wire_3_2(vertical_tile_30_1_to_tile_29_1_2),
		.out_wire_3_3(vertical_tile_30_1_to_tile_29_1_3),
		.in_wire_3_0(vertical_tile_29_1_to_tile_30_1_0),
		.in_wire_3_1(vertical_tile_29_1_to_tile_30_1_1),
		.in_wire_3_2(vertical_tile_29_1_to_tile_30_1_2),
		.in_wire_3_3(vertical_tile_29_1_to_tile_30_1_3),
		.out_wire_1_0(vertical_tile_30_1_to_tile_31_1_0),
		.out_wire_1_1(vertical_tile_30_1_to_tile_31_1_1),
		.out_wire_1_2(vertical_tile_30_1_to_tile_31_1_2),
		.out_wire_1_3(vertical_tile_30_1_to_tile_31_1_3),
		.in_wire_1_0(vertical_tile_31_1_to_tile_30_1_0),
		.in_wire_1_1(vertical_tile_31_1_to_tile_30_1_1),
		.in_wire_1_2(vertical_tile_31_1_to_tile_30_1_2),
		.in_wire_1_3(vertical_tile_31_1_to_tile_30_1_3),
		.out_wire_2_0(horizontal_tile_30_1_to_tile_30_0_0),
		.out_wire_2_1(horizontal_tile_30_1_to_tile_30_0_1),
		.out_wire_2_2(horizontal_tile_30_1_to_tile_30_0_2),
		.out_wire_2_3(horizontal_tile_30_1_to_tile_30_0_3),
		.in_wire_2_0(horizontal_tile_30_0_to_tile_30_1_0),
		.in_wire_2_1(horizontal_tile_30_0_to_tile_30_1_1),
		.in_wire_2_2(horizontal_tile_30_0_to_tile_30_1_2),
		.in_wire_2_3(horizontal_tile_30_0_to_tile_30_1_3),
		.out_wire_0_0(horizontal_tile_30_1_to_tile_30_2_0),
		.out_wire_0_1(horizontal_tile_30_1_to_tile_30_2_1),
		.out_wire_0_2(horizontal_tile_30_1_to_tile_30_2_2),
		.out_wire_0_3(horizontal_tile_30_1_to_tile_30_2_3),
		.in_wire_0_0(horizontal_tile_30_2_to_tile_30_1_0),
		.in_wire_0_1(horizontal_tile_30_2_to_tile_30_1_1),
		.in_wire_0_2(horizontal_tile_30_2_to_tile_30_1_2),
		.in_wire_0_3(horizontal_tile_30_2_to_tile_30_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(962)
	);

	pe_tile pe_tile_30_2(
		.out_wire_3_0(vertical_tile_30_2_to_tile_29_2_0),
		.out_wire_3_1(vertical_tile_30_2_to_tile_29_2_1),
		.out_wire_3_2(vertical_tile_30_2_to_tile_29_2_2),
		.out_wire_3_3(vertical_tile_30_2_to_tile_29_2_3),
		.in_wire_3_0(vertical_tile_29_2_to_tile_30_2_0),
		.in_wire_3_1(vertical_tile_29_2_to_tile_30_2_1),
		.in_wire_3_2(vertical_tile_29_2_to_tile_30_2_2),
		.in_wire_3_3(vertical_tile_29_2_to_tile_30_2_3),
		.out_wire_1_0(vertical_tile_30_2_to_tile_31_2_0),
		.out_wire_1_1(vertical_tile_30_2_to_tile_31_2_1),
		.out_wire_1_2(vertical_tile_30_2_to_tile_31_2_2),
		.out_wire_1_3(vertical_tile_30_2_to_tile_31_2_3),
		.in_wire_1_0(vertical_tile_31_2_to_tile_30_2_0),
		.in_wire_1_1(vertical_tile_31_2_to_tile_30_2_1),
		.in_wire_1_2(vertical_tile_31_2_to_tile_30_2_2),
		.in_wire_1_3(vertical_tile_31_2_to_tile_30_2_3),
		.out_wire_2_0(horizontal_tile_30_2_to_tile_30_1_0),
		.out_wire_2_1(horizontal_tile_30_2_to_tile_30_1_1),
		.out_wire_2_2(horizontal_tile_30_2_to_tile_30_1_2),
		.out_wire_2_3(horizontal_tile_30_2_to_tile_30_1_3),
		.in_wire_2_0(horizontal_tile_30_1_to_tile_30_2_0),
		.in_wire_2_1(horizontal_tile_30_1_to_tile_30_2_1),
		.in_wire_2_2(horizontal_tile_30_1_to_tile_30_2_2),
		.in_wire_2_3(horizontal_tile_30_1_to_tile_30_2_3),
		.out_wire_0_0(horizontal_tile_30_2_to_tile_30_3_0),
		.out_wire_0_1(horizontal_tile_30_2_to_tile_30_3_1),
		.out_wire_0_2(horizontal_tile_30_2_to_tile_30_3_2),
		.out_wire_0_3(horizontal_tile_30_2_to_tile_30_3_3),
		.in_wire_0_0(horizontal_tile_30_3_to_tile_30_2_0),
		.in_wire_0_1(horizontal_tile_30_3_to_tile_30_2_1),
		.in_wire_0_2(horizontal_tile_30_3_to_tile_30_2_2),
		.in_wire_0_3(horizontal_tile_30_3_to_tile_30_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(963)
	);

	pe_tile pe_tile_30_3(
		.out_wire_3_0(vertical_tile_30_3_to_tile_29_3_0),
		.out_wire_3_1(vertical_tile_30_3_to_tile_29_3_1),
		.out_wire_3_2(vertical_tile_30_3_to_tile_29_3_2),
		.out_wire_3_3(vertical_tile_30_3_to_tile_29_3_3),
		.in_wire_3_0(vertical_tile_29_3_to_tile_30_3_0),
		.in_wire_3_1(vertical_tile_29_3_to_tile_30_3_1),
		.in_wire_3_2(vertical_tile_29_3_to_tile_30_3_2),
		.in_wire_3_3(vertical_tile_29_3_to_tile_30_3_3),
		.out_wire_1_0(vertical_tile_30_3_to_tile_31_3_0),
		.out_wire_1_1(vertical_tile_30_3_to_tile_31_3_1),
		.out_wire_1_2(vertical_tile_30_3_to_tile_31_3_2),
		.out_wire_1_3(vertical_tile_30_3_to_tile_31_3_3),
		.in_wire_1_0(vertical_tile_31_3_to_tile_30_3_0),
		.in_wire_1_1(vertical_tile_31_3_to_tile_30_3_1),
		.in_wire_1_2(vertical_tile_31_3_to_tile_30_3_2),
		.in_wire_1_3(vertical_tile_31_3_to_tile_30_3_3),
		.out_wire_2_0(horizontal_tile_30_3_to_tile_30_2_0),
		.out_wire_2_1(horizontal_tile_30_3_to_tile_30_2_1),
		.out_wire_2_2(horizontal_tile_30_3_to_tile_30_2_2),
		.out_wire_2_3(horizontal_tile_30_3_to_tile_30_2_3),
		.in_wire_2_0(horizontal_tile_30_2_to_tile_30_3_0),
		.in_wire_2_1(horizontal_tile_30_2_to_tile_30_3_1),
		.in_wire_2_2(horizontal_tile_30_2_to_tile_30_3_2),
		.in_wire_2_3(horizontal_tile_30_2_to_tile_30_3_3),
		.out_wire_0_0(horizontal_tile_30_3_to_tile_30_4_0),
		.out_wire_0_1(horizontal_tile_30_3_to_tile_30_4_1),
		.out_wire_0_2(horizontal_tile_30_3_to_tile_30_4_2),
		.out_wire_0_3(horizontal_tile_30_3_to_tile_30_4_3),
		.in_wire_0_0(horizontal_tile_30_4_to_tile_30_3_0),
		.in_wire_0_1(horizontal_tile_30_4_to_tile_30_3_1),
		.in_wire_0_2(horizontal_tile_30_4_to_tile_30_3_2),
		.in_wire_0_3(horizontal_tile_30_4_to_tile_30_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(964)
	);

	pe_tile pe_tile_30_4(
		.out_wire_3_0(vertical_tile_30_4_to_tile_29_4_0),
		.out_wire_3_1(vertical_tile_30_4_to_tile_29_4_1),
		.out_wire_3_2(vertical_tile_30_4_to_tile_29_4_2),
		.out_wire_3_3(vertical_tile_30_4_to_tile_29_4_3),
		.in_wire_3_0(vertical_tile_29_4_to_tile_30_4_0),
		.in_wire_3_1(vertical_tile_29_4_to_tile_30_4_1),
		.in_wire_3_2(vertical_tile_29_4_to_tile_30_4_2),
		.in_wire_3_3(vertical_tile_29_4_to_tile_30_4_3),
		.out_wire_1_0(vertical_tile_30_4_to_tile_31_4_0),
		.out_wire_1_1(vertical_tile_30_4_to_tile_31_4_1),
		.out_wire_1_2(vertical_tile_30_4_to_tile_31_4_2),
		.out_wire_1_3(vertical_tile_30_4_to_tile_31_4_3),
		.in_wire_1_0(vertical_tile_31_4_to_tile_30_4_0),
		.in_wire_1_1(vertical_tile_31_4_to_tile_30_4_1),
		.in_wire_1_2(vertical_tile_31_4_to_tile_30_4_2),
		.in_wire_1_3(vertical_tile_31_4_to_tile_30_4_3),
		.out_wire_2_0(horizontal_tile_30_4_to_tile_30_3_0),
		.out_wire_2_1(horizontal_tile_30_4_to_tile_30_3_1),
		.out_wire_2_2(horizontal_tile_30_4_to_tile_30_3_2),
		.out_wire_2_3(horizontal_tile_30_4_to_tile_30_3_3),
		.in_wire_2_0(horizontal_tile_30_3_to_tile_30_4_0),
		.in_wire_2_1(horizontal_tile_30_3_to_tile_30_4_1),
		.in_wire_2_2(horizontal_tile_30_3_to_tile_30_4_2),
		.in_wire_2_3(horizontal_tile_30_3_to_tile_30_4_3),
		.out_wire_0_0(horizontal_tile_30_4_to_tile_30_5_0),
		.out_wire_0_1(horizontal_tile_30_4_to_tile_30_5_1),
		.out_wire_0_2(horizontal_tile_30_4_to_tile_30_5_2),
		.out_wire_0_3(horizontal_tile_30_4_to_tile_30_5_3),
		.in_wire_0_0(horizontal_tile_30_5_to_tile_30_4_0),
		.in_wire_0_1(horizontal_tile_30_5_to_tile_30_4_1),
		.in_wire_0_2(horizontal_tile_30_5_to_tile_30_4_2),
		.in_wire_0_3(horizontal_tile_30_5_to_tile_30_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(965)
	);

	pe_tile pe_tile_30_5(
		.out_wire_3_0(vertical_tile_30_5_to_tile_29_5_0),
		.out_wire_3_1(vertical_tile_30_5_to_tile_29_5_1),
		.out_wire_3_2(vertical_tile_30_5_to_tile_29_5_2),
		.out_wire_3_3(vertical_tile_30_5_to_tile_29_5_3),
		.in_wire_3_0(vertical_tile_29_5_to_tile_30_5_0),
		.in_wire_3_1(vertical_tile_29_5_to_tile_30_5_1),
		.in_wire_3_2(vertical_tile_29_5_to_tile_30_5_2),
		.in_wire_3_3(vertical_tile_29_5_to_tile_30_5_3),
		.out_wire_1_0(vertical_tile_30_5_to_tile_31_5_0),
		.out_wire_1_1(vertical_tile_30_5_to_tile_31_5_1),
		.out_wire_1_2(vertical_tile_30_5_to_tile_31_5_2),
		.out_wire_1_3(vertical_tile_30_5_to_tile_31_5_3),
		.in_wire_1_0(vertical_tile_31_5_to_tile_30_5_0),
		.in_wire_1_1(vertical_tile_31_5_to_tile_30_5_1),
		.in_wire_1_2(vertical_tile_31_5_to_tile_30_5_2),
		.in_wire_1_3(vertical_tile_31_5_to_tile_30_5_3),
		.out_wire_2_0(horizontal_tile_30_5_to_tile_30_4_0),
		.out_wire_2_1(horizontal_tile_30_5_to_tile_30_4_1),
		.out_wire_2_2(horizontal_tile_30_5_to_tile_30_4_2),
		.out_wire_2_3(horizontal_tile_30_5_to_tile_30_4_3),
		.in_wire_2_0(horizontal_tile_30_4_to_tile_30_5_0),
		.in_wire_2_1(horizontal_tile_30_4_to_tile_30_5_1),
		.in_wire_2_2(horizontal_tile_30_4_to_tile_30_5_2),
		.in_wire_2_3(horizontal_tile_30_4_to_tile_30_5_3),
		.out_wire_0_0(horizontal_tile_30_5_to_tile_30_6_0),
		.out_wire_0_1(horizontal_tile_30_5_to_tile_30_6_1),
		.out_wire_0_2(horizontal_tile_30_5_to_tile_30_6_2),
		.out_wire_0_3(horizontal_tile_30_5_to_tile_30_6_3),
		.in_wire_0_0(horizontal_tile_30_6_to_tile_30_5_0),
		.in_wire_0_1(horizontal_tile_30_6_to_tile_30_5_1),
		.in_wire_0_2(horizontal_tile_30_6_to_tile_30_5_2),
		.in_wire_0_3(horizontal_tile_30_6_to_tile_30_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(966)
	);

	pe_tile pe_tile_30_6(
		.out_wire_3_0(vertical_tile_30_6_to_tile_29_6_0),
		.out_wire_3_1(vertical_tile_30_6_to_tile_29_6_1),
		.out_wire_3_2(vertical_tile_30_6_to_tile_29_6_2),
		.out_wire_3_3(vertical_tile_30_6_to_tile_29_6_3),
		.in_wire_3_0(vertical_tile_29_6_to_tile_30_6_0),
		.in_wire_3_1(vertical_tile_29_6_to_tile_30_6_1),
		.in_wire_3_2(vertical_tile_29_6_to_tile_30_6_2),
		.in_wire_3_3(vertical_tile_29_6_to_tile_30_6_3),
		.out_wire_1_0(vertical_tile_30_6_to_tile_31_6_0),
		.out_wire_1_1(vertical_tile_30_6_to_tile_31_6_1),
		.out_wire_1_2(vertical_tile_30_6_to_tile_31_6_2),
		.out_wire_1_3(vertical_tile_30_6_to_tile_31_6_3),
		.in_wire_1_0(vertical_tile_31_6_to_tile_30_6_0),
		.in_wire_1_1(vertical_tile_31_6_to_tile_30_6_1),
		.in_wire_1_2(vertical_tile_31_6_to_tile_30_6_2),
		.in_wire_1_3(vertical_tile_31_6_to_tile_30_6_3),
		.out_wire_2_0(horizontal_tile_30_6_to_tile_30_5_0),
		.out_wire_2_1(horizontal_tile_30_6_to_tile_30_5_1),
		.out_wire_2_2(horizontal_tile_30_6_to_tile_30_5_2),
		.out_wire_2_3(horizontal_tile_30_6_to_tile_30_5_3),
		.in_wire_2_0(horizontal_tile_30_5_to_tile_30_6_0),
		.in_wire_2_1(horizontal_tile_30_5_to_tile_30_6_1),
		.in_wire_2_2(horizontal_tile_30_5_to_tile_30_6_2),
		.in_wire_2_3(horizontal_tile_30_5_to_tile_30_6_3),
		.out_wire_0_0(horizontal_tile_30_6_to_tile_30_7_0),
		.out_wire_0_1(horizontal_tile_30_6_to_tile_30_7_1),
		.out_wire_0_2(horizontal_tile_30_6_to_tile_30_7_2),
		.out_wire_0_3(horizontal_tile_30_6_to_tile_30_7_3),
		.in_wire_0_0(horizontal_tile_30_7_to_tile_30_6_0),
		.in_wire_0_1(horizontal_tile_30_7_to_tile_30_6_1),
		.in_wire_0_2(horizontal_tile_30_7_to_tile_30_6_2),
		.in_wire_0_3(horizontal_tile_30_7_to_tile_30_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(967)
	);

	pe_tile pe_tile_30_7(
		.out_wire_3_0(vertical_tile_30_7_to_tile_29_7_0),
		.out_wire_3_1(vertical_tile_30_7_to_tile_29_7_1),
		.out_wire_3_2(vertical_tile_30_7_to_tile_29_7_2),
		.out_wire_3_3(vertical_tile_30_7_to_tile_29_7_3),
		.in_wire_3_0(vertical_tile_29_7_to_tile_30_7_0),
		.in_wire_3_1(vertical_tile_29_7_to_tile_30_7_1),
		.in_wire_3_2(vertical_tile_29_7_to_tile_30_7_2),
		.in_wire_3_3(vertical_tile_29_7_to_tile_30_7_3),
		.out_wire_1_0(vertical_tile_30_7_to_tile_31_7_0),
		.out_wire_1_1(vertical_tile_30_7_to_tile_31_7_1),
		.out_wire_1_2(vertical_tile_30_7_to_tile_31_7_2),
		.out_wire_1_3(vertical_tile_30_7_to_tile_31_7_3),
		.in_wire_1_0(vertical_tile_31_7_to_tile_30_7_0),
		.in_wire_1_1(vertical_tile_31_7_to_tile_30_7_1),
		.in_wire_1_2(vertical_tile_31_7_to_tile_30_7_2),
		.in_wire_1_3(vertical_tile_31_7_to_tile_30_7_3),
		.out_wire_2_0(horizontal_tile_30_7_to_tile_30_6_0),
		.out_wire_2_1(horizontal_tile_30_7_to_tile_30_6_1),
		.out_wire_2_2(horizontal_tile_30_7_to_tile_30_6_2),
		.out_wire_2_3(horizontal_tile_30_7_to_tile_30_6_3),
		.in_wire_2_0(horizontal_tile_30_6_to_tile_30_7_0),
		.in_wire_2_1(horizontal_tile_30_6_to_tile_30_7_1),
		.in_wire_2_2(horizontal_tile_30_6_to_tile_30_7_2),
		.in_wire_2_3(horizontal_tile_30_6_to_tile_30_7_3),
		.out_wire_0_0(horizontal_tile_30_7_to_tile_30_8_0),
		.out_wire_0_1(horizontal_tile_30_7_to_tile_30_8_1),
		.out_wire_0_2(horizontal_tile_30_7_to_tile_30_8_2),
		.out_wire_0_3(horizontal_tile_30_7_to_tile_30_8_3),
		.in_wire_0_0(horizontal_tile_30_8_to_tile_30_7_0),
		.in_wire_0_1(horizontal_tile_30_8_to_tile_30_7_1),
		.in_wire_0_2(horizontal_tile_30_8_to_tile_30_7_2),
		.in_wire_0_3(horizontal_tile_30_8_to_tile_30_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(968)
	);

	pe_tile pe_tile_30_8(
		.out_wire_3_0(vertical_tile_30_8_to_tile_29_8_0),
		.out_wire_3_1(vertical_tile_30_8_to_tile_29_8_1),
		.out_wire_3_2(vertical_tile_30_8_to_tile_29_8_2),
		.out_wire_3_3(vertical_tile_30_8_to_tile_29_8_3),
		.in_wire_3_0(vertical_tile_29_8_to_tile_30_8_0),
		.in_wire_3_1(vertical_tile_29_8_to_tile_30_8_1),
		.in_wire_3_2(vertical_tile_29_8_to_tile_30_8_2),
		.in_wire_3_3(vertical_tile_29_8_to_tile_30_8_3),
		.out_wire_1_0(vertical_tile_30_8_to_tile_31_8_0),
		.out_wire_1_1(vertical_tile_30_8_to_tile_31_8_1),
		.out_wire_1_2(vertical_tile_30_8_to_tile_31_8_2),
		.out_wire_1_3(vertical_tile_30_8_to_tile_31_8_3),
		.in_wire_1_0(vertical_tile_31_8_to_tile_30_8_0),
		.in_wire_1_1(vertical_tile_31_8_to_tile_30_8_1),
		.in_wire_1_2(vertical_tile_31_8_to_tile_30_8_2),
		.in_wire_1_3(vertical_tile_31_8_to_tile_30_8_3),
		.out_wire_2_0(horizontal_tile_30_8_to_tile_30_7_0),
		.out_wire_2_1(horizontal_tile_30_8_to_tile_30_7_1),
		.out_wire_2_2(horizontal_tile_30_8_to_tile_30_7_2),
		.out_wire_2_3(horizontal_tile_30_8_to_tile_30_7_3),
		.in_wire_2_0(horizontal_tile_30_7_to_tile_30_8_0),
		.in_wire_2_1(horizontal_tile_30_7_to_tile_30_8_1),
		.in_wire_2_2(horizontal_tile_30_7_to_tile_30_8_2),
		.in_wire_2_3(horizontal_tile_30_7_to_tile_30_8_3),
		.out_wire_0_0(horizontal_tile_30_8_to_tile_30_9_0),
		.out_wire_0_1(horizontal_tile_30_8_to_tile_30_9_1),
		.out_wire_0_2(horizontal_tile_30_8_to_tile_30_9_2),
		.out_wire_0_3(horizontal_tile_30_8_to_tile_30_9_3),
		.in_wire_0_0(horizontal_tile_30_9_to_tile_30_8_0),
		.in_wire_0_1(horizontal_tile_30_9_to_tile_30_8_1),
		.in_wire_0_2(horizontal_tile_30_9_to_tile_30_8_2),
		.in_wire_0_3(horizontal_tile_30_9_to_tile_30_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(969)
	);

	pe_tile pe_tile_30_9(
		.out_wire_3_0(vertical_tile_30_9_to_tile_29_9_0),
		.out_wire_3_1(vertical_tile_30_9_to_tile_29_9_1),
		.out_wire_3_2(vertical_tile_30_9_to_tile_29_9_2),
		.out_wire_3_3(vertical_tile_30_9_to_tile_29_9_3),
		.in_wire_3_0(vertical_tile_29_9_to_tile_30_9_0),
		.in_wire_3_1(vertical_tile_29_9_to_tile_30_9_1),
		.in_wire_3_2(vertical_tile_29_9_to_tile_30_9_2),
		.in_wire_3_3(vertical_tile_29_9_to_tile_30_9_3),
		.out_wire_1_0(vertical_tile_30_9_to_tile_31_9_0),
		.out_wire_1_1(vertical_tile_30_9_to_tile_31_9_1),
		.out_wire_1_2(vertical_tile_30_9_to_tile_31_9_2),
		.out_wire_1_3(vertical_tile_30_9_to_tile_31_9_3),
		.in_wire_1_0(vertical_tile_31_9_to_tile_30_9_0),
		.in_wire_1_1(vertical_tile_31_9_to_tile_30_9_1),
		.in_wire_1_2(vertical_tile_31_9_to_tile_30_9_2),
		.in_wire_1_3(vertical_tile_31_9_to_tile_30_9_3),
		.out_wire_2_0(horizontal_tile_30_9_to_tile_30_8_0),
		.out_wire_2_1(horizontal_tile_30_9_to_tile_30_8_1),
		.out_wire_2_2(horizontal_tile_30_9_to_tile_30_8_2),
		.out_wire_2_3(horizontal_tile_30_9_to_tile_30_8_3),
		.in_wire_2_0(horizontal_tile_30_8_to_tile_30_9_0),
		.in_wire_2_1(horizontal_tile_30_8_to_tile_30_9_1),
		.in_wire_2_2(horizontal_tile_30_8_to_tile_30_9_2),
		.in_wire_2_3(horizontal_tile_30_8_to_tile_30_9_3),
		.out_wire_0_0(horizontal_tile_30_9_to_tile_30_10_0),
		.out_wire_0_1(horizontal_tile_30_9_to_tile_30_10_1),
		.out_wire_0_2(horizontal_tile_30_9_to_tile_30_10_2),
		.out_wire_0_3(horizontal_tile_30_9_to_tile_30_10_3),
		.in_wire_0_0(horizontal_tile_30_10_to_tile_30_9_0),
		.in_wire_0_1(horizontal_tile_30_10_to_tile_30_9_1),
		.in_wire_0_2(horizontal_tile_30_10_to_tile_30_9_2),
		.in_wire_0_3(horizontal_tile_30_10_to_tile_30_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(970)
	);

	pe_tile pe_tile_30_10(
		.out_wire_3_0(vertical_tile_30_10_to_tile_29_10_0),
		.out_wire_3_1(vertical_tile_30_10_to_tile_29_10_1),
		.out_wire_3_2(vertical_tile_30_10_to_tile_29_10_2),
		.out_wire_3_3(vertical_tile_30_10_to_tile_29_10_3),
		.in_wire_3_0(vertical_tile_29_10_to_tile_30_10_0),
		.in_wire_3_1(vertical_tile_29_10_to_tile_30_10_1),
		.in_wire_3_2(vertical_tile_29_10_to_tile_30_10_2),
		.in_wire_3_3(vertical_tile_29_10_to_tile_30_10_3),
		.out_wire_1_0(vertical_tile_30_10_to_tile_31_10_0),
		.out_wire_1_1(vertical_tile_30_10_to_tile_31_10_1),
		.out_wire_1_2(vertical_tile_30_10_to_tile_31_10_2),
		.out_wire_1_3(vertical_tile_30_10_to_tile_31_10_3),
		.in_wire_1_0(vertical_tile_31_10_to_tile_30_10_0),
		.in_wire_1_1(vertical_tile_31_10_to_tile_30_10_1),
		.in_wire_1_2(vertical_tile_31_10_to_tile_30_10_2),
		.in_wire_1_3(vertical_tile_31_10_to_tile_30_10_3),
		.out_wire_2_0(horizontal_tile_30_10_to_tile_30_9_0),
		.out_wire_2_1(horizontal_tile_30_10_to_tile_30_9_1),
		.out_wire_2_2(horizontal_tile_30_10_to_tile_30_9_2),
		.out_wire_2_3(horizontal_tile_30_10_to_tile_30_9_3),
		.in_wire_2_0(horizontal_tile_30_9_to_tile_30_10_0),
		.in_wire_2_1(horizontal_tile_30_9_to_tile_30_10_1),
		.in_wire_2_2(horizontal_tile_30_9_to_tile_30_10_2),
		.in_wire_2_3(horizontal_tile_30_9_to_tile_30_10_3),
		.out_wire_0_0(horizontal_tile_30_10_to_tile_30_11_0),
		.out_wire_0_1(horizontal_tile_30_10_to_tile_30_11_1),
		.out_wire_0_2(horizontal_tile_30_10_to_tile_30_11_2),
		.out_wire_0_3(horizontal_tile_30_10_to_tile_30_11_3),
		.in_wire_0_0(horizontal_tile_30_11_to_tile_30_10_0),
		.in_wire_0_1(horizontal_tile_30_11_to_tile_30_10_1),
		.in_wire_0_2(horizontal_tile_30_11_to_tile_30_10_2),
		.in_wire_0_3(horizontal_tile_30_11_to_tile_30_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(971)
	);

	pe_tile pe_tile_30_11(
		.out_wire_3_0(vertical_tile_30_11_to_tile_29_11_0),
		.out_wire_3_1(vertical_tile_30_11_to_tile_29_11_1),
		.out_wire_3_2(vertical_tile_30_11_to_tile_29_11_2),
		.out_wire_3_3(vertical_tile_30_11_to_tile_29_11_3),
		.in_wire_3_0(vertical_tile_29_11_to_tile_30_11_0),
		.in_wire_3_1(vertical_tile_29_11_to_tile_30_11_1),
		.in_wire_3_2(vertical_tile_29_11_to_tile_30_11_2),
		.in_wire_3_3(vertical_tile_29_11_to_tile_30_11_3),
		.out_wire_1_0(vertical_tile_30_11_to_tile_31_11_0),
		.out_wire_1_1(vertical_tile_30_11_to_tile_31_11_1),
		.out_wire_1_2(vertical_tile_30_11_to_tile_31_11_2),
		.out_wire_1_3(vertical_tile_30_11_to_tile_31_11_3),
		.in_wire_1_0(vertical_tile_31_11_to_tile_30_11_0),
		.in_wire_1_1(vertical_tile_31_11_to_tile_30_11_1),
		.in_wire_1_2(vertical_tile_31_11_to_tile_30_11_2),
		.in_wire_1_3(vertical_tile_31_11_to_tile_30_11_3),
		.out_wire_2_0(horizontal_tile_30_11_to_tile_30_10_0),
		.out_wire_2_1(horizontal_tile_30_11_to_tile_30_10_1),
		.out_wire_2_2(horizontal_tile_30_11_to_tile_30_10_2),
		.out_wire_2_3(horizontal_tile_30_11_to_tile_30_10_3),
		.in_wire_2_0(horizontal_tile_30_10_to_tile_30_11_0),
		.in_wire_2_1(horizontal_tile_30_10_to_tile_30_11_1),
		.in_wire_2_2(horizontal_tile_30_10_to_tile_30_11_2),
		.in_wire_2_3(horizontal_tile_30_10_to_tile_30_11_3),
		.out_wire_0_0(horizontal_tile_30_11_to_tile_30_12_0),
		.out_wire_0_1(horizontal_tile_30_11_to_tile_30_12_1),
		.out_wire_0_2(horizontal_tile_30_11_to_tile_30_12_2),
		.out_wire_0_3(horizontal_tile_30_11_to_tile_30_12_3),
		.in_wire_0_0(horizontal_tile_30_12_to_tile_30_11_0),
		.in_wire_0_1(horizontal_tile_30_12_to_tile_30_11_1),
		.in_wire_0_2(horizontal_tile_30_12_to_tile_30_11_2),
		.in_wire_0_3(horizontal_tile_30_12_to_tile_30_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(972)
	);

	pe_tile pe_tile_30_12(
		.out_wire_3_0(vertical_tile_30_12_to_tile_29_12_0),
		.out_wire_3_1(vertical_tile_30_12_to_tile_29_12_1),
		.out_wire_3_2(vertical_tile_30_12_to_tile_29_12_2),
		.out_wire_3_3(vertical_tile_30_12_to_tile_29_12_3),
		.in_wire_3_0(vertical_tile_29_12_to_tile_30_12_0),
		.in_wire_3_1(vertical_tile_29_12_to_tile_30_12_1),
		.in_wire_3_2(vertical_tile_29_12_to_tile_30_12_2),
		.in_wire_3_3(vertical_tile_29_12_to_tile_30_12_3),
		.out_wire_1_0(vertical_tile_30_12_to_tile_31_12_0),
		.out_wire_1_1(vertical_tile_30_12_to_tile_31_12_1),
		.out_wire_1_2(vertical_tile_30_12_to_tile_31_12_2),
		.out_wire_1_3(vertical_tile_30_12_to_tile_31_12_3),
		.in_wire_1_0(vertical_tile_31_12_to_tile_30_12_0),
		.in_wire_1_1(vertical_tile_31_12_to_tile_30_12_1),
		.in_wire_1_2(vertical_tile_31_12_to_tile_30_12_2),
		.in_wire_1_3(vertical_tile_31_12_to_tile_30_12_3),
		.out_wire_2_0(horizontal_tile_30_12_to_tile_30_11_0),
		.out_wire_2_1(horizontal_tile_30_12_to_tile_30_11_1),
		.out_wire_2_2(horizontal_tile_30_12_to_tile_30_11_2),
		.out_wire_2_3(horizontal_tile_30_12_to_tile_30_11_3),
		.in_wire_2_0(horizontal_tile_30_11_to_tile_30_12_0),
		.in_wire_2_1(horizontal_tile_30_11_to_tile_30_12_1),
		.in_wire_2_2(horizontal_tile_30_11_to_tile_30_12_2),
		.in_wire_2_3(horizontal_tile_30_11_to_tile_30_12_3),
		.out_wire_0_0(horizontal_tile_30_12_to_tile_30_13_0),
		.out_wire_0_1(horizontal_tile_30_12_to_tile_30_13_1),
		.out_wire_0_2(horizontal_tile_30_12_to_tile_30_13_2),
		.out_wire_0_3(horizontal_tile_30_12_to_tile_30_13_3),
		.in_wire_0_0(horizontal_tile_30_13_to_tile_30_12_0),
		.in_wire_0_1(horizontal_tile_30_13_to_tile_30_12_1),
		.in_wire_0_2(horizontal_tile_30_13_to_tile_30_12_2),
		.in_wire_0_3(horizontal_tile_30_13_to_tile_30_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(973)
	);

	pe_tile pe_tile_30_13(
		.out_wire_3_0(vertical_tile_30_13_to_tile_29_13_0),
		.out_wire_3_1(vertical_tile_30_13_to_tile_29_13_1),
		.out_wire_3_2(vertical_tile_30_13_to_tile_29_13_2),
		.out_wire_3_3(vertical_tile_30_13_to_tile_29_13_3),
		.in_wire_3_0(vertical_tile_29_13_to_tile_30_13_0),
		.in_wire_3_1(vertical_tile_29_13_to_tile_30_13_1),
		.in_wire_3_2(vertical_tile_29_13_to_tile_30_13_2),
		.in_wire_3_3(vertical_tile_29_13_to_tile_30_13_3),
		.out_wire_1_0(vertical_tile_30_13_to_tile_31_13_0),
		.out_wire_1_1(vertical_tile_30_13_to_tile_31_13_1),
		.out_wire_1_2(vertical_tile_30_13_to_tile_31_13_2),
		.out_wire_1_3(vertical_tile_30_13_to_tile_31_13_3),
		.in_wire_1_0(vertical_tile_31_13_to_tile_30_13_0),
		.in_wire_1_1(vertical_tile_31_13_to_tile_30_13_1),
		.in_wire_1_2(vertical_tile_31_13_to_tile_30_13_2),
		.in_wire_1_3(vertical_tile_31_13_to_tile_30_13_3),
		.out_wire_2_0(horizontal_tile_30_13_to_tile_30_12_0),
		.out_wire_2_1(horizontal_tile_30_13_to_tile_30_12_1),
		.out_wire_2_2(horizontal_tile_30_13_to_tile_30_12_2),
		.out_wire_2_3(horizontal_tile_30_13_to_tile_30_12_3),
		.in_wire_2_0(horizontal_tile_30_12_to_tile_30_13_0),
		.in_wire_2_1(horizontal_tile_30_12_to_tile_30_13_1),
		.in_wire_2_2(horizontal_tile_30_12_to_tile_30_13_2),
		.in_wire_2_3(horizontal_tile_30_12_to_tile_30_13_3),
		.out_wire_0_0(horizontal_tile_30_13_to_tile_30_14_0),
		.out_wire_0_1(horizontal_tile_30_13_to_tile_30_14_1),
		.out_wire_0_2(horizontal_tile_30_13_to_tile_30_14_2),
		.out_wire_0_3(horizontal_tile_30_13_to_tile_30_14_3),
		.in_wire_0_0(horizontal_tile_30_14_to_tile_30_13_0),
		.in_wire_0_1(horizontal_tile_30_14_to_tile_30_13_1),
		.in_wire_0_2(horizontal_tile_30_14_to_tile_30_13_2),
		.in_wire_0_3(horizontal_tile_30_14_to_tile_30_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(974)
	);

	pe_tile pe_tile_30_14(
		.out_wire_3_0(vertical_tile_30_14_to_tile_29_14_0),
		.out_wire_3_1(vertical_tile_30_14_to_tile_29_14_1),
		.out_wire_3_2(vertical_tile_30_14_to_tile_29_14_2),
		.out_wire_3_3(vertical_tile_30_14_to_tile_29_14_3),
		.in_wire_3_0(vertical_tile_29_14_to_tile_30_14_0),
		.in_wire_3_1(vertical_tile_29_14_to_tile_30_14_1),
		.in_wire_3_2(vertical_tile_29_14_to_tile_30_14_2),
		.in_wire_3_3(vertical_tile_29_14_to_tile_30_14_3),
		.out_wire_1_0(vertical_tile_30_14_to_tile_31_14_0),
		.out_wire_1_1(vertical_tile_30_14_to_tile_31_14_1),
		.out_wire_1_2(vertical_tile_30_14_to_tile_31_14_2),
		.out_wire_1_3(vertical_tile_30_14_to_tile_31_14_3),
		.in_wire_1_0(vertical_tile_31_14_to_tile_30_14_0),
		.in_wire_1_1(vertical_tile_31_14_to_tile_30_14_1),
		.in_wire_1_2(vertical_tile_31_14_to_tile_30_14_2),
		.in_wire_1_3(vertical_tile_31_14_to_tile_30_14_3),
		.out_wire_2_0(horizontal_tile_30_14_to_tile_30_13_0),
		.out_wire_2_1(horizontal_tile_30_14_to_tile_30_13_1),
		.out_wire_2_2(horizontal_tile_30_14_to_tile_30_13_2),
		.out_wire_2_3(horizontal_tile_30_14_to_tile_30_13_3),
		.in_wire_2_0(horizontal_tile_30_13_to_tile_30_14_0),
		.in_wire_2_1(horizontal_tile_30_13_to_tile_30_14_1),
		.in_wire_2_2(horizontal_tile_30_13_to_tile_30_14_2),
		.in_wire_2_3(horizontal_tile_30_13_to_tile_30_14_3),
		.out_wire_0_0(horizontal_tile_30_14_to_tile_30_15_0),
		.out_wire_0_1(horizontal_tile_30_14_to_tile_30_15_1),
		.out_wire_0_2(horizontal_tile_30_14_to_tile_30_15_2),
		.out_wire_0_3(horizontal_tile_30_14_to_tile_30_15_3),
		.in_wire_0_0(horizontal_tile_30_15_to_tile_30_14_0),
		.in_wire_0_1(horizontal_tile_30_15_to_tile_30_14_1),
		.in_wire_0_2(horizontal_tile_30_15_to_tile_30_14_2),
		.in_wire_0_3(horizontal_tile_30_15_to_tile_30_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(975)
	);

	pe_tile pe_tile_30_15(
		.out_wire_3_0(vertical_tile_30_15_to_tile_29_15_0),
		.out_wire_3_1(vertical_tile_30_15_to_tile_29_15_1),
		.out_wire_3_2(vertical_tile_30_15_to_tile_29_15_2),
		.out_wire_3_3(vertical_tile_30_15_to_tile_29_15_3),
		.in_wire_3_0(vertical_tile_29_15_to_tile_30_15_0),
		.in_wire_3_1(vertical_tile_29_15_to_tile_30_15_1),
		.in_wire_3_2(vertical_tile_29_15_to_tile_30_15_2),
		.in_wire_3_3(vertical_tile_29_15_to_tile_30_15_3),
		.out_wire_1_0(vertical_tile_30_15_to_tile_31_15_0),
		.out_wire_1_1(vertical_tile_30_15_to_tile_31_15_1),
		.out_wire_1_2(vertical_tile_30_15_to_tile_31_15_2),
		.out_wire_1_3(vertical_tile_30_15_to_tile_31_15_3),
		.in_wire_1_0(vertical_tile_31_15_to_tile_30_15_0),
		.in_wire_1_1(vertical_tile_31_15_to_tile_30_15_1),
		.in_wire_1_2(vertical_tile_31_15_to_tile_30_15_2),
		.in_wire_1_3(vertical_tile_31_15_to_tile_30_15_3),
		.out_wire_2_0(horizontal_tile_30_15_to_tile_30_14_0),
		.out_wire_2_1(horizontal_tile_30_15_to_tile_30_14_1),
		.out_wire_2_2(horizontal_tile_30_15_to_tile_30_14_2),
		.out_wire_2_3(horizontal_tile_30_15_to_tile_30_14_3),
		.in_wire_2_0(horizontal_tile_30_14_to_tile_30_15_0),
		.in_wire_2_1(horizontal_tile_30_14_to_tile_30_15_1),
		.in_wire_2_2(horizontal_tile_30_14_to_tile_30_15_2),
		.in_wire_2_3(horizontal_tile_30_14_to_tile_30_15_3),
		.out_wire_0_0(horizontal_tile_30_15_to_tile_30_16_0),
		.out_wire_0_1(horizontal_tile_30_15_to_tile_30_16_1),
		.out_wire_0_2(horizontal_tile_30_15_to_tile_30_16_2),
		.out_wire_0_3(horizontal_tile_30_15_to_tile_30_16_3),
		.in_wire_0_0(horizontal_tile_30_16_to_tile_30_15_0),
		.in_wire_0_1(horizontal_tile_30_16_to_tile_30_15_1),
		.in_wire_0_2(horizontal_tile_30_16_to_tile_30_15_2),
		.in_wire_0_3(horizontal_tile_30_16_to_tile_30_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(976)
	);

	pe_tile pe_tile_30_16(
		.out_wire_3_0(vertical_tile_30_16_to_tile_29_16_0),
		.out_wire_3_1(vertical_tile_30_16_to_tile_29_16_1),
		.out_wire_3_2(vertical_tile_30_16_to_tile_29_16_2),
		.out_wire_3_3(vertical_tile_30_16_to_tile_29_16_3),
		.in_wire_3_0(vertical_tile_29_16_to_tile_30_16_0),
		.in_wire_3_1(vertical_tile_29_16_to_tile_30_16_1),
		.in_wire_3_2(vertical_tile_29_16_to_tile_30_16_2),
		.in_wire_3_3(vertical_tile_29_16_to_tile_30_16_3),
		.out_wire_1_0(vertical_tile_30_16_to_tile_31_16_0),
		.out_wire_1_1(vertical_tile_30_16_to_tile_31_16_1),
		.out_wire_1_2(vertical_tile_30_16_to_tile_31_16_2),
		.out_wire_1_3(vertical_tile_30_16_to_tile_31_16_3),
		.in_wire_1_0(vertical_tile_31_16_to_tile_30_16_0),
		.in_wire_1_1(vertical_tile_31_16_to_tile_30_16_1),
		.in_wire_1_2(vertical_tile_31_16_to_tile_30_16_2),
		.in_wire_1_3(vertical_tile_31_16_to_tile_30_16_3),
		.out_wire_2_0(horizontal_tile_30_16_to_tile_30_15_0),
		.out_wire_2_1(horizontal_tile_30_16_to_tile_30_15_1),
		.out_wire_2_2(horizontal_tile_30_16_to_tile_30_15_2),
		.out_wire_2_3(horizontal_tile_30_16_to_tile_30_15_3),
		.in_wire_2_0(horizontal_tile_30_15_to_tile_30_16_0),
		.in_wire_2_1(horizontal_tile_30_15_to_tile_30_16_1),
		.in_wire_2_2(horizontal_tile_30_15_to_tile_30_16_2),
		.in_wire_2_3(horizontal_tile_30_15_to_tile_30_16_3),
		.out_wire_0_0(horizontal_tile_30_16_to_tile_30_17_0),
		.out_wire_0_1(horizontal_tile_30_16_to_tile_30_17_1),
		.out_wire_0_2(horizontal_tile_30_16_to_tile_30_17_2),
		.out_wire_0_3(horizontal_tile_30_16_to_tile_30_17_3),
		.in_wire_0_0(horizontal_tile_30_17_to_tile_30_16_0),
		.in_wire_0_1(horizontal_tile_30_17_to_tile_30_16_1),
		.in_wire_0_2(horizontal_tile_30_17_to_tile_30_16_2),
		.in_wire_0_3(horizontal_tile_30_17_to_tile_30_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(977)
	);

	pe_tile pe_tile_30_17(
		.out_wire_3_0(vertical_tile_30_17_to_tile_29_17_0),
		.out_wire_3_1(vertical_tile_30_17_to_tile_29_17_1),
		.out_wire_3_2(vertical_tile_30_17_to_tile_29_17_2),
		.out_wire_3_3(vertical_tile_30_17_to_tile_29_17_3),
		.in_wire_3_0(vertical_tile_29_17_to_tile_30_17_0),
		.in_wire_3_1(vertical_tile_29_17_to_tile_30_17_1),
		.in_wire_3_2(vertical_tile_29_17_to_tile_30_17_2),
		.in_wire_3_3(vertical_tile_29_17_to_tile_30_17_3),
		.out_wire_1_0(vertical_tile_30_17_to_tile_31_17_0),
		.out_wire_1_1(vertical_tile_30_17_to_tile_31_17_1),
		.out_wire_1_2(vertical_tile_30_17_to_tile_31_17_2),
		.out_wire_1_3(vertical_tile_30_17_to_tile_31_17_3),
		.in_wire_1_0(vertical_tile_31_17_to_tile_30_17_0),
		.in_wire_1_1(vertical_tile_31_17_to_tile_30_17_1),
		.in_wire_1_2(vertical_tile_31_17_to_tile_30_17_2),
		.in_wire_1_3(vertical_tile_31_17_to_tile_30_17_3),
		.out_wire_2_0(horizontal_tile_30_17_to_tile_30_16_0),
		.out_wire_2_1(horizontal_tile_30_17_to_tile_30_16_1),
		.out_wire_2_2(horizontal_tile_30_17_to_tile_30_16_2),
		.out_wire_2_3(horizontal_tile_30_17_to_tile_30_16_3),
		.in_wire_2_0(horizontal_tile_30_16_to_tile_30_17_0),
		.in_wire_2_1(horizontal_tile_30_16_to_tile_30_17_1),
		.in_wire_2_2(horizontal_tile_30_16_to_tile_30_17_2),
		.in_wire_2_3(horizontal_tile_30_16_to_tile_30_17_3),
		.out_wire_0_0(horizontal_tile_30_17_to_tile_30_18_0),
		.out_wire_0_1(horizontal_tile_30_17_to_tile_30_18_1),
		.out_wire_0_2(horizontal_tile_30_17_to_tile_30_18_2),
		.out_wire_0_3(horizontal_tile_30_17_to_tile_30_18_3),
		.in_wire_0_0(horizontal_tile_30_18_to_tile_30_17_0),
		.in_wire_0_1(horizontal_tile_30_18_to_tile_30_17_1),
		.in_wire_0_2(horizontal_tile_30_18_to_tile_30_17_2),
		.in_wire_0_3(horizontal_tile_30_18_to_tile_30_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(978)
	);

	pe_tile pe_tile_30_18(
		.out_wire_3_0(vertical_tile_30_18_to_tile_29_18_0),
		.out_wire_3_1(vertical_tile_30_18_to_tile_29_18_1),
		.out_wire_3_2(vertical_tile_30_18_to_tile_29_18_2),
		.out_wire_3_3(vertical_tile_30_18_to_tile_29_18_3),
		.in_wire_3_0(vertical_tile_29_18_to_tile_30_18_0),
		.in_wire_3_1(vertical_tile_29_18_to_tile_30_18_1),
		.in_wire_3_2(vertical_tile_29_18_to_tile_30_18_2),
		.in_wire_3_3(vertical_tile_29_18_to_tile_30_18_3),
		.out_wire_1_0(vertical_tile_30_18_to_tile_31_18_0),
		.out_wire_1_1(vertical_tile_30_18_to_tile_31_18_1),
		.out_wire_1_2(vertical_tile_30_18_to_tile_31_18_2),
		.out_wire_1_3(vertical_tile_30_18_to_tile_31_18_3),
		.in_wire_1_0(vertical_tile_31_18_to_tile_30_18_0),
		.in_wire_1_1(vertical_tile_31_18_to_tile_30_18_1),
		.in_wire_1_2(vertical_tile_31_18_to_tile_30_18_2),
		.in_wire_1_3(vertical_tile_31_18_to_tile_30_18_3),
		.out_wire_2_0(horizontal_tile_30_18_to_tile_30_17_0),
		.out_wire_2_1(horizontal_tile_30_18_to_tile_30_17_1),
		.out_wire_2_2(horizontal_tile_30_18_to_tile_30_17_2),
		.out_wire_2_3(horizontal_tile_30_18_to_tile_30_17_3),
		.in_wire_2_0(horizontal_tile_30_17_to_tile_30_18_0),
		.in_wire_2_1(horizontal_tile_30_17_to_tile_30_18_1),
		.in_wire_2_2(horizontal_tile_30_17_to_tile_30_18_2),
		.in_wire_2_3(horizontal_tile_30_17_to_tile_30_18_3),
		.out_wire_0_0(horizontal_tile_30_18_to_tile_30_19_0),
		.out_wire_0_1(horizontal_tile_30_18_to_tile_30_19_1),
		.out_wire_0_2(horizontal_tile_30_18_to_tile_30_19_2),
		.out_wire_0_3(horizontal_tile_30_18_to_tile_30_19_3),
		.in_wire_0_0(horizontal_tile_30_19_to_tile_30_18_0),
		.in_wire_0_1(horizontal_tile_30_19_to_tile_30_18_1),
		.in_wire_0_2(horizontal_tile_30_19_to_tile_30_18_2),
		.in_wire_0_3(horizontal_tile_30_19_to_tile_30_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(979)
	);

	pe_tile pe_tile_30_19(
		.out_wire_3_0(vertical_tile_30_19_to_tile_29_19_0),
		.out_wire_3_1(vertical_tile_30_19_to_tile_29_19_1),
		.out_wire_3_2(vertical_tile_30_19_to_tile_29_19_2),
		.out_wire_3_3(vertical_tile_30_19_to_tile_29_19_3),
		.in_wire_3_0(vertical_tile_29_19_to_tile_30_19_0),
		.in_wire_3_1(vertical_tile_29_19_to_tile_30_19_1),
		.in_wire_3_2(vertical_tile_29_19_to_tile_30_19_2),
		.in_wire_3_3(vertical_tile_29_19_to_tile_30_19_3),
		.out_wire_1_0(vertical_tile_30_19_to_tile_31_19_0),
		.out_wire_1_1(vertical_tile_30_19_to_tile_31_19_1),
		.out_wire_1_2(vertical_tile_30_19_to_tile_31_19_2),
		.out_wire_1_3(vertical_tile_30_19_to_tile_31_19_3),
		.in_wire_1_0(vertical_tile_31_19_to_tile_30_19_0),
		.in_wire_1_1(vertical_tile_31_19_to_tile_30_19_1),
		.in_wire_1_2(vertical_tile_31_19_to_tile_30_19_2),
		.in_wire_1_3(vertical_tile_31_19_to_tile_30_19_3),
		.out_wire_2_0(horizontal_tile_30_19_to_tile_30_18_0),
		.out_wire_2_1(horizontal_tile_30_19_to_tile_30_18_1),
		.out_wire_2_2(horizontal_tile_30_19_to_tile_30_18_2),
		.out_wire_2_3(horizontal_tile_30_19_to_tile_30_18_3),
		.in_wire_2_0(horizontal_tile_30_18_to_tile_30_19_0),
		.in_wire_2_1(horizontal_tile_30_18_to_tile_30_19_1),
		.in_wire_2_2(horizontal_tile_30_18_to_tile_30_19_2),
		.in_wire_2_3(horizontal_tile_30_18_to_tile_30_19_3),
		.out_wire_0_0(horizontal_tile_30_19_to_tile_30_20_0),
		.out_wire_0_1(horizontal_tile_30_19_to_tile_30_20_1),
		.out_wire_0_2(horizontal_tile_30_19_to_tile_30_20_2),
		.out_wire_0_3(horizontal_tile_30_19_to_tile_30_20_3),
		.in_wire_0_0(horizontal_tile_30_20_to_tile_30_19_0),
		.in_wire_0_1(horizontal_tile_30_20_to_tile_30_19_1),
		.in_wire_0_2(horizontal_tile_30_20_to_tile_30_19_2),
		.in_wire_0_3(horizontal_tile_30_20_to_tile_30_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(980)
	);

	pe_tile pe_tile_30_20(
		.out_wire_3_0(vertical_tile_30_20_to_tile_29_20_0),
		.out_wire_3_1(vertical_tile_30_20_to_tile_29_20_1),
		.out_wire_3_2(vertical_tile_30_20_to_tile_29_20_2),
		.out_wire_3_3(vertical_tile_30_20_to_tile_29_20_3),
		.in_wire_3_0(vertical_tile_29_20_to_tile_30_20_0),
		.in_wire_3_1(vertical_tile_29_20_to_tile_30_20_1),
		.in_wire_3_2(vertical_tile_29_20_to_tile_30_20_2),
		.in_wire_3_3(vertical_tile_29_20_to_tile_30_20_3),
		.out_wire_1_0(vertical_tile_30_20_to_tile_31_20_0),
		.out_wire_1_1(vertical_tile_30_20_to_tile_31_20_1),
		.out_wire_1_2(vertical_tile_30_20_to_tile_31_20_2),
		.out_wire_1_3(vertical_tile_30_20_to_tile_31_20_3),
		.in_wire_1_0(vertical_tile_31_20_to_tile_30_20_0),
		.in_wire_1_1(vertical_tile_31_20_to_tile_30_20_1),
		.in_wire_1_2(vertical_tile_31_20_to_tile_30_20_2),
		.in_wire_1_3(vertical_tile_31_20_to_tile_30_20_3),
		.out_wire_2_0(horizontal_tile_30_20_to_tile_30_19_0),
		.out_wire_2_1(horizontal_tile_30_20_to_tile_30_19_1),
		.out_wire_2_2(horizontal_tile_30_20_to_tile_30_19_2),
		.out_wire_2_3(horizontal_tile_30_20_to_tile_30_19_3),
		.in_wire_2_0(horizontal_tile_30_19_to_tile_30_20_0),
		.in_wire_2_1(horizontal_tile_30_19_to_tile_30_20_1),
		.in_wire_2_2(horizontal_tile_30_19_to_tile_30_20_2),
		.in_wire_2_3(horizontal_tile_30_19_to_tile_30_20_3),
		.out_wire_0_0(horizontal_tile_30_20_to_tile_30_21_0),
		.out_wire_0_1(horizontal_tile_30_20_to_tile_30_21_1),
		.out_wire_0_2(horizontal_tile_30_20_to_tile_30_21_2),
		.out_wire_0_3(horizontal_tile_30_20_to_tile_30_21_3),
		.in_wire_0_0(horizontal_tile_30_21_to_tile_30_20_0),
		.in_wire_0_1(horizontal_tile_30_21_to_tile_30_20_1),
		.in_wire_0_2(horizontal_tile_30_21_to_tile_30_20_2),
		.in_wire_0_3(horizontal_tile_30_21_to_tile_30_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(981)
	);

	pe_tile pe_tile_30_21(
		.out_wire_3_0(vertical_tile_30_21_to_tile_29_21_0),
		.out_wire_3_1(vertical_tile_30_21_to_tile_29_21_1),
		.out_wire_3_2(vertical_tile_30_21_to_tile_29_21_2),
		.out_wire_3_3(vertical_tile_30_21_to_tile_29_21_3),
		.in_wire_3_0(vertical_tile_29_21_to_tile_30_21_0),
		.in_wire_3_1(vertical_tile_29_21_to_tile_30_21_1),
		.in_wire_3_2(vertical_tile_29_21_to_tile_30_21_2),
		.in_wire_3_3(vertical_tile_29_21_to_tile_30_21_3),
		.out_wire_1_0(vertical_tile_30_21_to_tile_31_21_0),
		.out_wire_1_1(vertical_tile_30_21_to_tile_31_21_1),
		.out_wire_1_2(vertical_tile_30_21_to_tile_31_21_2),
		.out_wire_1_3(vertical_tile_30_21_to_tile_31_21_3),
		.in_wire_1_0(vertical_tile_31_21_to_tile_30_21_0),
		.in_wire_1_1(vertical_tile_31_21_to_tile_30_21_1),
		.in_wire_1_2(vertical_tile_31_21_to_tile_30_21_2),
		.in_wire_1_3(vertical_tile_31_21_to_tile_30_21_3),
		.out_wire_2_0(horizontal_tile_30_21_to_tile_30_20_0),
		.out_wire_2_1(horizontal_tile_30_21_to_tile_30_20_1),
		.out_wire_2_2(horizontal_tile_30_21_to_tile_30_20_2),
		.out_wire_2_3(horizontal_tile_30_21_to_tile_30_20_3),
		.in_wire_2_0(horizontal_tile_30_20_to_tile_30_21_0),
		.in_wire_2_1(horizontal_tile_30_20_to_tile_30_21_1),
		.in_wire_2_2(horizontal_tile_30_20_to_tile_30_21_2),
		.in_wire_2_3(horizontal_tile_30_20_to_tile_30_21_3),
		.out_wire_0_0(horizontal_tile_30_21_to_tile_30_22_0),
		.out_wire_0_1(horizontal_tile_30_21_to_tile_30_22_1),
		.out_wire_0_2(horizontal_tile_30_21_to_tile_30_22_2),
		.out_wire_0_3(horizontal_tile_30_21_to_tile_30_22_3),
		.in_wire_0_0(horizontal_tile_30_22_to_tile_30_21_0),
		.in_wire_0_1(horizontal_tile_30_22_to_tile_30_21_1),
		.in_wire_0_2(horizontal_tile_30_22_to_tile_30_21_2),
		.in_wire_0_3(horizontal_tile_30_22_to_tile_30_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(982)
	);

	pe_tile pe_tile_30_22(
		.out_wire_3_0(vertical_tile_30_22_to_tile_29_22_0),
		.out_wire_3_1(vertical_tile_30_22_to_tile_29_22_1),
		.out_wire_3_2(vertical_tile_30_22_to_tile_29_22_2),
		.out_wire_3_3(vertical_tile_30_22_to_tile_29_22_3),
		.in_wire_3_0(vertical_tile_29_22_to_tile_30_22_0),
		.in_wire_3_1(vertical_tile_29_22_to_tile_30_22_1),
		.in_wire_3_2(vertical_tile_29_22_to_tile_30_22_2),
		.in_wire_3_3(vertical_tile_29_22_to_tile_30_22_3),
		.out_wire_1_0(vertical_tile_30_22_to_tile_31_22_0),
		.out_wire_1_1(vertical_tile_30_22_to_tile_31_22_1),
		.out_wire_1_2(vertical_tile_30_22_to_tile_31_22_2),
		.out_wire_1_3(vertical_tile_30_22_to_tile_31_22_3),
		.in_wire_1_0(vertical_tile_31_22_to_tile_30_22_0),
		.in_wire_1_1(vertical_tile_31_22_to_tile_30_22_1),
		.in_wire_1_2(vertical_tile_31_22_to_tile_30_22_2),
		.in_wire_1_3(vertical_tile_31_22_to_tile_30_22_3),
		.out_wire_2_0(horizontal_tile_30_22_to_tile_30_21_0),
		.out_wire_2_1(horizontal_tile_30_22_to_tile_30_21_1),
		.out_wire_2_2(horizontal_tile_30_22_to_tile_30_21_2),
		.out_wire_2_3(horizontal_tile_30_22_to_tile_30_21_3),
		.in_wire_2_0(horizontal_tile_30_21_to_tile_30_22_0),
		.in_wire_2_1(horizontal_tile_30_21_to_tile_30_22_1),
		.in_wire_2_2(horizontal_tile_30_21_to_tile_30_22_2),
		.in_wire_2_3(horizontal_tile_30_21_to_tile_30_22_3),
		.out_wire_0_0(horizontal_tile_30_22_to_tile_30_23_0),
		.out_wire_0_1(horizontal_tile_30_22_to_tile_30_23_1),
		.out_wire_0_2(horizontal_tile_30_22_to_tile_30_23_2),
		.out_wire_0_3(horizontal_tile_30_22_to_tile_30_23_3),
		.in_wire_0_0(horizontal_tile_30_23_to_tile_30_22_0),
		.in_wire_0_1(horizontal_tile_30_23_to_tile_30_22_1),
		.in_wire_0_2(horizontal_tile_30_23_to_tile_30_22_2),
		.in_wire_0_3(horizontal_tile_30_23_to_tile_30_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(983)
	);

	pe_tile pe_tile_30_23(
		.out_wire_3_0(vertical_tile_30_23_to_tile_29_23_0),
		.out_wire_3_1(vertical_tile_30_23_to_tile_29_23_1),
		.out_wire_3_2(vertical_tile_30_23_to_tile_29_23_2),
		.out_wire_3_3(vertical_tile_30_23_to_tile_29_23_3),
		.in_wire_3_0(vertical_tile_29_23_to_tile_30_23_0),
		.in_wire_3_1(vertical_tile_29_23_to_tile_30_23_1),
		.in_wire_3_2(vertical_tile_29_23_to_tile_30_23_2),
		.in_wire_3_3(vertical_tile_29_23_to_tile_30_23_3),
		.out_wire_1_0(vertical_tile_30_23_to_tile_31_23_0),
		.out_wire_1_1(vertical_tile_30_23_to_tile_31_23_1),
		.out_wire_1_2(vertical_tile_30_23_to_tile_31_23_2),
		.out_wire_1_3(vertical_tile_30_23_to_tile_31_23_3),
		.in_wire_1_0(vertical_tile_31_23_to_tile_30_23_0),
		.in_wire_1_1(vertical_tile_31_23_to_tile_30_23_1),
		.in_wire_1_2(vertical_tile_31_23_to_tile_30_23_2),
		.in_wire_1_3(vertical_tile_31_23_to_tile_30_23_3),
		.out_wire_2_0(horizontal_tile_30_23_to_tile_30_22_0),
		.out_wire_2_1(horizontal_tile_30_23_to_tile_30_22_1),
		.out_wire_2_2(horizontal_tile_30_23_to_tile_30_22_2),
		.out_wire_2_3(horizontal_tile_30_23_to_tile_30_22_3),
		.in_wire_2_0(horizontal_tile_30_22_to_tile_30_23_0),
		.in_wire_2_1(horizontal_tile_30_22_to_tile_30_23_1),
		.in_wire_2_2(horizontal_tile_30_22_to_tile_30_23_2),
		.in_wire_2_3(horizontal_tile_30_22_to_tile_30_23_3),
		.out_wire_0_0(horizontal_tile_30_23_to_tile_30_24_0),
		.out_wire_0_1(horizontal_tile_30_23_to_tile_30_24_1),
		.out_wire_0_2(horizontal_tile_30_23_to_tile_30_24_2),
		.out_wire_0_3(horizontal_tile_30_23_to_tile_30_24_3),
		.in_wire_0_0(horizontal_tile_30_24_to_tile_30_23_0),
		.in_wire_0_1(horizontal_tile_30_24_to_tile_30_23_1),
		.in_wire_0_2(horizontal_tile_30_24_to_tile_30_23_2),
		.in_wire_0_3(horizontal_tile_30_24_to_tile_30_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(984)
	);

	pe_tile pe_tile_30_24(
		.out_wire_3_0(vertical_tile_30_24_to_tile_29_24_0),
		.out_wire_3_1(vertical_tile_30_24_to_tile_29_24_1),
		.out_wire_3_2(vertical_tile_30_24_to_tile_29_24_2),
		.out_wire_3_3(vertical_tile_30_24_to_tile_29_24_3),
		.in_wire_3_0(vertical_tile_29_24_to_tile_30_24_0),
		.in_wire_3_1(vertical_tile_29_24_to_tile_30_24_1),
		.in_wire_3_2(vertical_tile_29_24_to_tile_30_24_2),
		.in_wire_3_3(vertical_tile_29_24_to_tile_30_24_3),
		.out_wire_1_0(vertical_tile_30_24_to_tile_31_24_0),
		.out_wire_1_1(vertical_tile_30_24_to_tile_31_24_1),
		.out_wire_1_2(vertical_tile_30_24_to_tile_31_24_2),
		.out_wire_1_3(vertical_tile_30_24_to_tile_31_24_3),
		.in_wire_1_0(vertical_tile_31_24_to_tile_30_24_0),
		.in_wire_1_1(vertical_tile_31_24_to_tile_30_24_1),
		.in_wire_1_2(vertical_tile_31_24_to_tile_30_24_2),
		.in_wire_1_3(vertical_tile_31_24_to_tile_30_24_3),
		.out_wire_2_0(horizontal_tile_30_24_to_tile_30_23_0),
		.out_wire_2_1(horizontal_tile_30_24_to_tile_30_23_1),
		.out_wire_2_2(horizontal_tile_30_24_to_tile_30_23_2),
		.out_wire_2_3(horizontal_tile_30_24_to_tile_30_23_3),
		.in_wire_2_0(horizontal_tile_30_23_to_tile_30_24_0),
		.in_wire_2_1(horizontal_tile_30_23_to_tile_30_24_1),
		.in_wire_2_2(horizontal_tile_30_23_to_tile_30_24_2),
		.in_wire_2_3(horizontal_tile_30_23_to_tile_30_24_3),
		.out_wire_0_0(horizontal_tile_30_24_to_tile_30_25_0),
		.out_wire_0_1(horizontal_tile_30_24_to_tile_30_25_1),
		.out_wire_0_2(horizontal_tile_30_24_to_tile_30_25_2),
		.out_wire_0_3(horizontal_tile_30_24_to_tile_30_25_3),
		.in_wire_0_0(horizontal_tile_30_25_to_tile_30_24_0),
		.in_wire_0_1(horizontal_tile_30_25_to_tile_30_24_1),
		.in_wire_0_2(horizontal_tile_30_25_to_tile_30_24_2),
		.in_wire_0_3(horizontal_tile_30_25_to_tile_30_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(985)
	);

	pe_tile pe_tile_30_25(
		.out_wire_3_0(vertical_tile_30_25_to_tile_29_25_0),
		.out_wire_3_1(vertical_tile_30_25_to_tile_29_25_1),
		.out_wire_3_2(vertical_tile_30_25_to_tile_29_25_2),
		.out_wire_3_3(vertical_tile_30_25_to_tile_29_25_3),
		.in_wire_3_0(vertical_tile_29_25_to_tile_30_25_0),
		.in_wire_3_1(vertical_tile_29_25_to_tile_30_25_1),
		.in_wire_3_2(vertical_tile_29_25_to_tile_30_25_2),
		.in_wire_3_3(vertical_tile_29_25_to_tile_30_25_3),
		.out_wire_1_0(vertical_tile_30_25_to_tile_31_25_0),
		.out_wire_1_1(vertical_tile_30_25_to_tile_31_25_1),
		.out_wire_1_2(vertical_tile_30_25_to_tile_31_25_2),
		.out_wire_1_3(vertical_tile_30_25_to_tile_31_25_3),
		.in_wire_1_0(vertical_tile_31_25_to_tile_30_25_0),
		.in_wire_1_1(vertical_tile_31_25_to_tile_30_25_1),
		.in_wire_1_2(vertical_tile_31_25_to_tile_30_25_2),
		.in_wire_1_3(vertical_tile_31_25_to_tile_30_25_3),
		.out_wire_2_0(horizontal_tile_30_25_to_tile_30_24_0),
		.out_wire_2_1(horizontal_tile_30_25_to_tile_30_24_1),
		.out_wire_2_2(horizontal_tile_30_25_to_tile_30_24_2),
		.out_wire_2_3(horizontal_tile_30_25_to_tile_30_24_3),
		.in_wire_2_0(horizontal_tile_30_24_to_tile_30_25_0),
		.in_wire_2_1(horizontal_tile_30_24_to_tile_30_25_1),
		.in_wire_2_2(horizontal_tile_30_24_to_tile_30_25_2),
		.in_wire_2_3(horizontal_tile_30_24_to_tile_30_25_3),
		.out_wire_0_0(horizontal_tile_30_25_to_tile_30_26_0),
		.out_wire_0_1(horizontal_tile_30_25_to_tile_30_26_1),
		.out_wire_0_2(horizontal_tile_30_25_to_tile_30_26_2),
		.out_wire_0_3(horizontal_tile_30_25_to_tile_30_26_3),
		.in_wire_0_0(horizontal_tile_30_26_to_tile_30_25_0),
		.in_wire_0_1(horizontal_tile_30_26_to_tile_30_25_1),
		.in_wire_0_2(horizontal_tile_30_26_to_tile_30_25_2),
		.in_wire_0_3(horizontal_tile_30_26_to_tile_30_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(986)
	);

	pe_tile pe_tile_30_26(
		.out_wire_3_0(vertical_tile_30_26_to_tile_29_26_0),
		.out_wire_3_1(vertical_tile_30_26_to_tile_29_26_1),
		.out_wire_3_2(vertical_tile_30_26_to_tile_29_26_2),
		.out_wire_3_3(vertical_tile_30_26_to_tile_29_26_3),
		.in_wire_3_0(vertical_tile_29_26_to_tile_30_26_0),
		.in_wire_3_1(vertical_tile_29_26_to_tile_30_26_1),
		.in_wire_3_2(vertical_tile_29_26_to_tile_30_26_2),
		.in_wire_3_3(vertical_tile_29_26_to_tile_30_26_3),
		.out_wire_1_0(vertical_tile_30_26_to_tile_31_26_0),
		.out_wire_1_1(vertical_tile_30_26_to_tile_31_26_1),
		.out_wire_1_2(vertical_tile_30_26_to_tile_31_26_2),
		.out_wire_1_3(vertical_tile_30_26_to_tile_31_26_3),
		.in_wire_1_0(vertical_tile_31_26_to_tile_30_26_0),
		.in_wire_1_1(vertical_tile_31_26_to_tile_30_26_1),
		.in_wire_1_2(vertical_tile_31_26_to_tile_30_26_2),
		.in_wire_1_3(vertical_tile_31_26_to_tile_30_26_3),
		.out_wire_2_0(horizontal_tile_30_26_to_tile_30_25_0),
		.out_wire_2_1(horizontal_tile_30_26_to_tile_30_25_1),
		.out_wire_2_2(horizontal_tile_30_26_to_tile_30_25_2),
		.out_wire_2_3(horizontal_tile_30_26_to_tile_30_25_3),
		.in_wire_2_0(horizontal_tile_30_25_to_tile_30_26_0),
		.in_wire_2_1(horizontal_tile_30_25_to_tile_30_26_1),
		.in_wire_2_2(horizontal_tile_30_25_to_tile_30_26_2),
		.in_wire_2_3(horizontal_tile_30_25_to_tile_30_26_3),
		.out_wire_0_0(horizontal_tile_30_26_to_tile_30_27_0),
		.out_wire_0_1(horizontal_tile_30_26_to_tile_30_27_1),
		.out_wire_0_2(horizontal_tile_30_26_to_tile_30_27_2),
		.out_wire_0_3(horizontal_tile_30_26_to_tile_30_27_3),
		.in_wire_0_0(horizontal_tile_30_27_to_tile_30_26_0),
		.in_wire_0_1(horizontal_tile_30_27_to_tile_30_26_1),
		.in_wire_0_2(horizontal_tile_30_27_to_tile_30_26_2),
		.in_wire_0_3(horizontal_tile_30_27_to_tile_30_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(987)
	);

	pe_tile pe_tile_30_27(
		.out_wire_3_0(vertical_tile_30_27_to_tile_29_27_0),
		.out_wire_3_1(vertical_tile_30_27_to_tile_29_27_1),
		.out_wire_3_2(vertical_tile_30_27_to_tile_29_27_2),
		.out_wire_3_3(vertical_tile_30_27_to_tile_29_27_3),
		.in_wire_3_0(vertical_tile_29_27_to_tile_30_27_0),
		.in_wire_3_1(vertical_tile_29_27_to_tile_30_27_1),
		.in_wire_3_2(vertical_tile_29_27_to_tile_30_27_2),
		.in_wire_3_3(vertical_tile_29_27_to_tile_30_27_3),
		.out_wire_1_0(vertical_tile_30_27_to_tile_31_27_0),
		.out_wire_1_1(vertical_tile_30_27_to_tile_31_27_1),
		.out_wire_1_2(vertical_tile_30_27_to_tile_31_27_2),
		.out_wire_1_3(vertical_tile_30_27_to_tile_31_27_3),
		.in_wire_1_0(vertical_tile_31_27_to_tile_30_27_0),
		.in_wire_1_1(vertical_tile_31_27_to_tile_30_27_1),
		.in_wire_1_2(vertical_tile_31_27_to_tile_30_27_2),
		.in_wire_1_3(vertical_tile_31_27_to_tile_30_27_3),
		.out_wire_2_0(horizontal_tile_30_27_to_tile_30_26_0),
		.out_wire_2_1(horizontal_tile_30_27_to_tile_30_26_1),
		.out_wire_2_2(horizontal_tile_30_27_to_tile_30_26_2),
		.out_wire_2_3(horizontal_tile_30_27_to_tile_30_26_3),
		.in_wire_2_0(horizontal_tile_30_26_to_tile_30_27_0),
		.in_wire_2_1(horizontal_tile_30_26_to_tile_30_27_1),
		.in_wire_2_2(horizontal_tile_30_26_to_tile_30_27_2),
		.in_wire_2_3(horizontal_tile_30_26_to_tile_30_27_3),
		.out_wire_0_0(horizontal_tile_30_27_to_tile_30_28_0),
		.out_wire_0_1(horizontal_tile_30_27_to_tile_30_28_1),
		.out_wire_0_2(horizontal_tile_30_27_to_tile_30_28_2),
		.out_wire_0_3(horizontal_tile_30_27_to_tile_30_28_3),
		.in_wire_0_0(horizontal_tile_30_28_to_tile_30_27_0),
		.in_wire_0_1(horizontal_tile_30_28_to_tile_30_27_1),
		.in_wire_0_2(horizontal_tile_30_28_to_tile_30_27_2),
		.in_wire_0_3(horizontal_tile_30_28_to_tile_30_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(988)
	);

	pe_tile pe_tile_30_28(
		.out_wire_3_0(vertical_tile_30_28_to_tile_29_28_0),
		.out_wire_3_1(vertical_tile_30_28_to_tile_29_28_1),
		.out_wire_3_2(vertical_tile_30_28_to_tile_29_28_2),
		.out_wire_3_3(vertical_tile_30_28_to_tile_29_28_3),
		.in_wire_3_0(vertical_tile_29_28_to_tile_30_28_0),
		.in_wire_3_1(vertical_tile_29_28_to_tile_30_28_1),
		.in_wire_3_2(vertical_tile_29_28_to_tile_30_28_2),
		.in_wire_3_3(vertical_tile_29_28_to_tile_30_28_3),
		.out_wire_1_0(vertical_tile_30_28_to_tile_31_28_0),
		.out_wire_1_1(vertical_tile_30_28_to_tile_31_28_1),
		.out_wire_1_2(vertical_tile_30_28_to_tile_31_28_2),
		.out_wire_1_3(vertical_tile_30_28_to_tile_31_28_3),
		.in_wire_1_0(vertical_tile_31_28_to_tile_30_28_0),
		.in_wire_1_1(vertical_tile_31_28_to_tile_30_28_1),
		.in_wire_1_2(vertical_tile_31_28_to_tile_30_28_2),
		.in_wire_1_3(vertical_tile_31_28_to_tile_30_28_3),
		.out_wire_2_0(horizontal_tile_30_28_to_tile_30_27_0),
		.out_wire_2_1(horizontal_tile_30_28_to_tile_30_27_1),
		.out_wire_2_2(horizontal_tile_30_28_to_tile_30_27_2),
		.out_wire_2_3(horizontal_tile_30_28_to_tile_30_27_3),
		.in_wire_2_0(horizontal_tile_30_27_to_tile_30_28_0),
		.in_wire_2_1(horizontal_tile_30_27_to_tile_30_28_1),
		.in_wire_2_2(horizontal_tile_30_27_to_tile_30_28_2),
		.in_wire_2_3(horizontal_tile_30_27_to_tile_30_28_3),
		.out_wire_0_0(horizontal_tile_30_28_to_tile_30_29_0),
		.out_wire_0_1(horizontal_tile_30_28_to_tile_30_29_1),
		.out_wire_0_2(horizontal_tile_30_28_to_tile_30_29_2),
		.out_wire_0_3(horizontal_tile_30_28_to_tile_30_29_3),
		.in_wire_0_0(horizontal_tile_30_29_to_tile_30_28_0),
		.in_wire_0_1(horizontal_tile_30_29_to_tile_30_28_1),
		.in_wire_0_2(horizontal_tile_30_29_to_tile_30_28_2),
		.in_wire_0_3(horizontal_tile_30_29_to_tile_30_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(989)
	);

	pe_tile pe_tile_30_29(
		.out_wire_3_0(vertical_tile_30_29_to_tile_29_29_0),
		.out_wire_3_1(vertical_tile_30_29_to_tile_29_29_1),
		.out_wire_3_2(vertical_tile_30_29_to_tile_29_29_2),
		.out_wire_3_3(vertical_tile_30_29_to_tile_29_29_3),
		.in_wire_3_0(vertical_tile_29_29_to_tile_30_29_0),
		.in_wire_3_1(vertical_tile_29_29_to_tile_30_29_1),
		.in_wire_3_2(vertical_tile_29_29_to_tile_30_29_2),
		.in_wire_3_3(vertical_tile_29_29_to_tile_30_29_3),
		.out_wire_1_0(vertical_tile_30_29_to_tile_31_29_0),
		.out_wire_1_1(vertical_tile_30_29_to_tile_31_29_1),
		.out_wire_1_2(vertical_tile_30_29_to_tile_31_29_2),
		.out_wire_1_3(vertical_tile_30_29_to_tile_31_29_3),
		.in_wire_1_0(vertical_tile_31_29_to_tile_30_29_0),
		.in_wire_1_1(vertical_tile_31_29_to_tile_30_29_1),
		.in_wire_1_2(vertical_tile_31_29_to_tile_30_29_2),
		.in_wire_1_3(vertical_tile_31_29_to_tile_30_29_3),
		.out_wire_2_0(horizontal_tile_30_29_to_tile_30_28_0),
		.out_wire_2_1(horizontal_tile_30_29_to_tile_30_28_1),
		.out_wire_2_2(horizontal_tile_30_29_to_tile_30_28_2),
		.out_wire_2_3(horizontal_tile_30_29_to_tile_30_28_3),
		.in_wire_2_0(horizontal_tile_30_28_to_tile_30_29_0),
		.in_wire_2_1(horizontal_tile_30_28_to_tile_30_29_1),
		.in_wire_2_2(horizontal_tile_30_28_to_tile_30_29_2),
		.in_wire_2_3(horizontal_tile_30_28_to_tile_30_29_3),
		.out_wire_0_0(horizontal_tile_30_29_to_tile_30_30_0),
		.out_wire_0_1(horizontal_tile_30_29_to_tile_30_30_1),
		.out_wire_0_2(horizontal_tile_30_29_to_tile_30_30_2),
		.out_wire_0_3(horizontal_tile_30_29_to_tile_30_30_3),
		.in_wire_0_0(horizontal_tile_30_30_to_tile_30_29_0),
		.in_wire_0_1(horizontal_tile_30_30_to_tile_30_29_1),
		.in_wire_0_2(horizontal_tile_30_30_to_tile_30_29_2),
		.in_wire_0_3(horizontal_tile_30_30_to_tile_30_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(990)
	);

	pe_tile pe_tile_30_30(
		.out_wire_3_0(vertical_tile_30_30_to_tile_29_30_0),
		.out_wire_3_1(vertical_tile_30_30_to_tile_29_30_1),
		.out_wire_3_2(vertical_tile_30_30_to_tile_29_30_2),
		.out_wire_3_3(vertical_tile_30_30_to_tile_29_30_3),
		.in_wire_3_0(vertical_tile_29_30_to_tile_30_30_0),
		.in_wire_3_1(vertical_tile_29_30_to_tile_30_30_1),
		.in_wire_3_2(vertical_tile_29_30_to_tile_30_30_2),
		.in_wire_3_3(vertical_tile_29_30_to_tile_30_30_3),
		.out_wire_1_0(vertical_tile_30_30_to_tile_31_30_0),
		.out_wire_1_1(vertical_tile_30_30_to_tile_31_30_1),
		.out_wire_1_2(vertical_tile_30_30_to_tile_31_30_2),
		.out_wire_1_3(vertical_tile_30_30_to_tile_31_30_3),
		.in_wire_1_0(vertical_tile_31_30_to_tile_30_30_0),
		.in_wire_1_1(vertical_tile_31_30_to_tile_30_30_1),
		.in_wire_1_2(vertical_tile_31_30_to_tile_30_30_2),
		.in_wire_1_3(vertical_tile_31_30_to_tile_30_30_3),
		.out_wire_2_0(horizontal_tile_30_30_to_tile_30_29_0),
		.out_wire_2_1(horizontal_tile_30_30_to_tile_30_29_1),
		.out_wire_2_2(horizontal_tile_30_30_to_tile_30_29_2),
		.out_wire_2_3(horizontal_tile_30_30_to_tile_30_29_3),
		.in_wire_2_0(horizontal_tile_30_29_to_tile_30_30_0),
		.in_wire_2_1(horizontal_tile_30_29_to_tile_30_30_1),
		.in_wire_2_2(horizontal_tile_30_29_to_tile_30_30_2),
		.in_wire_2_3(horizontal_tile_30_29_to_tile_30_30_3),
		.out_wire_0_0(horizontal_tile_30_30_to_tile_30_31_0),
		.out_wire_0_1(horizontal_tile_30_30_to_tile_30_31_1),
		.out_wire_0_2(horizontal_tile_30_30_to_tile_30_31_2),
		.out_wire_0_3(horizontal_tile_30_30_to_tile_30_31_3),
		.in_wire_0_0(horizontal_tile_30_31_to_tile_30_30_0),
		.in_wire_0_1(horizontal_tile_30_31_to_tile_30_30_1),
		.in_wire_0_2(horizontal_tile_30_31_to_tile_30_30_2),
		.in_wire_0_3(horizontal_tile_30_31_to_tile_30_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(991)
	);

	pe_tile_right pe_tile_30_31(
		.out_wire_3_0(vertical_tile_30_31_to_tile_29_31_0),
		.out_wire_3_1(vertical_tile_30_31_to_tile_29_31_1),
		.out_wire_3_2(vertical_tile_30_31_to_tile_29_31_2),
		.out_wire_3_3(vertical_tile_30_31_to_tile_29_31_3),
		.in_wire_3_0(vertical_tile_29_31_to_tile_30_31_0),
		.in_wire_3_1(vertical_tile_29_31_to_tile_30_31_1),
		.in_wire_3_2(vertical_tile_29_31_to_tile_30_31_2),
		.in_wire_3_3(vertical_tile_29_31_to_tile_30_31_3),
		.out_wire_1_0(vertical_tile_30_31_to_tile_31_31_0),
		.out_wire_1_1(vertical_tile_30_31_to_tile_31_31_1),
		.out_wire_1_2(vertical_tile_30_31_to_tile_31_31_2),
		.out_wire_1_3(vertical_tile_30_31_to_tile_31_31_3),
		.in_wire_1_0(vertical_tile_31_31_to_tile_30_31_0),
		.in_wire_1_1(vertical_tile_31_31_to_tile_30_31_1),
		.in_wire_1_2(vertical_tile_31_31_to_tile_30_31_2),
		.in_wire_1_3(vertical_tile_31_31_to_tile_30_31_3),
		.out_wire_2_0(horizontal_tile_30_31_to_tile_30_30_0),
		.out_wire_2_1(horizontal_tile_30_31_to_tile_30_30_1),
		.out_wire_2_2(horizontal_tile_30_31_to_tile_30_30_2),
		.out_wire_2_3(horizontal_tile_30_31_to_tile_30_30_3),
		.in_wire_2_0(horizontal_tile_30_30_to_tile_30_31_0),
		.in_wire_2_1(horizontal_tile_30_30_to_tile_30_31_1),
		.in_wire_2_2(horizontal_tile_30_30_to_tile_30_31_2),
		.in_wire_2_3(horizontal_tile_30_30_to_tile_30_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(992)
	);

	pe_tile_bottom_left pe_tile_31_0(
		.out_wire_3_0(vertical_tile_31_0_to_tile_30_0_0),
		.out_wire_3_1(vertical_tile_31_0_to_tile_30_0_1),
		.out_wire_3_2(vertical_tile_31_0_to_tile_30_0_2),
		.out_wire_3_3(vertical_tile_31_0_to_tile_30_0_3),
		.in_wire_3_0(vertical_tile_30_0_to_tile_31_0_0),
		.in_wire_3_1(vertical_tile_30_0_to_tile_31_0_1),
		.in_wire_3_2(vertical_tile_30_0_to_tile_31_0_2),
		.in_wire_3_3(vertical_tile_30_0_to_tile_31_0_3),
		.out_wire_1_0(grid_to_output_0),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.in_wire_2_0(1'b0),
		.in_wire_2_1(1'b0),
		.in_wire_2_2(1'b0),
		.in_wire_2_3(1'b0),
		.out_wire_0_0(horizontal_tile_31_0_to_tile_31_1_0),
		.out_wire_0_1(horizontal_tile_31_0_to_tile_31_1_1),
		.out_wire_0_2(horizontal_tile_31_0_to_tile_31_1_2),
		.out_wire_0_3(horizontal_tile_31_0_to_tile_31_1_3),
		.in_wire_0_0(horizontal_tile_31_1_to_tile_31_0_0),
		.in_wire_0_1(horizontal_tile_31_1_to_tile_31_0_1),
		.in_wire_0_2(horizontal_tile_31_1_to_tile_31_0_2),
		.in_wire_0_3(horizontal_tile_31_1_to_tile_31_0_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(993)
	);

	pe_tile_bottom pe_tile_31_1(
		.out_wire_3_0(vertical_tile_31_1_to_tile_30_1_0),
		.out_wire_3_1(vertical_tile_31_1_to_tile_30_1_1),
		.out_wire_3_2(vertical_tile_31_1_to_tile_30_1_2),
		.out_wire_3_3(vertical_tile_31_1_to_tile_30_1_3),
		.in_wire_3_0(vertical_tile_30_1_to_tile_31_1_0),
		.in_wire_3_1(vertical_tile_30_1_to_tile_31_1_1),
		.in_wire_3_2(vertical_tile_30_1_to_tile_31_1_2),
		.in_wire_3_3(vertical_tile_30_1_to_tile_31_1_3),
		.out_wire_1_0(grid_to_output_1),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_1_to_tile_31_0_0),
		.out_wire_2_1(horizontal_tile_31_1_to_tile_31_0_1),
		.out_wire_2_2(horizontal_tile_31_1_to_tile_31_0_2),
		.out_wire_2_3(horizontal_tile_31_1_to_tile_31_0_3),
		.in_wire_2_0(horizontal_tile_31_0_to_tile_31_1_0),
		.in_wire_2_1(horizontal_tile_31_0_to_tile_31_1_1),
		.in_wire_2_2(horizontal_tile_31_0_to_tile_31_1_2),
		.in_wire_2_3(horizontal_tile_31_0_to_tile_31_1_3),
		.out_wire_0_0(horizontal_tile_31_1_to_tile_31_2_0),
		.out_wire_0_1(horizontal_tile_31_1_to_tile_31_2_1),
		.out_wire_0_2(horizontal_tile_31_1_to_tile_31_2_2),
		.out_wire_0_3(horizontal_tile_31_1_to_tile_31_2_3),
		.in_wire_0_0(horizontal_tile_31_2_to_tile_31_1_0),
		.in_wire_0_1(horizontal_tile_31_2_to_tile_31_1_1),
		.in_wire_0_2(horizontal_tile_31_2_to_tile_31_1_2),
		.in_wire_0_3(horizontal_tile_31_2_to_tile_31_1_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(994)
	);

	pe_tile_bottom pe_tile_31_2(
		.out_wire_3_0(vertical_tile_31_2_to_tile_30_2_0),
		.out_wire_3_1(vertical_tile_31_2_to_tile_30_2_1),
		.out_wire_3_2(vertical_tile_31_2_to_tile_30_2_2),
		.out_wire_3_3(vertical_tile_31_2_to_tile_30_2_3),
		.in_wire_3_0(vertical_tile_30_2_to_tile_31_2_0),
		.in_wire_3_1(vertical_tile_30_2_to_tile_31_2_1),
		.in_wire_3_2(vertical_tile_30_2_to_tile_31_2_2),
		.in_wire_3_3(vertical_tile_30_2_to_tile_31_2_3),
		.out_wire_1_0(grid_to_output_2),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_2_to_tile_31_1_0),
		.out_wire_2_1(horizontal_tile_31_2_to_tile_31_1_1),
		.out_wire_2_2(horizontal_tile_31_2_to_tile_31_1_2),
		.out_wire_2_3(horizontal_tile_31_2_to_tile_31_1_3),
		.in_wire_2_0(horizontal_tile_31_1_to_tile_31_2_0),
		.in_wire_2_1(horizontal_tile_31_1_to_tile_31_2_1),
		.in_wire_2_2(horizontal_tile_31_1_to_tile_31_2_2),
		.in_wire_2_3(horizontal_tile_31_1_to_tile_31_2_3),
		.out_wire_0_0(horizontal_tile_31_2_to_tile_31_3_0),
		.out_wire_0_1(horizontal_tile_31_2_to_tile_31_3_1),
		.out_wire_0_2(horizontal_tile_31_2_to_tile_31_3_2),
		.out_wire_0_3(horizontal_tile_31_2_to_tile_31_3_3),
		.in_wire_0_0(horizontal_tile_31_3_to_tile_31_2_0),
		.in_wire_0_1(horizontal_tile_31_3_to_tile_31_2_1),
		.in_wire_0_2(horizontal_tile_31_3_to_tile_31_2_2),
		.in_wire_0_3(horizontal_tile_31_3_to_tile_31_2_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(995)
	);

	pe_tile_bottom pe_tile_31_3(
		.out_wire_3_0(vertical_tile_31_3_to_tile_30_3_0),
		.out_wire_3_1(vertical_tile_31_3_to_tile_30_3_1),
		.out_wire_3_2(vertical_tile_31_3_to_tile_30_3_2),
		.out_wire_3_3(vertical_tile_31_3_to_tile_30_3_3),
		.in_wire_3_0(vertical_tile_30_3_to_tile_31_3_0),
		.in_wire_3_1(vertical_tile_30_3_to_tile_31_3_1),
		.in_wire_3_2(vertical_tile_30_3_to_tile_31_3_2),
		.in_wire_3_3(vertical_tile_30_3_to_tile_31_3_3),
		.out_wire_1_0(grid_to_output_3),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_3_to_tile_31_2_0),
		.out_wire_2_1(horizontal_tile_31_3_to_tile_31_2_1),
		.out_wire_2_2(horizontal_tile_31_3_to_tile_31_2_2),
		.out_wire_2_3(horizontal_tile_31_3_to_tile_31_2_3),
		.in_wire_2_0(horizontal_tile_31_2_to_tile_31_3_0),
		.in_wire_2_1(horizontal_tile_31_2_to_tile_31_3_1),
		.in_wire_2_2(horizontal_tile_31_2_to_tile_31_3_2),
		.in_wire_2_3(horizontal_tile_31_2_to_tile_31_3_3),
		.out_wire_0_0(horizontal_tile_31_3_to_tile_31_4_0),
		.out_wire_0_1(horizontal_tile_31_3_to_tile_31_4_1),
		.out_wire_0_2(horizontal_tile_31_3_to_tile_31_4_2),
		.out_wire_0_3(horizontal_tile_31_3_to_tile_31_4_3),
		.in_wire_0_0(horizontal_tile_31_4_to_tile_31_3_0),
		.in_wire_0_1(horizontal_tile_31_4_to_tile_31_3_1),
		.in_wire_0_2(horizontal_tile_31_4_to_tile_31_3_2),
		.in_wire_0_3(horizontal_tile_31_4_to_tile_31_3_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(996)
	);

	pe_tile_bottom pe_tile_31_4(
		.out_wire_3_0(vertical_tile_31_4_to_tile_30_4_0),
		.out_wire_3_1(vertical_tile_31_4_to_tile_30_4_1),
		.out_wire_3_2(vertical_tile_31_4_to_tile_30_4_2),
		.out_wire_3_3(vertical_tile_31_4_to_tile_30_4_3),
		.in_wire_3_0(vertical_tile_30_4_to_tile_31_4_0),
		.in_wire_3_1(vertical_tile_30_4_to_tile_31_4_1),
		.in_wire_3_2(vertical_tile_30_4_to_tile_31_4_2),
		.in_wire_3_3(vertical_tile_30_4_to_tile_31_4_3),
		.out_wire_1_0(grid_to_output_4),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_4_to_tile_31_3_0),
		.out_wire_2_1(horizontal_tile_31_4_to_tile_31_3_1),
		.out_wire_2_2(horizontal_tile_31_4_to_tile_31_3_2),
		.out_wire_2_3(horizontal_tile_31_4_to_tile_31_3_3),
		.in_wire_2_0(horizontal_tile_31_3_to_tile_31_4_0),
		.in_wire_2_1(horizontal_tile_31_3_to_tile_31_4_1),
		.in_wire_2_2(horizontal_tile_31_3_to_tile_31_4_2),
		.in_wire_2_3(horizontal_tile_31_3_to_tile_31_4_3),
		.out_wire_0_0(horizontal_tile_31_4_to_tile_31_5_0),
		.out_wire_0_1(horizontal_tile_31_4_to_tile_31_5_1),
		.out_wire_0_2(horizontal_tile_31_4_to_tile_31_5_2),
		.out_wire_0_3(horizontal_tile_31_4_to_tile_31_5_3),
		.in_wire_0_0(horizontal_tile_31_5_to_tile_31_4_0),
		.in_wire_0_1(horizontal_tile_31_5_to_tile_31_4_1),
		.in_wire_0_2(horizontal_tile_31_5_to_tile_31_4_2),
		.in_wire_0_3(horizontal_tile_31_5_to_tile_31_4_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(997)
	);

	pe_tile_bottom pe_tile_31_5(
		.out_wire_3_0(vertical_tile_31_5_to_tile_30_5_0),
		.out_wire_3_1(vertical_tile_31_5_to_tile_30_5_1),
		.out_wire_3_2(vertical_tile_31_5_to_tile_30_5_2),
		.out_wire_3_3(vertical_tile_31_5_to_tile_30_5_3),
		.in_wire_3_0(vertical_tile_30_5_to_tile_31_5_0),
		.in_wire_3_1(vertical_tile_30_5_to_tile_31_5_1),
		.in_wire_3_2(vertical_tile_30_5_to_tile_31_5_2),
		.in_wire_3_3(vertical_tile_30_5_to_tile_31_5_3),
		.out_wire_1_0(grid_to_output_5),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_5_to_tile_31_4_0),
		.out_wire_2_1(horizontal_tile_31_5_to_tile_31_4_1),
		.out_wire_2_2(horizontal_tile_31_5_to_tile_31_4_2),
		.out_wire_2_3(horizontal_tile_31_5_to_tile_31_4_3),
		.in_wire_2_0(horizontal_tile_31_4_to_tile_31_5_0),
		.in_wire_2_1(horizontal_tile_31_4_to_tile_31_5_1),
		.in_wire_2_2(horizontal_tile_31_4_to_tile_31_5_2),
		.in_wire_2_3(horizontal_tile_31_4_to_tile_31_5_3),
		.out_wire_0_0(horizontal_tile_31_5_to_tile_31_6_0),
		.out_wire_0_1(horizontal_tile_31_5_to_tile_31_6_1),
		.out_wire_0_2(horizontal_tile_31_5_to_tile_31_6_2),
		.out_wire_0_3(horizontal_tile_31_5_to_tile_31_6_3),
		.in_wire_0_0(horizontal_tile_31_6_to_tile_31_5_0),
		.in_wire_0_1(horizontal_tile_31_6_to_tile_31_5_1),
		.in_wire_0_2(horizontal_tile_31_6_to_tile_31_5_2),
		.in_wire_0_3(horizontal_tile_31_6_to_tile_31_5_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(998)
	);

	pe_tile_bottom pe_tile_31_6(
		.out_wire_3_0(vertical_tile_31_6_to_tile_30_6_0),
		.out_wire_3_1(vertical_tile_31_6_to_tile_30_6_1),
		.out_wire_3_2(vertical_tile_31_6_to_tile_30_6_2),
		.out_wire_3_3(vertical_tile_31_6_to_tile_30_6_3),
		.in_wire_3_0(vertical_tile_30_6_to_tile_31_6_0),
		.in_wire_3_1(vertical_tile_30_6_to_tile_31_6_1),
		.in_wire_3_2(vertical_tile_30_6_to_tile_31_6_2),
		.in_wire_3_3(vertical_tile_30_6_to_tile_31_6_3),
		.out_wire_1_0(grid_to_output_6),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_6_to_tile_31_5_0),
		.out_wire_2_1(horizontal_tile_31_6_to_tile_31_5_1),
		.out_wire_2_2(horizontal_tile_31_6_to_tile_31_5_2),
		.out_wire_2_3(horizontal_tile_31_6_to_tile_31_5_3),
		.in_wire_2_0(horizontal_tile_31_5_to_tile_31_6_0),
		.in_wire_2_1(horizontal_tile_31_5_to_tile_31_6_1),
		.in_wire_2_2(horizontal_tile_31_5_to_tile_31_6_2),
		.in_wire_2_3(horizontal_tile_31_5_to_tile_31_6_3),
		.out_wire_0_0(horizontal_tile_31_6_to_tile_31_7_0),
		.out_wire_0_1(horizontal_tile_31_6_to_tile_31_7_1),
		.out_wire_0_2(horizontal_tile_31_6_to_tile_31_7_2),
		.out_wire_0_3(horizontal_tile_31_6_to_tile_31_7_3),
		.in_wire_0_0(horizontal_tile_31_7_to_tile_31_6_0),
		.in_wire_0_1(horizontal_tile_31_7_to_tile_31_6_1),
		.in_wire_0_2(horizontal_tile_31_7_to_tile_31_6_2),
		.in_wire_0_3(horizontal_tile_31_7_to_tile_31_6_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(999)
	);

	pe_tile_bottom pe_tile_31_7(
		.out_wire_3_0(vertical_tile_31_7_to_tile_30_7_0),
		.out_wire_3_1(vertical_tile_31_7_to_tile_30_7_1),
		.out_wire_3_2(vertical_tile_31_7_to_tile_30_7_2),
		.out_wire_3_3(vertical_tile_31_7_to_tile_30_7_3),
		.in_wire_3_0(vertical_tile_30_7_to_tile_31_7_0),
		.in_wire_3_1(vertical_tile_30_7_to_tile_31_7_1),
		.in_wire_3_2(vertical_tile_30_7_to_tile_31_7_2),
		.in_wire_3_3(vertical_tile_30_7_to_tile_31_7_3),
		.out_wire_1_0(grid_to_output_7),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_7_to_tile_31_6_0),
		.out_wire_2_1(horizontal_tile_31_7_to_tile_31_6_1),
		.out_wire_2_2(horizontal_tile_31_7_to_tile_31_6_2),
		.out_wire_2_3(horizontal_tile_31_7_to_tile_31_6_3),
		.in_wire_2_0(horizontal_tile_31_6_to_tile_31_7_0),
		.in_wire_2_1(horizontal_tile_31_6_to_tile_31_7_1),
		.in_wire_2_2(horizontal_tile_31_6_to_tile_31_7_2),
		.in_wire_2_3(horizontal_tile_31_6_to_tile_31_7_3),
		.out_wire_0_0(horizontal_tile_31_7_to_tile_31_8_0),
		.out_wire_0_1(horizontal_tile_31_7_to_tile_31_8_1),
		.out_wire_0_2(horizontal_tile_31_7_to_tile_31_8_2),
		.out_wire_0_3(horizontal_tile_31_7_to_tile_31_8_3),
		.in_wire_0_0(horizontal_tile_31_8_to_tile_31_7_0),
		.in_wire_0_1(horizontal_tile_31_8_to_tile_31_7_1),
		.in_wire_0_2(horizontal_tile_31_8_to_tile_31_7_2),
		.in_wire_0_3(horizontal_tile_31_8_to_tile_31_7_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1000)
	);

	pe_tile_bottom pe_tile_31_8(
		.out_wire_3_0(vertical_tile_31_8_to_tile_30_8_0),
		.out_wire_3_1(vertical_tile_31_8_to_tile_30_8_1),
		.out_wire_3_2(vertical_tile_31_8_to_tile_30_8_2),
		.out_wire_3_3(vertical_tile_31_8_to_tile_30_8_3),
		.in_wire_3_0(vertical_tile_30_8_to_tile_31_8_0),
		.in_wire_3_1(vertical_tile_30_8_to_tile_31_8_1),
		.in_wire_3_2(vertical_tile_30_8_to_tile_31_8_2),
		.in_wire_3_3(vertical_tile_30_8_to_tile_31_8_3),
		.out_wire_1_0(grid_to_output_8),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_8_to_tile_31_7_0),
		.out_wire_2_1(horizontal_tile_31_8_to_tile_31_7_1),
		.out_wire_2_2(horizontal_tile_31_8_to_tile_31_7_2),
		.out_wire_2_3(horizontal_tile_31_8_to_tile_31_7_3),
		.in_wire_2_0(horizontal_tile_31_7_to_tile_31_8_0),
		.in_wire_2_1(horizontal_tile_31_7_to_tile_31_8_1),
		.in_wire_2_2(horizontal_tile_31_7_to_tile_31_8_2),
		.in_wire_2_3(horizontal_tile_31_7_to_tile_31_8_3),
		.out_wire_0_0(horizontal_tile_31_8_to_tile_31_9_0),
		.out_wire_0_1(horizontal_tile_31_8_to_tile_31_9_1),
		.out_wire_0_2(horizontal_tile_31_8_to_tile_31_9_2),
		.out_wire_0_3(horizontal_tile_31_8_to_tile_31_9_3),
		.in_wire_0_0(horizontal_tile_31_9_to_tile_31_8_0),
		.in_wire_0_1(horizontal_tile_31_9_to_tile_31_8_1),
		.in_wire_0_2(horizontal_tile_31_9_to_tile_31_8_2),
		.in_wire_0_3(horizontal_tile_31_9_to_tile_31_8_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1001)
	);

	pe_tile_bottom pe_tile_31_9(
		.out_wire_3_0(vertical_tile_31_9_to_tile_30_9_0),
		.out_wire_3_1(vertical_tile_31_9_to_tile_30_9_1),
		.out_wire_3_2(vertical_tile_31_9_to_tile_30_9_2),
		.out_wire_3_3(vertical_tile_31_9_to_tile_30_9_3),
		.in_wire_3_0(vertical_tile_30_9_to_tile_31_9_0),
		.in_wire_3_1(vertical_tile_30_9_to_tile_31_9_1),
		.in_wire_3_2(vertical_tile_30_9_to_tile_31_9_2),
		.in_wire_3_3(vertical_tile_30_9_to_tile_31_9_3),
		.out_wire_1_0(grid_to_output_9),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_9_to_tile_31_8_0),
		.out_wire_2_1(horizontal_tile_31_9_to_tile_31_8_1),
		.out_wire_2_2(horizontal_tile_31_9_to_tile_31_8_2),
		.out_wire_2_3(horizontal_tile_31_9_to_tile_31_8_3),
		.in_wire_2_0(horizontal_tile_31_8_to_tile_31_9_0),
		.in_wire_2_1(horizontal_tile_31_8_to_tile_31_9_1),
		.in_wire_2_2(horizontal_tile_31_8_to_tile_31_9_2),
		.in_wire_2_3(horizontal_tile_31_8_to_tile_31_9_3),
		.out_wire_0_0(horizontal_tile_31_9_to_tile_31_10_0),
		.out_wire_0_1(horizontal_tile_31_9_to_tile_31_10_1),
		.out_wire_0_2(horizontal_tile_31_9_to_tile_31_10_2),
		.out_wire_0_3(horizontal_tile_31_9_to_tile_31_10_3),
		.in_wire_0_0(horizontal_tile_31_10_to_tile_31_9_0),
		.in_wire_0_1(horizontal_tile_31_10_to_tile_31_9_1),
		.in_wire_0_2(horizontal_tile_31_10_to_tile_31_9_2),
		.in_wire_0_3(horizontal_tile_31_10_to_tile_31_9_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1002)
	);

	pe_tile_bottom pe_tile_31_10(
		.out_wire_3_0(vertical_tile_31_10_to_tile_30_10_0),
		.out_wire_3_1(vertical_tile_31_10_to_tile_30_10_1),
		.out_wire_3_2(vertical_tile_31_10_to_tile_30_10_2),
		.out_wire_3_3(vertical_tile_31_10_to_tile_30_10_3),
		.in_wire_3_0(vertical_tile_30_10_to_tile_31_10_0),
		.in_wire_3_1(vertical_tile_30_10_to_tile_31_10_1),
		.in_wire_3_2(vertical_tile_30_10_to_tile_31_10_2),
		.in_wire_3_3(vertical_tile_30_10_to_tile_31_10_3),
		.out_wire_1_0(grid_to_output_10),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_10_to_tile_31_9_0),
		.out_wire_2_1(horizontal_tile_31_10_to_tile_31_9_1),
		.out_wire_2_2(horizontal_tile_31_10_to_tile_31_9_2),
		.out_wire_2_3(horizontal_tile_31_10_to_tile_31_9_3),
		.in_wire_2_0(horizontal_tile_31_9_to_tile_31_10_0),
		.in_wire_2_1(horizontal_tile_31_9_to_tile_31_10_1),
		.in_wire_2_2(horizontal_tile_31_9_to_tile_31_10_2),
		.in_wire_2_3(horizontal_tile_31_9_to_tile_31_10_3),
		.out_wire_0_0(horizontal_tile_31_10_to_tile_31_11_0),
		.out_wire_0_1(horizontal_tile_31_10_to_tile_31_11_1),
		.out_wire_0_2(horizontal_tile_31_10_to_tile_31_11_2),
		.out_wire_0_3(horizontal_tile_31_10_to_tile_31_11_3),
		.in_wire_0_0(horizontal_tile_31_11_to_tile_31_10_0),
		.in_wire_0_1(horizontal_tile_31_11_to_tile_31_10_1),
		.in_wire_0_2(horizontal_tile_31_11_to_tile_31_10_2),
		.in_wire_0_3(horizontal_tile_31_11_to_tile_31_10_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1003)
	);

	pe_tile_bottom pe_tile_31_11(
		.out_wire_3_0(vertical_tile_31_11_to_tile_30_11_0),
		.out_wire_3_1(vertical_tile_31_11_to_tile_30_11_1),
		.out_wire_3_2(vertical_tile_31_11_to_tile_30_11_2),
		.out_wire_3_3(vertical_tile_31_11_to_tile_30_11_3),
		.in_wire_3_0(vertical_tile_30_11_to_tile_31_11_0),
		.in_wire_3_1(vertical_tile_30_11_to_tile_31_11_1),
		.in_wire_3_2(vertical_tile_30_11_to_tile_31_11_2),
		.in_wire_3_3(vertical_tile_30_11_to_tile_31_11_3),
		.out_wire_1_0(grid_to_output_11),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_11_to_tile_31_10_0),
		.out_wire_2_1(horizontal_tile_31_11_to_tile_31_10_1),
		.out_wire_2_2(horizontal_tile_31_11_to_tile_31_10_2),
		.out_wire_2_3(horizontal_tile_31_11_to_tile_31_10_3),
		.in_wire_2_0(horizontal_tile_31_10_to_tile_31_11_0),
		.in_wire_2_1(horizontal_tile_31_10_to_tile_31_11_1),
		.in_wire_2_2(horizontal_tile_31_10_to_tile_31_11_2),
		.in_wire_2_3(horizontal_tile_31_10_to_tile_31_11_3),
		.out_wire_0_0(horizontal_tile_31_11_to_tile_31_12_0),
		.out_wire_0_1(horizontal_tile_31_11_to_tile_31_12_1),
		.out_wire_0_2(horizontal_tile_31_11_to_tile_31_12_2),
		.out_wire_0_3(horizontal_tile_31_11_to_tile_31_12_3),
		.in_wire_0_0(horizontal_tile_31_12_to_tile_31_11_0),
		.in_wire_0_1(horizontal_tile_31_12_to_tile_31_11_1),
		.in_wire_0_2(horizontal_tile_31_12_to_tile_31_11_2),
		.in_wire_0_3(horizontal_tile_31_12_to_tile_31_11_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1004)
	);

	pe_tile_bottom pe_tile_31_12(
		.out_wire_3_0(vertical_tile_31_12_to_tile_30_12_0),
		.out_wire_3_1(vertical_tile_31_12_to_tile_30_12_1),
		.out_wire_3_2(vertical_tile_31_12_to_tile_30_12_2),
		.out_wire_3_3(vertical_tile_31_12_to_tile_30_12_3),
		.in_wire_3_0(vertical_tile_30_12_to_tile_31_12_0),
		.in_wire_3_1(vertical_tile_30_12_to_tile_31_12_1),
		.in_wire_3_2(vertical_tile_30_12_to_tile_31_12_2),
		.in_wire_3_3(vertical_tile_30_12_to_tile_31_12_3),
		.out_wire_1_0(grid_to_output_12),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_12_to_tile_31_11_0),
		.out_wire_2_1(horizontal_tile_31_12_to_tile_31_11_1),
		.out_wire_2_2(horizontal_tile_31_12_to_tile_31_11_2),
		.out_wire_2_3(horizontal_tile_31_12_to_tile_31_11_3),
		.in_wire_2_0(horizontal_tile_31_11_to_tile_31_12_0),
		.in_wire_2_1(horizontal_tile_31_11_to_tile_31_12_1),
		.in_wire_2_2(horizontal_tile_31_11_to_tile_31_12_2),
		.in_wire_2_3(horizontal_tile_31_11_to_tile_31_12_3),
		.out_wire_0_0(horizontal_tile_31_12_to_tile_31_13_0),
		.out_wire_0_1(horizontal_tile_31_12_to_tile_31_13_1),
		.out_wire_0_2(horizontal_tile_31_12_to_tile_31_13_2),
		.out_wire_0_3(horizontal_tile_31_12_to_tile_31_13_3),
		.in_wire_0_0(horizontal_tile_31_13_to_tile_31_12_0),
		.in_wire_0_1(horizontal_tile_31_13_to_tile_31_12_1),
		.in_wire_0_2(horizontal_tile_31_13_to_tile_31_12_2),
		.in_wire_0_3(horizontal_tile_31_13_to_tile_31_12_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1005)
	);

	pe_tile_bottom pe_tile_31_13(
		.out_wire_3_0(vertical_tile_31_13_to_tile_30_13_0),
		.out_wire_3_1(vertical_tile_31_13_to_tile_30_13_1),
		.out_wire_3_2(vertical_tile_31_13_to_tile_30_13_2),
		.out_wire_3_3(vertical_tile_31_13_to_tile_30_13_3),
		.in_wire_3_0(vertical_tile_30_13_to_tile_31_13_0),
		.in_wire_3_1(vertical_tile_30_13_to_tile_31_13_1),
		.in_wire_3_2(vertical_tile_30_13_to_tile_31_13_2),
		.in_wire_3_3(vertical_tile_30_13_to_tile_31_13_3),
		.out_wire_1_0(grid_to_output_13),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_13_to_tile_31_12_0),
		.out_wire_2_1(horizontal_tile_31_13_to_tile_31_12_1),
		.out_wire_2_2(horizontal_tile_31_13_to_tile_31_12_2),
		.out_wire_2_3(horizontal_tile_31_13_to_tile_31_12_3),
		.in_wire_2_0(horizontal_tile_31_12_to_tile_31_13_0),
		.in_wire_2_1(horizontal_tile_31_12_to_tile_31_13_1),
		.in_wire_2_2(horizontal_tile_31_12_to_tile_31_13_2),
		.in_wire_2_3(horizontal_tile_31_12_to_tile_31_13_3),
		.out_wire_0_0(horizontal_tile_31_13_to_tile_31_14_0),
		.out_wire_0_1(horizontal_tile_31_13_to_tile_31_14_1),
		.out_wire_0_2(horizontal_tile_31_13_to_tile_31_14_2),
		.out_wire_0_3(horizontal_tile_31_13_to_tile_31_14_3),
		.in_wire_0_0(horizontal_tile_31_14_to_tile_31_13_0),
		.in_wire_0_1(horizontal_tile_31_14_to_tile_31_13_1),
		.in_wire_0_2(horizontal_tile_31_14_to_tile_31_13_2),
		.in_wire_0_3(horizontal_tile_31_14_to_tile_31_13_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1006)
	);

	pe_tile_bottom pe_tile_31_14(
		.out_wire_3_0(vertical_tile_31_14_to_tile_30_14_0),
		.out_wire_3_1(vertical_tile_31_14_to_tile_30_14_1),
		.out_wire_3_2(vertical_tile_31_14_to_tile_30_14_2),
		.out_wire_3_3(vertical_tile_31_14_to_tile_30_14_3),
		.in_wire_3_0(vertical_tile_30_14_to_tile_31_14_0),
		.in_wire_3_1(vertical_tile_30_14_to_tile_31_14_1),
		.in_wire_3_2(vertical_tile_30_14_to_tile_31_14_2),
		.in_wire_3_3(vertical_tile_30_14_to_tile_31_14_3),
		.out_wire_1_0(grid_to_output_14),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_14_to_tile_31_13_0),
		.out_wire_2_1(horizontal_tile_31_14_to_tile_31_13_1),
		.out_wire_2_2(horizontal_tile_31_14_to_tile_31_13_2),
		.out_wire_2_3(horizontal_tile_31_14_to_tile_31_13_3),
		.in_wire_2_0(horizontal_tile_31_13_to_tile_31_14_0),
		.in_wire_2_1(horizontal_tile_31_13_to_tile_31_14_1),
		.in_wire_2_2(horizontal_tile_31_13_to_tile_31_14_2),
		.in_wire_2_3(horizontal_tile_31_13_to_tile_31_14_3),
		.out_wire_0_0(horizontal_tile_31_14_to_tile_31_15_0),
		.out_wire_0_1(horizontal_tile_31_14_to_tile_31_15_1),
		.out_wire_0_2(horizontal_tile_31_14_to_tile_31_15_2),
		.out_wire_0_3(horizontal_tile_31_14_to_tile_31_15_3),
		.in_wire_0_0(horizontal_tile_31_15_to_tile_31_14_0),
		.in_wire_0_1(horizontal_tile_31_15_to_tile_31_14_1),
		.in_wire_0_2(horizontal_tile_31_15_to_tile_31_14_2),
		.in_wire_0_3(horizontal_tile_31_15_to_tile_31_14_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1007)
	);

	pe_tile_bottom pe_tile_31_15(
		.out_wire_3_0(vertical_tile_31_15_to_tile_30_15_0),
		.out_wire_3_1(vertical_tile_31_15_to_tile_30_15_1),
		.out_wire_3_2(vertical_tile_31_15_to_tile_30_15_2),
		.out_wire_3_3(vertical_tile_31_15_to_tile_30_15_3),
		.in_wire_3_0(vertical_tile_30_15_to_tile_31_15_0),
		.in_wire_3_1(vertical_tile_30_15_to_tile_31_15_1),
		.in_wire_3_2(vertical_tile_30_15_to_tile_31_15_2),
		.in_wire_3_3(vertical_tile_30_15_to_tile_31_15_3),
		.out_wire_1_0(grid_to_output_15),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_15_to_tile_31_14_0),
		.out_wire_2_1(horizontal_tile_31_15_to_tile_31_14_1),
		.out_wire_2_2(horizontal_tile_31_15_to_tile_31_14_2),
		.out_wire_2_3(horizontal_tile_31_15_to_tile_31_14_3),
		.in_wire_2_0(horizontal_tile_31_14_to_tile_31_15_0),
		.in_wire_2_1(horizontal_tile_31_14_to_tile_31_15_1),
		.in_wire_2_2(horizontal_tile_31_14_to_tile_31_15_2),
		.in_wire_2_3(horizontal_tile_31_14_to_tile_31_15_3),
		.out_wire_0_0(horizontal_tile_31_15_to_tile_31_16_0),
		.out_wire_0_1(horizontal_tile_31_15_to_tile_31_16_1),
		.out_wire_0_2(horizontal_tile_31_15_to_tile_31_16_2),
		.out_wire_0_3(horizontal_tile_31_15_to_tile_31_16_3),
		.in_wire_0_0(horizontal_tile_31_16_to_tile_31_15_0),
		.in_wire_0_1(horizontal_tile_31_16_to_tile_31_15_1),
		.in_wire_0_2(horizontal_tile_31_16_to_tile_31_15_2),
		.in_wire_0_3(horizontal_tile_31_16_to_tile_31_15_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1008)
	);

	pe_tile_bottom pe_tile_31_16(
		.out_wire_3_0(vertical_tile_31_16_to_tile_30_16_0),
		.out_wire_3_1(vertical_tile_31_16_to_tile_30_16_1),
		.out_wire_3_2(vertical_tile_31_16_to_tile_30_16_2),
		.out_wire_3_3(vertical_tile_31_16_to_tile_30_16_3),
		.in_wire_3_0(vertical_tile_30_16_to_tile_31_16_0),
		.in_wire_3_1(vertical_tile_30_16_to_tile_31_16_1),
		.in_wire_3_2(vertical_tile_30_16_to_tile_31_16_2),
		.in_wire_3_3(vertical_tile_30_16_to_tile_31_16_3),
		.out_wire_1_0(grid_to_output_16),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_16_to_tile_31_15_0),
		.out_wire_2_1(horizontal_tile_31_16_to_tile_31_15_1),
		.out_wire_2_2(horizontal_tile_31_16_to_tile_31_15_2),
		.out_wire_2_3(horizontal_tile_31_16_to_tile_31_15_3),
		.in_wire_2_0(horizontal_tile_31_15_to_tile_31_16_0),
		.in_wire_2_1(horizontal_tile_31_15_to_tile_31_16_1),
		.in_wire_2_2(horizontal_tile_31_15_to_tile_31_16_2),
		.in_wire_2_3(horizontal_tile_31_15_to_tile_31_16_3),
		.out_wire_0_0(horizontal_tile_31_16_to_tile_31_17_0),
		.out_wire_0_1(horizontal_tile_31_16_to_tile_31_17_1),
		.out_wire_0_2(horizontal_tile_31_16_to_tile_31_17_2),
		.out_wire_0_3(horizontal_tile_31_16_to_tile_31_17_3),
		.in_wire_0_0(horizontal_tile_31_17_to_tile_31_16_0),
		.in_wire_0_1(horizontal_tile_31_17_to_tile_31_16_1),
		.in_wire_0_2(horizontal_tile_31_17_to_tile_31_16_2),
		.in_wire_0_3(horizontal_tile_31_17_to_tile_31_16_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1009)
	);

	pe_tile_bottom pe_tile_31_17(
		.out_wire_3_0(vertical_tile_31_17_to_tile_30_17_0),
		.out_wire_3_1(vertical_tile_31_17_to_tile_30_17_1),
		.out_wire_3_2(vertical_tile_31_17_to_tile_30_17_2),
		.out_wire_3_3(vertical_tile_31_17_to_tile_30_17_3),
		.in_wire_3_0(vertical_tile_30_17_to_tile_31_17_0),
		.in_wire_3_1(vertical_tile_30_17_to_tile_31_17_1),
		.in_wire_3_2(vertical_tile_30_17_to_tile_31_17_2),
		.in_wire_3_3(vertical_tile_30_17_to_tile_31_17_3),
		.out_wire_1_0(grid_to_output_17),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_17_to_tile_31_16_0),
		.out_wire_2_1(horizontal_tile_31_17_to_tile_31_16_1),
		.out_wire_2_2(horizontal_tile_31_17_to_tile_31_16_2),
		.out_wire_2_3(horizontal_tile_31_17_to_tile_31_16_3),
		.in_wire_2_0(horizontal_tile_31_16_to_tile_31_17_0),
		.in_wire_2_1(horizontal_tile_31_16_to_tile_31_17_1),
		.in_wire_2_2(horizontal_tile_31_16_to_tile_31_17_2),
		.in_wire_2_3(horizontal_tile_31_16_to_tile_31_17_3),
		.out_wire_0_0(horizontal_tile_31_17_to_tile_31_18_0),
		.out_wire_0_1(horizontal_tile_31_17_to_tile_31_18_1),
		.out_wire_0_2(horizontal_tile_31_17_to_tile_31_18_2),
		.out_wire_0_3(horizontal_tile_31_17_to_tile_31_18_3),
		.in_wire_0_0(horizontal_tile_31_18_to_tile_31_17_0),
		.in_wire_0_1(horizontal_tile_31_18_to_tile_31_17_1),
		.in_wire_0_2(horizontal_tile_31_18_to_tile_31_17_2),
		.in_wire_0_3(horizontal_tile_31_18_to_tile_31_17_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1010)
	);

	pe_tile_bottom pe_tile_31_18(
		.out_wire_3_0(vertical_tile_31_18_to_tile_30_18_0),
		.out_wire_3_1(vertical_tile_31_18_to_tile_30_18_1),
		.out_wire_3_2(vertical_tile_31_18_to_tile_30_18_2),
		.out_wire_3_3(vertical_tile_31_18_to_tile_30_18_3),
		.in_wire_3_0(vertical_tile_30_18_to_tile_31_18_0),
		.in_wire_3_1(vertical_tile_30_18_to_tile_31_18_1),
		.in_wire_3_2(vertical_tile_30_18_to_tile_31_18_2),
		.in_wire_3_3(vertical_tile_30_18_to_tile_31_18_3),
		.out_wire_1_0(grid_to_output_18),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_18_to_tile_31_17_0),
		.out_wire_2_1(horizontal_tile_31_18_to_tile_31_17_1),
		.out_wire_2_2(horizontal_tile_31_18_to_tile_31_17_2),
		.out_wire_2_3(horizontal_tile_31_18_to_tile_31_17_3),
		.in_wire_2_0(horizontal_tile_31_17_to_tile_31_18_0),
		.in_wire_2_1(horizontal_tile_31_17_to_tile_31_18_1),
		.in_wire_2_2(horizontal_tile_31_17_to_tile_31_18_2),
		.in_wire_2_3(horizontal_tile_31_17_to_tile_31_18_3),
		.out_wire_0_0(horizontal_tile_31_18_to_tile_31_19_0),
		.out_wire_0_1(horizontal_tile_31_18_to_tile_31_19_1),
		.out_wire_0_2(horizontal_tile_31_18_to_tile_31_19_2),
		.out_wire_0_3(horizontal_tile_31_18_to_tile_31_19_3),
		.in_wire_0_0(horizontal_tile_31_19_to_tile_31_18_0),
		.in_wire_0_1(horizontal_tile_31_19_to_tile_31_18_1),
		.in_wire_0_2(horizontal_tile_31_19_to_tile_31_18_2),
		.in_wire_0_3(horizontal_tile_31_19_to_tile_31_18_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1011)
	);

	pe_tile_bottom pe_tile_31_19(
		.out_wire_3_0(vertical_tile_31_19_to_tile_30_19_0),
		.out_wire_3_1(vertical_tile_31_19_to_tile_30_19_1),
		.out_wire_3_2(vertical_tile_31_19_to_tile_30_19_2),
		.out_wire_3_3(vertical_tile_31_19_to_tile_30_19_3),
		.in_wire_3_0(vertical_tile_30_19_to_tile_31_19_0),
		.in_wire_3_1(vertical_tile_30_19_to_tile_31_19_1),
		.in_wire_3_2(vertical_tile_30_19_to_tile_31_19_2),
		.in_wire_3_3(vertical_tile_30_19_to_tile_31_19_3),
		.out_wire_1_0(grid_to_output_19),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_19_to_tile_31_18_0),
		.out_wire_2_1(horizontal_tile_31_19_to_tile_31_18_1),
		.out_wire_2_2(horizontal_tile_31_19_to_tile_31_18_2),
		.out_wire_2_3(horizontal_tile_31_19_to_tile_31_18_3),
		.in_wire_2_0(horizontal_tile_31_18_to_tile_31_19_0),
		.in_wire_2_1(horizontal_tile_31_18_to_tile_31_19_1),
		.in_wire_2_2(horizontal_tile_31_18_to_tile_31_19_2),
		.in_wire_2_3(horizontal_tile_31_18_to_tile_31_19_3),
		.out_wire_0_0(horizontal_tile_31_19_to_tile_31_20_0),
		.out_wire_0_1(horizontal_tile_31_19_to_tile_31_20_1),
		.out_wire_0_2(horizontal_tile_31_19_to_tile_31_20_2),
		.out_wire_0_3(horizontal_tile_31_19_to_tile_31_20_3),
		.in_wire_0_0(horizontal_tile_31_20_to_tile_31_19_0),
		.in_wire_0_1(horizontal_tile_31_20_to_tile_31_19_1),
		.in_wire_0_2(horizontal_tile_31_20_to_tile_31_19_2),
		.in_wire_0_3(horizontal_tile_31_20_to_tile_31_19_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1012)
	);

	pe_tile_bottom pe_tile_31_20(
		.out_wire_3_0(vertical_tile_31_20_to_tile_30_20_0),
		.out_wire_3_1(vertical_tile_31_20_to_tile_30_20_1),
		.out_wire_3_2(vertical_tile_31_20_to_tile_30_20_2),
		.out_wire_3_3(vertical_tile_31_20_to_tile_30_20_3),
		.in_wire_3_0(vertical_tile_30_20_to_tile_31_20_0),
		.in_wire_3_1(vertical_tile_30_20_to_tile_31_20_1),
		.in_wire_3_2(vertical_tile_30_20_to_tile_31_20_2),
		.in_wire_3_3(vertical_tile_30_20_to_tile_31_20_3),
		.out_wire_1_0(grid_to_output_20),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_20_to_tile_31_19_0),
		.out_wire_2_1(horizontal_tile_31_20_to_tile_31_19_1),
		.out_wire_2_2(horizontal_tile_31_20_to_tile_31_19_2),
		.out_wire_2_3(horizontal_tile_31_20_to_tile_31_19_3),
		.in_wire_2_0(horizontal_tile_31_19_to_tile_31_20_0),
		.in_wire_2_1(horizontal_tile_31_19_to_tile_31_20_1),
		.in_wire_2_2(horizontal_tile_31_19_to_tile_31_20_2),
		.in_wire_2_3(horizontal_tile_31_19_to_tile_31_20_3),
		.out_wire_0_0(horizontal_tile_31_20_to_tile_31_21_0),
		.out_wire_0_1(horizontal_tile_31_20_to_tile_31_21_1),
		.out_wire_0_2(horizontal_tile_31_20_to_tile_31_21_2),
		.out_wire_0_3(horizontal_tile_31_20_to_tile_31_21_3),
		.in_wire_0_0(horizontal_tile_31_21_to_tile_31_20_0),
		.in_wire_0_1(horizontal_tile_31_21_to_tile_31_20_1),
		.in_wire_0_2(horizontal_tile_31_21_to_tile_31_20_2),
		.in_wire_0_3(horizontal_tile_31_21_to_tile_31_20_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1013)
	);

	pe_tile_bottom pe_tile_31_21(
		.out_wire_3_0(vertical_tile_31_21_to_tile_30_21_0),
		.out_wire_3_1(vertical_tile_31_21_to_tile_30_21_1),
		.out_wire_3_2(vertical_tile_31_21_to_tile_30_21_2),
		.out_wire_3_3(vertical_tile_31_21_to_tile_30_21_3),
		.in_wire_3_0(vertical_tile_30_21_to_tile_31_21_0),
		.in_wire_3_1(vertical_tile_30_21_to_tile_31_21_1),
		.in_wire_3_2(vertical_tile_30_21_to_tile_31_21_2),
		.in_wire_3_3(vertical_tile_30_21_to_tile_31_21_3),
		.out_wire_1_0(grid_to_output_21),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_21_to_tile_31_20_0),
		.out_wire_2_1(horizontal_tile_31_21_to_tile_31_20_1),
		.out_wire_2_2(horizontal_tile_31_21_to_tile_31_20_2),
		.out_wire_2_3(horizontal_tile_31_21_to_tile_31_20_3),
		.in_wire_2_0(horizontal_tile_31_20_to_tile_31_21_0),
		.in_wire_2_1(horizontal_tile_31_20_to_tile_31_21_1),
		.in_wire_2_2(horizontal_tile_31_20_to_tile_31_21_2),
		.in_wire_2_3(horizontal_tile_31_20_to_tile_31_21_3),
		.out_wire_0_0(horizontal_tile_31_21_to_tile_31_22_0),
		.out_wire_0_1(horizontal_tile_31_21_to_tile_31_22_1),
		.out_wire_0_2(horizontal_tile_31_21_to_tile_31_22_2),
		.out_wire_0_3(horizontal_tile_31_21_to_tile_31_22_3),
		.in_wire_0_0(horizontal_tile_31_22_to_tile_31_21_0),
		.in_wire_0_1(horizontal_tile_31_22_to_tile_31_21_1),
		.in_wire_0_2(horizontal_tile_31_22_to_tile_31_21_2),
		.in_wire_0_3(horizontal_tile_31_22_to_tile_31_21_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1014)
	);

	pe_tile_bottom pe_tile_31_22(
		.out_wire_3_0(vertical_tile_31_22_to_tile_30_22_0),
		.out_wire_3_1(vertical_tile_31_22_to_tile_30_22_1),
		.out_wire_3_2(vertical_tile_31_22_to_tile_30_22_2),
		.out_wire_3_3(vertical_tile_31_22_to_tile_30_22_3),
		.in_wire_3_0(vertical_tile_30_22_to_tile_31_22_0),
		.in_wire_3_1(vertical_tile_30_22_to_tile_31_22_1),
		.in_wire_3_2(vertical_tile_30_22_to_tile_31_22_2),
		.in_wire_3_3(vertical_tile_30_22_to_tile_31_22_3),
		.out_wire_1_0(grid_to_output_22),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_22_to_tile_31_21_0),
		.out_wire_2_1(horizontal_tile_31_22_to_tile_31_21_1),
		.out_wire_2_2(horizontal_tile_31_22_to_tile_31_21_2),
		.out_wire_2_3(horizontal_tile_31_22_to_tile_31_21_3),
		.in_wire_2_0(horizontal_tile_31_21_to_tile_31_22_0),
		.in_wire_2_1(horizontal_tile_31_21_to_tile_31_22_1),
		.in_wire_2_2(horizontal_tile_31_21_to_tile_31_22_2),
		.in_wire_2_3(horizontal_tile_31_21_to_tile_31_22_3),
		.out_wire_0_0(horizontal_tile_31_22_to_tile_31_23_0),
		.out_wire_0_1(horizontal_tile_31_22_to_tile_31_23_1),
		.out_wire_0_2(horizontal_tile_31_22_to_tile_31_23_2),
		.out_wire_0_3(horizontal_tile_31_22_to_tile_31_23_3),
		.in_wire_0_0(horizontal_tile_31_23_to_tile_31_22_0),
		.in_wire_0_1(horizontal_tile_31_23_to_tile_31_22_1),
		.in_wire_0_2(horizontal_tile_31_23_to_tile_31_22_2),
		.in_wire_0_3(horizontal_tile_31_23_to_tile_31_22_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1015)
	);

	pe_tile_bottom pe_tile_31_23(
		.out_wire_3_0(vertical_tile_31_23_to_tile_30_23_0),
		.out_wire_3_1(vertical_tile_31_23_to_tile_30_23_1),
		.out_wire_3_2(vertical_tile_31_23_to_tile_30_23_2),
		.out_wire_3_3(vertical_tile_31_23_to_tile_30_23_3),
		.in_wire_3_0(vertical_tile_30_23_to_tile_31_23_0),
		.in_wire_3_1(vertical_tile_30_23_to_tile_31_23_1),
		.in_wire_3_2(vertical_tile_30_23_to_tile_31_23_2),
		.in_wire_3_3(vertical_tile_30_23_to_tile_31_23_3),
		.out_wire_1_0(grid_to_output_23),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_23_to_tile_31_22_0),
		.out_wire_2_1(horizontal_tile_31_23_to_tile_31_22_1),
		.out_wire_2_2(horizontal_tile_31_23_to_tile_31_22_2),
		.out_wire_2_3(horizontal_tile_31_23_to_tile_31_22_3),
		.in_wire_2_0(horizontal_tile_31_22_to_tile_31_23_0),
		.in_wire_2_1(horizontal_tile_31_22_to_tile_31_23_1),
		.in_wire_2_2(horizontal_tile_31_22_to_tile_31_23_2),
		.in_wire_2_3(horizontal_tile_31_22_to_tile_31_23_3),
		.out_wire_0_0(horizontal_tile_31_23_to_tile_31_24_0),
		.out_wire_0_1(horizontal_tile_31_23_to_tile_31_24_1),
		.out_wire_0_2(horizontal_tile_31_23_to_tile_31_24_2),
		.out_wire_0_3(horizontal_tile_31_23_to_tile_31_24_3),
		.in_wire_0_0(horizontal_tile_31_24_to_tile_31_23_0),
		.in_wire_0_1(horizontal_tile_31_24_to_tile_31_23_1),
		.in_wire_0_2(horizontal_tile_31_24_to_tile_31_23_2),
		.in_wire_0_3(horizontal_tile_31_24_to_tile_31_23_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1016)
	);

	pe_tile_bottom pe_tile_31_24(
		.out_wire_3_0(vertical_tile_31_24_to_tile_30_24_0),
		.out_wire_3_1(vertical_tile_31_24_to_tile_30_24_1),
		.out_wire_3_2(vertical_tile_31_24_to_tile_30_24_2),
		.out_wire_3_3(vertical_tile_31_24_to_tile_30_24_3),
		.in_wire_3_0(vertical_tile_30_24_to_tile_31_24_0),
		.in_wire_3_1(vertical_tile_30_24_to_tile_31_24_1),
		.in_wire_3_2(vertical_tile_30_24_to_tile_31_24_2),
		.in_wire_3_3(vertical_tile_30_24_to_tile_31_24_3),
		.out_wire_1_0(grid_to_output_24),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_24_to_tile_31_23_0),
		.out_wire_2_1(horizontal_tile_31_24_to_tile_31_23_1),
		.out_wire_2_2(horizontal_tile_31_24_to_tile_31_23_2),
		.out_wire_2_3(horizontal_tile_31_24_to_tile_31_23_3),
		.in_wire_2_0(horizontal_tile_31_23_to_tile_31_24_0),
		.in_wire_2_1(horizontal_tile_31_23_to_tile_31_24_1),
		.in_wire_2_2(horizontal_tile_31_23_to_tile_31_24_2),
		.in_wire_2_3(horizontal_tile_31_23_to_tile_31_24_3),
		.out_wire_0_0(horizontal_tile_31_24_to_tile_31_25_0),
		.out_wire_0_1(horizontal_tile_31_24_to_tile_31_25_1),
		.out_wire_0_2(horizontal_tile_31_24_to_tile_31_25_2),
		.out_wire_0_3(horizontal_tile_31_24_to_tile_31_25_3),
		.in_wire_0_0(horizontal_tile_31_25_to_tile_31_24_0),
		.in_wire_0_1(horizontal_tile_31_25_to_tile_31_24_1),
		.in_wire_0_2(horizontal_tile_31_25_to_tile_31_24_2),
		.in_wire_0_3(horizontal_tile_31_25_to_tile_31_24_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1017)
	);

	pe_tile_bottom pe_tile_31_25(
		.out_wire_3_0(vertical_tile_31_25_to_tile_30_25_0),
		.out_wire_3_1(vertical_tile_31_25_to_tile_30_25_1),
		.out_wire_3_2(vertical_tile_31_25_to_tile_30_25_2),
		.out_wire_3_3(vertical_tile_31_25_to_tile_30_25_3),
		.in_wire_3_0(vertical_tile_30_25_to_tile_31_25_0),
		.in_wire_3_1(vertical_tile_30_25_to_tile_31_25_1),
		.in_wire_3_2(vertical_tile_30_25_to_tile_31_25_2),
		.in_wire_3_3(vertical_tile_30_25_to_tile_31_25_3),
		.out_wire_1_0(grid_to_output_25),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_25_to_tile_31_24_0),
		.out_wire_2_1(horizontal_tile_31_25_to_tile_31_24_1),
		.out_wire_2_2(horizontal_tile_31_25_to_tile_31_24_2),
		.out_wire_2_3(horizontal_tile_31_25_to_tile_31_24_3),
		.in_wire_2_0(horizontal_tile_31_24_to_tile_31_25_0),
		.in_wire_2_1(horizontal_tile_31_24_to_tile_31_25_1),
		.in_wire_2_2(horizontal_tile_31_24_to_tile_31_25_2),
		.in_wire_2_3(horizontal_tile_31_24_to_tile_31_25_3),
		.out_wire_0_0(horizontal_tile_31_25_to_tile_31_26_0),
		.out_wire_0_1(horizontal_tile_31_25_to_tile_31_26_1),
		.out_wire_0_2(horizontal_tile_31_25_to_tile_31_26_2),
		.out_wire_0_3(horizontal_tile_31_25_to_tile_31_26_3),
		.in_wire_0_0(horizontal_tile_31_26_to_tile_31_25_0),
		.in_wire_0_1(horizontal_tile_31_26_to_tile_31_25_1),
		.in_wire_0_2(horizontal_tile_31_26_to_tile_31_25_2),
		.in_wire_0_3(horizontal_tile_31_26_to_tile_31_25_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1018)
	);

	pe_tile_bottom pe_tile_31_26(
		.out_wire_3_0(vertical_tile_31_26_to_tile_30_26_0),
		.out_wire_3_1(vertical_tile_31_26_to_tile_30_26_1),
		.out_wire_3_2(vertical_tile_31_26_to_tile_30_26_2),
		.out_wire_3_3(vertical_tile_31_26_to_tile_30_26_3),
		.in_wire_3_0(vertical_tile_30_26_to_tile_31_26_0),
		.in_wire_3_1(vertical_tile_30_26_to_tile_31_26_1),
		.in_wire_3_2(vertical_tile_30_26_to_tile_31_26_2),
		.in_wire_3_3(vertical_tile_30_26_to_tile_31_26_3),
		.out_wire_1_0(grid_to_output_26),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_26_to_tile_31_25_0),
		.out_wire_2_1(horizontal_tile_31_26_to_tile_31_25_1),
		.out_wire_2_2(horizontal_tile_31_26_to_tile_31_25_2),
		.out_wire_2_3(horizontal_tile_31_26_to_tile_31_25_3),
		.in_wire_2_0(horizontal_tile_31_25_to_tile_31_26_0),
		.in_wire_2_1(horizontal_tile_31_25_to_tile_31_26_1),
		.in_wire_2_2(horizontal_tile_31_25_to_tile_31_26_2),
		.in_wire_2_3(horizontal_tile_31_25_to_tile_31_26_3),
		.out_wire_0_0(horizontal_tile_31_26_to_tile_31_27_0),
		.out_wire_0_1(horizontal_tile_31_26_to_tile_31_27_1),
		.out_wire_0_2(horizontal_tile_31_26_to_tile_31_27_2),
		.out_wire_0_3(horizontal_tile_31_26_to_tile_31_27_3),
		.in_wire_0_0(horizontal_tile_31_27_to_tile_31_26_0),
		.in_wire_0_1(horizontal_tile_31_27_to_tile_31_26_1),
		.in_wire_0_2(horizontal_tile_31_27_to_tile_31_26_2),
		.in_wire_0_3(horizontal_tile_31_27_to_tile_31_26_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1019)
	);

	pe_tile_bottom pe_tile_31_27(
		.out_wire_3_0(vertical_tile_31_27_to_tile_30_27_0),
		.out_wire_3_1(vertical_tile_31_27_to_tile_30_27_1),
		.out_wire_3_2(vertical_tile_31_27_to_tile_30_27_2),
		.out_wire_3_3(vertical_tile_31_27_to_tile_30_27_3),
		.in_wire_3_0(vertical_tile_30_27_to_tile_31_27_0),
		.in_wire_3_1(vertical_tile_30_27_to_tile_31_27_1),
		.in_wire_3_2(vertical_tile_30_27_to_tile_31_27_2),
		.in_wire_3_3(vertical_tile_30_27_to_tile_31_27_3),
		.out_wire_1_0(grid_to_output_27),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_27_to_tile_31_26_0),
		.out_wire_2_1(horizontal_tile_31_27_to_tile_31_26_1),
		.out_wire_2_2(horizontal_tile_31_27_to_tile_31_26_2),
		.out_wire_2_3(horizontal_tile_31_27_to_tile_31_26_3),
		.in_wire_2_0(horizontal_tile_31_26_to_tile_31_27_0),
		.in_wire_2_1(horizontal_tile_31_26_to_tile_31_27_1),
		.in_wire_2_2(horizontal_tile_31_26_to_tile_31_27_2),
		.in_wire_2_3(horizontal_tile_31_26_to_tile_31_27_3),
		.out_wire_0_0(horizontal_tile_31_27_to_tile_31_28_0),
		.out_wire_0_1(horizontal_tile_31_27_to_tile_31_28_1),
		.out_wire_0_2(horizontal_tile_31_27_to_tile_31_28_2),
		.out_wire_0_3(horizontal_tile_31_27_to_tile_31_28_3),
		.in_wire_0_0(horizontal_tile_31_28_to_tile_31_27_0),
		.in_wire_0_1(horizontal_tile_31_28_to_tile_31_27_1),
		.in_wire_0_2(horizontal_tile_31_28_to_tile_31_27_2),
		.in_wire_0_3(horizontal_tile_31_28_to_tile_31_27_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1020)
	);

	pe_tile_bottom pe_tile_31_28(
		.out_wire_3_0(vertical_tile_31_28_to_tile_30_28_0),
		.out_wire_3_1(vertical_tile_31_28_to_tile_30_28_1),
		.out_wire_3_2(vertical_tile_31_28_to_tile_30_28_2),
		.out_wire_3_3(vertical_tile_31_28_to_tile_30_28_3),
		.in_wire_3_0(vertical_tile_30_28_to_tile_31_28_0),
		.in_wire_3_1(vertical_tile_30_28_to_tile_31_28_1),
		.in_wire_3_2(vertical_tile_30_28_to_tile_31_28_2),
		.in_wire_3_3(vertical_tile_30_28_to_tile_31_28_3),
		.out_wire_1_0(grid_to_output_28),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_28_to_tile_31_27_0),
		.out_wire_2_1(horizontal_tile_31_28_to_tile_31_27_1),
		.out_wire_2_2(horizontal_tile_31_28_to_tile_31_27_2),
		.out_wire_2_3(horizontal_tile_31_28_to_tile_31_27_3),
		.in_wire_2_0(horizontal_tile_31_27_to_tile_31_28_0),
		.in_wire_2_1(horizontal_tile_31_27_to_tile_31_28_1),
		.in_wire_2_2(horizontal_tile_31_27_to_tile_31_28_2),
		.in_wire_2_3(horizontal_tile_31_27_to_tile_31_28_3),
		.out_wire_0_0(horizontal_tile_31_28_to_tile_31_29_0),
		.out_wire_0_1(horizontal_tile_31_28_to_tile_31_29_1),
		.out_wire_0_2(horizontal_tile_31_28_to_tile_31_29_2),
		.out_wire_0_3(horizontal_tile_31_28_to_tile_31_29_3),
		.in_wire_0_0(horizontal_tile_31_29_to_tile_31_28_0),
		.in_wire_0_1(horizontal_tile_31_29_to_tile_31_28_1),
		.in_wire_0_2(horizontal_tile_31_29_to_tile_31_28_2),
		.in_wire_0_3(horizontal_tile_31_29_to_tile_31_28_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1021)
	);

	pe_tile_bottom pe_tile_31_29(
		.out_wire_3_0(vertical_tile_31_29_to_tile_30_29_0),
		.out_wire_3_1(vertical_tile_31_29_to_tile_30_29_1),
		.out_wire_3_2(vertical_tile_31_29_to_tile_30_29_2),
		.out_wire_3_3(vertical_tile_31_29_to_tile_30_29_3),
		.in_wire_3_0(vertical_tile_30_29_to_tile_31_29_0),
		.in_wire_3_1(vertical_tile_30_29_to_tile_31_29_1),
		.in_wire_3_2(vertical_tile_30_29_to_tile_31_29_2),
		.in_wire_3_3(vertical_tile_30_29_to_tile_31_29_3),
		.out_wire_1_0(grid_to_output_29),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_29_to_tile_31_28_0),
		.out_wire_2_1(horizontal_tile_31_29_to_tile_31_28_1),
		.out_wire_2_2(horizontal_tile_31_29_to_tile_31_28_2),
		.out_wire_2_3(horizontal_tile_31_29_to_tile_31_28_3),
		.in_wire_2_0(horizontal_tile_31_28_to_tile_31_29_0),
		.in_wire_2_1(horizontal_tile_31_28_to_tile_31_29_1),
		.in_wire_2_2(horizontal_tile_31_28_to_tile_31_29_2),
		.in_wire_2_3(horizontal_tile_31_28_to_tile_31_29_3),
		.out_wire_0_0(horizontal_tile_31_29_to_tile_31_30_0),
		.out_wire_0_1(horizontal_tile_31_29_to_tile_31_30_1),
		.out_wire_0_2(horizontal_tile_31_29_to_tile_31_30_2),
		.out_wire_0_3(horizontal_tile_31_29_to_tile_31_30_3),
		.in_wire_0_0(horizontal_tile_31_30_to_tile_31_29_0),
		.in_wire_0_1(horizontal_tile_31_30_to_tile_31_29_1),
		.in_wire_0_2(horizontal_tile_31_30_to_tile_31_29_2),
		.in_wire_0_3(horizontal_tile_31_30_to_tile_31_29_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1022)
	);

	pe_tile_bottom pe_tile_31_30(
		.out_wire_3_0(vertical_tile_31_30_to_tile_30_30_0),
		.out_wire_3_1(vertical_tile_31_30_to_tile_30_30_1),
		.out_wire_3_2(vertical_tile_31_30_to_tile_30_30_2),
		.out_wire_3_3(vertical_tile_31_30_to_tile_30_30_3),
		.in_wire_3_0(vertical_tile_30_30_to_tile_31_30_0),
		.in_wire_3_1(vertical_tile_30_30_to_tile_31_30_1),
		.in_wire_3_2(vertical_tile_30_30_to_tile_31_30_2),
		.in_wire_3_3(vertical_tile_30_30_to_tile_31_30_3),
		.out_wire_1_0(grid_to_output_30),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_30_to_tile_31_29_0),
		.out_wire_2_1(horizontal_tile_31_30_to_tile_31_29_1),
		.out_wire_2_2(horizontal_tile_31_30_to_tile_31_29_2),
		.out_wire_2_3(horizontal_tile_31_30_to_tile_31_29_3),
		.in_wire_2_0(horizontal_tile_31_29_to_tile_31_30_0),
		.in_wire_2_1(horizontal_tile_31_29_to_tile_31_30_1),
		.in_wire_2_2(horizontal_tile_31_29_to_tile_31_30_2),
		.in_wire_2_3(horizontal_tile_31_29_to_tile_31_30_3),
		.out_wire_0_0(horizontal_tile_31_30_to_tile_31_31_0),
		.out_wire_0_1(horizontal_tile_31_30_to_tile_31_31_1),
		.out_wire_0_2(horizontal_tile_31_30_to_tile_31_31_2),
		.out_wire_0_3(horizontal_tile_31_30_to_tile_31_31_3),
		.in_wire_0_0(horizontal_tile_31_31_to_tile_31_30_0),
		.in_wire_0_1(horizontal_tile_31_31_to_tile_31_30_1),
		.in_wire_0_2(horizontal_tile_31_31_to_tile_31_30_2),
		.in_wire_0_3(horizontal_tile_31_31_to_tile_31_30_3),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1023)
	);

	pe_tile_bottom_right pe_tile_31_31(
		.out_wire_3_0(vertical_tile_31_31_to_tile_30_31_0),
		.out_wire_3_1(vertical_tile_31_31_to_tile_30_31_1),
		.out_wire_3_2(vertical_tile_31_31_to_tile_30_31_2),
		.out_wire_3_3(vertical_tile_31_31_to_tile_30_31_3),
		.in_wire_3_0(vertical_tile_30_31_to_tile_31_31_0),
		.in_wire_3_1(vertical_tile_30_31_to_tile_31_31_1),
		.in_wire_3_2(vertical_tile_30_31_to_tile_31_31_2),
		.in_wire_3_3(vertical_tile_30_31_to_tile_31_31_3),
		.out_wire_1_0(grid_to_output_31),
		.in_wire_1_0(1'b0),
		.in_wire_1_1(1'b0),
		.in_wire_1_2(1'b0),
		.in_wire_1_3(1'b0),
		.out_wire_2_0(horizontal_tile_31_31_to_tile_31_30_0),
		.out_wire_2_1(horizontal_tile_31_31_to_tile_31_30_1),
		.out_wire_2_2(horizontal_tile_31_31_to_tile_31_30_2),
		.out_wire_2_3(horizontal_tile_31_31_to_tile_31_30_3),
		.in_wire_2_0(horizontal_tile_31_30_to_tile_31_31_0),
		.in_wire_2_1(horizontal_tile_31_30_to_tile_31_31_1),
		.in_wire_2_2(horizontal_tile_31_30_to_tile_31_31_2),
		.in_wire_2_3(horizontal_tile_31_30_to_tile_31_31_3),
		.in_wire_0_0(1'b0),
		.in_wire_0_1(1'b0),
		.in_wire_0_2(1'b0),
		.in_wire_0_3(1'b0),
		.clk(clk),
		.reset(reset),
		.config_addr(config_addr),
		.config_data(config_data),
		.tile_id(1024)
	);



endmodule