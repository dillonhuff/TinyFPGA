module connect_box();


endmodule; // connect_box
