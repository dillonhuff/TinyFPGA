
//                2
//
// 
//  3        switch_box        1
//
//                
//                0

module switch_box(input clk,
                  input rst,

                  // Vertical tracks
                  input side_0_track_0_in,
                  input side_0_track_1_in,
                  input side_0_track_2_in,
                  input side_0_track_3_in,

                  input side_1_track_0_in,
                  input side_1_track_1_in,
                  input side_1_track_2_in,
                  input side_1_track_3_in,

                  input side_2_track_0_in,
                  input side_2_track_1_in,
                  input side_2_track_2_in,
                  input side_2_track_3_in,

                  input side_3_track_0_in,
                  input side_3_track_1_in,
                  input side_3_track_2_in,
                  input side_3_track_3_in,

                  );

   
endmodule
