module connect_box(
                   input  track0_in,
                   input  track1_in,
                   input  track2_in,
                   input  track3_in,

                   input  track0_out,
                   input  track1_out,
                   input  track2_out,
                   input  track3_out,
                   
                   output block_out
                   
                   );

   
   
   
endmodule; // connect_box
